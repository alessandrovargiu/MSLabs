
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_top_entity is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_top_entity;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_entity.all;

entity register_file_nbit32_addr_bits5 is

   port( CLK, RESET, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
         ADD_RD2 : in std_logic_vector (4 downto 0);  DATAIN : in 
         std_logic_vector (31 downto 0);  OUT1, OUT2 : out std_logic_vector (31
         downto 0));

end register_file_nbit32_addr_bits5;

architecture SYN_Behavioral of register_file_nbit32_addr_bits5 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X4
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component TBUF_X1
      port( A, EN : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal REGISTERS_0_31_port, REGISTERS_0_30_port, REGISTERS_0_29_port, 
      REGISTERS_0_28_port, REGISTERS_0_27_port, REGISTERS_0_26_port, 
      REGISTERS_0_25_port, REGISTERS_0_24_port, REGISTERS_0_23_port, 
      REGISTERS_0_22_port, REGISTERS_0_21_port, REGISTERS_0_20_port, 
      REGISTERS_0_19_port, REGISTERS_0_18_port, REGISTERS_0_17_port, 
      REGISTERS_0_16_port, REGISTERS_0_15_port, REGISTERS_0_14_port, 
      REGISTERS_0_13_port, REGISTERS_0_12_port, REGISTERS_0_11_port, 
      REGISTERS_0_10_port, REGISTERS_0_9_port, REGISTERS_0_8_port, 
      REGISTERS_0_7_port, REGISTERS_0_6_port, REGISTERS_0_5_port, 
      REGISTERS_0_4_port, REGISTERS_0_3_port, REGISTERS_0_2_port, 
      REGISTERS_0_1_port, REGISTERS_0_0_port, REGISTERS_1_31_port, 
      REGISTERS_1_30_port, REGISTERS_1_29_port, REGISTERS_1_28_port, 
      REGISTERS_1_27_port, REGISTERS_1_26_port, REGISTERS_1_25_port, 
      REGISTERS_1_24_port, REGISTERS_1_23_port, REGISTERS_1_22_port, 
      REGISTERS_1_21_port, REGISTERS_1_20_port, REGISTERS_1_19_port, 
      REGISTERS_1_18_port, REGISTERS_1_17_port, REGISTERS_1_16_port, 
      REGISTERS_1_15_port, REGISTERS_1_14_port, REGISTERS_1_13_port, 
      REGISTERS_1_12_port, REGISTERS_1_11_port, REGISTERS_1_10_port, 
      REGISTERS_1_9_port, REGISTERS_1_8_port, REGISTERS_1_7_port, 
      REGISTERS_1_6_port, REGISTERS_1_5_port, REGISTERS_1_4_port, 
      REGISTERS_1_3_port, REGISTERS_1_2_port, REGISTERS_1_1_port, 
      REGISTERS_1_0_port, REGISTERS_2_31_port, REGISTERS_2_30_port, 
      REGISTERS_2_29_port, REGISTERS_2_28_port, REGISTERS_2_27_port, 
      REGISTERS_2_26_port, REGISTERS_2_25_port, REGISTERS_2_24_port, 
      REGISTERS_2_23_port, REGISTERS_2_22_port, REGISTERS_2_21_port, 
      REGISTERS_2_20_port, REGISTERS_2_19_port, REGISTERS_2_18_port, 
      REGISTERS_2_17_port, REGISTERS_2_16_port, REGISTERS_2_15_port, 
      REGISTERS_2_14_port, REGISTERS_2_13_port, REGISTERS_2_12_port, 
      REGISTERS_2_11_port, REGISTERS_2_10_port, REGISTERS_2_9_port, 
      REGISTERS_2_8_port, REGISTERS_2_7_port, REGISTERS_2_6_port, 
      REGISTERS_2_5_port, REGISTERS_2_4_port, REGISTERS_2_3_port, 
      REGISTERS_2_2_port, REGISTERS_2_1_port, REGISTERS_2_0_port, 
      REGISTERS_3_31_port, REGISTERS_3_30_port, REGISTERS_3_29_port, 
      REGISTERS_3_28_port, REGISTERS_3_27_port, REGISTERS_3_26_port, 
      REGISTERS_3_25_port, REGISTERS_3_24_port, REGISTERS_3_23_port, 
      REGISTERS_3_22_port, REGISTERS_3_21_port, REGISTERS_3_20_port, 
      REGISTERS_3_19_port, REGISTERS_3_18_port, REGISTERS_3_17_port, 
      REGISTERS_3_16_port, REGISTERS_3_15_port, REGISTERS_3_14_port, 
      REGISTERS_3_13_port, REGISTERS_3_12_port, REGISTERS_3_11_port, 
      REGISTERS_3_10_port, REGISTERS_3_9_port, REGISTERS_3_8_port, 
      REGISTERS_3_7_port, REGISTERS_3_6_port, REGISTERS_3_5_port, 
      REGISTERS_3_4_port, REGISTERS_3_3_port, REGISTERS_3_2_port, 
      REGISTERS_3_1_port, REGISTERS_3_0_port, REGISTERS_4_31_port, 
      REGISTERS_4_30_port, REGISTERS_4_29_port, REGISTERS_4_28_port, 
      REGISTERS_4_27_port, REGISTERS_4_26_port, REGISTERS_4_25_port, 
      REGISTERS_4_24_port, REGISTERS_4_23_port, REGISTERS_4_22_port, 
      REGISTERS_4_21_port, REGISTERS_4_20_port, REGISTERS_4_19_port, 
      REGISTERS_4_18_port, REGISTERS_4_17_port, REGISTERS_4_16_port, 
      REGISTERS_4_15_port, REGISTERS_4_14_port, REGISTERS_4_13_port, 
      REGISTERS_4_12_port, REGISTERS_4_11_port, REGISTERS_4_10_port, 
      REGISTERS_4_9_port, REGISTERS_4_8_port, REGISTERS_4_7_port, 
      REGISTERS_4_6_port, REGISTERS_4_5_port, REGISTERS_4_4_port, 
      REGISTERS_4_3_port, REGISTERS_4_2_port, REGISTERS_4_1_port, 
      REGISTERS_4_0_port, REGISTERS_5_31_port, REGISTERS_5_30_port, 
      REGISTERS_5_29_port, REGISTERS_5_28_port, REGISTERS_5_27_port, 
      REGISTERS_5_26_port, REGISTERS_5_25_port, REGISTERS_5_24_port, 
      REGISTERS_5_23_port, REGISTERS_5_22_port, REGISTERS_5_21_port, 
      REGISTERS_5_20_port, REGISTERS_5_19_port, REGISTERS_5_18_port, 
      REGISTERS_5_17_port, REGISTERS_5_16_port, REGISTERS_5_15_port, 
      REGISTERS_5_14_port, REGISTERS_5_13_port, REGISTERS_5_12_port, 
      REGISTERS_5_11_port, REGISTERS_5_10_port, REGISTERS_5_9_port, 
      REGISTERS_5_8_port, REGISTERS_5_7_port, REGISTERS_5_6_port, 
      REGISTERS_5_5_port, REGISTERS_5_4_port, REGISTERS_5_3_port, 
      REGISTERS_5_2_port, REGISTERS_5_1_port, REGISTERS_5_0_port, 
      REGISTERS_6_31_port, REGISTERS_6_30_port, REGISTERS_6_29_port, 
      REGISTERS_6_28_port, REGISTERS_6_27_port, REGISTERS_6_26_port, 
      REGISTERS_6_25_port, REGISTERS_6_24_port, REGISTERS_6_23_port, 
      REGISTERS_6_22_port, REGISTERS_6_21_port, REGISTERS_6_20_port, 
      REGISTERS_6_19_port, REGISTERS_6_18_port, REGISTERS_6_17_port, 
      REGISTERS_6_16_port, REGISTERS_6_15_port, REGISTERS_6_14_port, 
      REGISTERS_6_13_port, REGISTERS_6_12_port, REGISTERS_6_11_port, 
      REGISTERS_6_10_port, REGISTERS_6_9_port, REGISTERS_6_8_port, 
      REGISTERS_6_7_port, REGISTERS_6_6_port, REGISTERS_6_5_port, 
      REGISTERS_6_4_port, REGISTERS_6_3_port, REGISTERS_6_2_port, 
      REGISTERS_6_1_port, REGISTERS_6_0_port, REGISTERS_7_31_port, 
      REGISTERS_7_30_port, REGISTERS_7_29_port, REGISTERS_7_28_port, 
      REGISTERS_7_27_port, REGISTERS_7_26_port, REGISTERS_7_25_port, 
      REGISTERS_7_24_port, REGISTERS_7_23_port, REGISTERS_7_22_port, 
      REGISTERS_7_21_port, REGISTERS_7_20_port, REGISTERS_7_19_port, 
      REGISTERS_7_18_port, REGISTERS_7_17_port, REGISTERS_7_16_port, 
      REGISTERS_7_15_port, REGISTERS_7_14_port, REGISTERS_7_13_port, 
      REGISTERS_7_12_port, REGISTERS_7_11_port, REGISTERS_7_10_port, 
      REGISTERS_7_9_port, REGISTERS_7_8_port, REGISTERS_7_7_port, 
      REGISTERS_7_6_port, REGISTERS_7_5_port, REGISTERS_7_4_port, 
      REGISTERS_7_3_port, REGISTERS_7_2_port, REGISTERS_7_1_port, 
      REGISTERS_7_0_port, REGISTERS_8_31_port, REGISTERS_8_30_port, 
      REGISTERS_8_29_port, REGISTERS_8_28_port, REGISTERS_8_27_port, 
      REGISTERS_8_26_port, REGISTERS_8_25_port, REGISTERS_8_24_port, 
      REGISTERS_8_23_port, REGISTERS_8_22_port, REGISTERS_8_21_port, 
      REGISTERS_8_20_port, REGISTERS_8_19_port, REGISTERS_8_18_port, 
      REGISTERS_8_17_port, REGISTERS_8_16_port, REGISTERS_8_15_port, 
      REGISTERS_8_14_port, REGISTERS_8_13_port, REGISTERS_8_12_port, 
      REGISTERS_8_11_port, REGISTERS_8_10_port, REGISTERS_8_9_port, 
      REGISTERS_8_8_port, REGISTERS_8_7_port, REGISTERS_8_6_port, 
      REGISTERS_8_5_port, REGISTERS_8_4_port, REGISTERS_8_3_port, 
      REGISTERS_8_2_port, REGISTERS_8_1_port, REGISTERS_8_0_port, 
      REGISTERS_9_31_port, REGISTERS_9_30_port, REGISTERS_9_29_port, 
      REGISTERS_9_28_port, REGISTERS_9_27_port, REGISTERS_9_26_port, 
      REGISTERS_9_25_port, REGISTERS_9_24_port, REGISTERS_9_23_port, 
      REGISTERS_9_22_port, REGISTERS_9_21_port, REGISTERS_9_20_port, 
      REGISTERS_9_19_port, REGISTERS_9_18_port, REGISTERS_9_17_port, 
      REGISTERS_9_16_port, REGISTERS_9_15_port, REGISTERS_9_14_port, 
      REGISTERS_9_13_port, REGISTERS_9_12_port, REGISTERS_9_11_port, 
      REGISTERS_9_10_port, REGISTERS_9_9_port, REGISTERS_9_8_port, 
      REGISTERS_9_7_port, REGISTERS_9_6_port, REGISTERS_9_5_port, 
      REGISTERS_9_4_port, REGISTERS_9_3_port, REGISTERS_9_2_port, 
      REGISTERS_9_1_port, REGISTERS_9_0_port, REGISTERS_10_31_port, 
      REGISTERS_10_30_port, REGISTERS_10_29_port, REGISTERS_10_28_port, 
      REGISTERS_10_27_port, REGISTERS_10_26_port, REGISTERS_10_25_port, 
      REGISTERS_10_24_port, REGISTERS_10_23_port, REGISTERS_10_22_port, 
      REGISTERS_10_21_port, REGISTERS_10_20_port, REGISTERS_10_19_port, 
      REGISTERS_10_18_port, REGISTERS_10_17_port, REGISTERS_10_16_port, 
      REGISTERS_10_15_port, REGISTERS_10_14_port, REGISTERS_10_13_port, 
      REGISTERS_10_12_port, REGISTERS_10_11_port, REGISTERS_10_10_port, 
      REGISTERS_10_9_port, REGISTERS_10_8_port, REGISTERS_10_7_port, 
      REGISTERS_10_6_port, REGISTERS_10_5_port, REGISTERS_10_4_port, 
      REGISTERS_10_3_port, REGISTERS_10_2_port, REGISTERS_10_1_port, 
      REGISTERS_10_0_port, REGISTERS_11_31_port, REGISTERS_11_30_port, 
      REGISTERS_11_29_port, REGISTERS_11_28_port, REGISTERS_11_27_port, 
      REGISTERS_11_26_port, REGISTERS_11_25_port, REGISTERS_11_24_port, 
      REGISTERS_11_23_port, REGISTERS_11_22_port, REGISTERS_11_21_port, 
      REGISTERS_11_20_port, REGISTERS_11_19_port, REGISTERS_11_18_port, 
      REGISTERS_11_17_port, REGISTERS_11_16_port, REGISTERS_11_15_port, 
      REGISTERS_11_14_port, REGISTERS_11_13_port, REGISTERS_11_12_port, 
      REGISTERS_11_11_port, REGISTERS_11_10_port, REGISTERS_11_9_port, 
      REGISTERS_11_8_port, REGISTERS_11_7_port, REGISTERS_11_6_port, 
      REGISTERS_11_5_port, REGISTERS_11_4_port, REGISTERS_11_3_port, 
      REGISTERS_11_2_port, REGISTERS_11_1_port, REGISTERS_11_0_port, 
      REGISTERS_12_31_port, REGISTERS_12_30_port, REGISTERS_12_29_port, 
      REGISTERS_12_28_port, REGISTERS_12_27_port, REGISTERS_12_26_port, 
      REGISTERS_12_25_port, REGISTERS_12_24_port, REGISTERS_12_23_port, 
      REGISTERS_12_22_port, REGISTERS_12_21_port, REGISTERS_12_20_port, 
      REGISTERS_12_19_port, REGISTERS_12_18_port, REGISTERS_12_17_port, 
      REGISTERS_12_16_port, REGISTERS_12_15_port, REGISTERS_12_14_port, 
      REGISTERS_12_13_port, REGISTERS_12_12_port, REGISTERS_12_11_port, 
      REGISTERS_12_10_port, REGISTERS_12_9_port, REGISTERS_12_8_port, 
      REGISTERS_12_7_port, REGISTERS_12_6_port, REGISTERS_12_5_port, 
      REGISTERS_12_4_port, REGISTERS_12_3_port, REGISTERS_12_2_port, 
      REGISTERS_12_1_port, REGISTERS_12_0_port, REGISTERS_13_31_port, 
      REGISTERS_13_30_port, REGISTERS_13_29_port, REGISTERS_13_28_port, 
      REGISTERS_13_27_port, REGISTERS_13_26_port, REGISTERS_13_25_port, 
      REGISTERS_13_24_port, REGISTERS_13_23_port, REGISTERS_13_22_port, 
      REGISTERS_13_21_port, REGISTERS_13_20_port, REGISTERS_13_19_port, 
      REGISTERS_13_18_port, REGISTERS_13_17_port, REGISTERS_13_16_port, 
      REGISTERS_13_15_port, REGISTERS_13_14_port, REGISTERS_13_13_port, 
      REGISTERS_13_12_port, REGISTERS_13_11_port, REGISTERS_13_10_port, 
      REGISTERS_13_9_port, REGISTERS_13_8_port, REGISTERS_13_7_port, 
      REGISTERS_13_6_port, REGISTERS_13_5_port, REGISTERS_13_4_port, 
      REGISTERS_13_3_port, REGISTERS_13_2_port, REGISTERS_13_1_port, 
      REGISTERS_13_0_port, REGISTERS_14_31_port, REGISTERS_14_30_port, 
      REGISTERS_14_29_port, REGISTERS_14_28_port, REGISTERS_14_27_port, 
      REGISTERS_14_26_port, REGISTERS_14_25_port, REGISTERS_14_24_port, 
      REGISTERS_14_23_port, REGISTERS_14_22_port, REGISTERS_14_21_port, 
      REGISTERS_14_20_port, REGISTERS_14_19_port, REGISTERS_14_18_port, 
      REGISTERS_14_17_port, REGISTERS_14_16_port, REGISTERS_14_15_port, 
      REGISTERS_14_14_port, REGISTERS_14_13_port, REGISTERS_14_12_port, 
      REGISTERS_14_11_port, REGISTERS_14_10_port, REGISTERS_14_9_port, 
      REGISTERS_14_8_port, REGISTERS_14_7_port, REGISTERS_14_6_port, 
      REGISTERS_14_5_port, REGISTERS_14_4_port, REGISTERS_14_3_port, 
      REGISTERS_14_2_port, REGISTERS_14_1_port, REGISTERS_14_0_port, 
      REGISTERS_15_31_port, REGISTERS_15_30_port, REGISTERS_15_29_port, 
      REGISTERS_15_28_port, REGISTERS_15_27_port, REGISTERS_15_26_port, 
      REGISTERS_15_25_port, REGISTERS_15_24_port, REGISTERS_15_23_port, 
      REGISTERS_15_22_port, REGISTERS_15_21_port, REGISTERS_15_20_port, 
      REGISTERS_15_19_port, REGISTERS_15_18_port, REGISTERS_15_17_port, 
      REGISTERS_15_16_port, REGISTERS_15_15_port, REGISTERS_15_14_port, 
      REGISTERS_15_13_port, REGISTERS_15_12_port, REGISTERS_15_11_port, 
      REGISTERS_15_10_port, REGISTERS_15_9_port, REGISTERS_15_8_port, 
      REGISTERS_15_7_port, REGISTERS_15_6_port, REGISTERS_15_5_port, 
      REGISTERS_15_4_port, REGISTERS_15_3_port, REGISTERS_15_2_port, 
      REGISTERS_15_1_port, REGISTERS_15_0_port, REGISTERS_16_31_port, 
      REGISTERS_16_30_port, REGISTERS_16_29_port, REGISTERS_16_28_port, 
      REGISTERS_16_27_port, REGISTERS_16_26_port, REGISTERS_16_25_port, 
      REGISTERS_16_24_port, REGISTERS_16_23_port, REGISTERS_16_22_port, 
      REGISTERS_16_21_port, REGISTERS_16_20_port, REGISTERS_16_19_port, 
      REGISTERS_16_18_port, REGISTERS_16_17_port, REGISTERS_16_16_port, 
      REGISTERS_16_15_port, REGISTERS_16_14_port, REGISTERS_16_13_port, 
      REGISTERS_16_12_port, REGISTERS_16_11_port, REGISTERS_16_10_port, 
      REGISTERS_16_9_port, REGISTERS_16_8_port, REGISTERS_16_7_port, 
      REGISTERS_16_6_port, REGISTERS_16_5_port, REGISTERS_16_4_port, 
      REGISTERS_16_3_port, REGISTERS_16_2_port, REGISTERS_16_1_port, 
      REGISTERS_16_0_port, REGISTERS_17_31_port, REGISTERS_17_30_port, 
      REGISTERS_17_29_port, REGISTERS_17_28_port, REGISTERS_17_27_port, 
      REGISTERS_17_26_port, REGISTERS_17_25_port, REGISTERS_17_24_port, 
      REGISTERS_17_23_port, REGISTERS_17_22_port, REGISTERS_17_21_port, 
      REGISTERS_17_20_port, REGISTERS_17_19_port, REGISTERS_17_18_port, 
      REGISTERS_17_17_port, REGISTERS_17_16_port, REGISTERS_17_15_port, 
      REGISTERS_17_14_port, REGISTERS_17_13_port, REGISTERS_17_12_port, 
      REGISTERS_17_11_port, REGISTERS_17_10_port, REGISTERS_17_9_port, 
      REGISTERS_17_8_port, REGISTERS_17_7_port, REGISTERS_17_6_port, 
      REGISTERS_17_5_port, REGISTERS_17_4_port, REGISTERS_17_3_port, 
      REGISTERS_17_2_port, REGISTERS_17_1_port, REGISTERS_17_0_port, 
      REGISTERS_18_31_port, REGISTERS_18_30_port, REGISTERS_18_29_port, 
      REGISTERS_18_28_port, REGISTERS_18_27_port, REGISTERS_18_26_port, 
      REGISTERS_18_25_port, REGISTERS_18_24_port, REGISTERS_18_23_port, 
      REGISTERS_18_22_port, REGISTERS_18_21_port, REGISTERS_18_20_port, 
      REGISTERS_18_19_port, REGISTERS_18_18_port, REGISTERS_18_17_port, 
      REGISTERS_18_16_port, REGISTERS_18_15_port, REGISTERS_18_14_port, 
      REGISTERS_18_13_port, REGISTERS_18_12_port, REGISTERS_18_11_port, 
      REGISTERS_18_10_port, REGISTERS_18_9_port, REGISTERS_18_8_port, 
      REGISTERS_18_7_port, REGISTERS_18_6_port, REGISTERS_18_5_port, 
      REGISTERS_18_4_port, REGISTERS_18_3_port, REGISTERS_18_2_port, 
      REGISTERS_18_1_port, REGISTERS_18_0_port, REGISTERS_19_31_port, 
      REGISTERS_19_30_port, REGISTERS_19_29_port, REGISTERS_19_28_port, 
      REGISTERS_19_27_port, REGISTERS_19_26_port, REGISTERS_19_25_port, 
      REGISTERS_19_24_port, REGISTERS_19_23_port, REGISTERS_19_22_port, 
      REGISTERS_19_21_port, REGISTERS_19_20_port, REGISTERS_19_19_port, 
      REGISTERS_19_18_port, REGISTERS_19_17_port, REGISTERS_19_16_port, 
      REGISTERS_19_15_port, REGISTERS_19_14_port, REGISTERS_19_13_port, 
      REGISTERS_19_12_port, REGISTERS_19_11_port, REGISTERS_19_10_port, 
      REGISTERS_19_9_port, REGISTERS_19_8_port, REGISTERS_19_7_port, 
      REGISTERS_19_6_port, REGISTERS_19_5_port, REGISTERS_19_4_port, 
      REGISTERS_19_3_port, REGISTERS_19_2_port, REGISTERS_19_1_port, 
      REGISTERS_19_0_port, REGISTERS_20_31_port, REGISTERS_20_30_port, 
      REGISTERS_20_29_port, REGISTERS_20_28_port, REGISTERS_20_27_port, 
      REGISTERS_20_26_port, REGISTERS_20_25_port, REGISTERS_20_24_port, 
      REGISTERS_20_23_port, REGISTERS_20_22_port, REGISTERS_20_21_port, 
      REGISTERS_20_20_port, REGISTERS_20_19_port, REGISTERS_20_18_port, 
      REGISTERS_20_17_port, REGISTERS_20_16_port, REGISTERS_20_15_port, 
      REGISTERS_20_14_port, REGISTERS_20_13_port, REGISTERS_20_12_port, 
      REGISTERS_20_11_port, REGISTERS_20_10_port, REGISTERS_20_9_port, 
      REGISTERS_20_8_port, REGISTERS_20_7_port, REGISTERS_20_6_port, 
      REGISTERS_20_5_port, REGISTERS_20_4_port, REGISTERS_20_3_port, 
      REGISTERS_20_2_port, REGISTERS_20_1_port, REGISTERS_20_0_port, 
      REGISTERS_21_31_port, REGISTERS_21_30_port, REGISTERS_21_29_port, 
      REGISTERS_21_28_port, REGISTERS_21_27_port, REGISTERS_21_26_port, 
      REGISTERS_21_25_port, REGISTERS_21_24_port, REGISTERS_21_23_port, 
      REGISTERS_21_22_port, REGISTERS_21_21_port, REGISTERS_21_20_port, 
      REGISTERS_21_19_port, REGISTERS_21_18_port, REGISTERS_21_17_port, 
      REGISTERS_21_16_port, REGISTERS_21_15_port, REGISTERS_21_14_port, 
      REGISTERS_21_13_port, REGISTERS_21_12_port, REGISTERS_21_11_port, 
      REGISTERS_21_10_port, REGISTERS_21_9_port, REGISTERS_21_8_port, 
      REGISTERS_21_7_port, REGISTERS_21_6_port, REGISTERS_21_5_port, 
      REGISTERS_21_4_port, REGISTERS_21_3_port, REGISTERS_21_2_port, 
      REGISTERS_21_1_port, REGISTERS_21_0_port, REGISTERS_22_31_port, 
      REGISTERS_22_30_port, REGISTERS_22_29_port, REGISTERS_22_28_port, 
      REGISTERS_22_27_port, REGISTERS_22_26_port, REGISTERS_22_25_port, 
      REGISTERS_22_24_port, REGISTERS_22_23_port, REGISTERS_22_22_port, 
      REGISTERS_22_21_port, REGISTERS_22_20_port, REGISTERS_22_19_port, 
      REGISTERS_22_18_port, REGISTERS_22_17_port, REGISTERS_22_16_port, 
      REGISTERS_22_15_port, REGISTERS_22_14_port, REGISTERS_22_13_port, 
      REGISTERS_22_12_port, REGISTERS_22_11_port, REGISTERS_22_10_port, 
      REGISTERS_22_9_port, REGISTERS_22_8_port, REGISTERS_22_7_port, 
      REGISTERS_22_6_port, REGISTERS_22_5_port, REGISTERS_22_4_port, 
      REGISTERS_22_3_port, REGISTERS_22_2_port, REGISTERS_22_1_port, 
      REGISTERS_22_0_port, REGISTERS_23_31_port, REGISTERS_23_30_port, 
      REGISTERS_23_29_port, REGISTERS_23_28_port, REGISTERS_23_27_port, 
      REGISTERS_23_26_port, REGISTERS_23_25_port, REGISTERS_23_24_port, 
      REGISTERS_23_23_port, REGISTERS_23_22_port, REGISTERS_23_21_port, 
      REGISTERS_23_20_port, REGISTERS_23_19_port, REGISTERS_23_18_port, 
      REGISTERS_23_17_port, REGISTERS_23_16_port, REGISTERS_23_15_port, 
      REGISTERS_23_14_port, REGISTERS_23_13_port, REGISTERS_23_12_port, 
      REGISTERS_23_11_port, REGISTERS_23_10_port, REGISTERS_23_9_port, 
      REGISTERS_23_8_port, REGISTERS_23_7_port, REGISTERS_23_6_port, 
      REGISTERS_23_5_port, REGISTERS_23_4_port, REGISTERS_23_3_port, 
      REGISTERS_23_2_port, REGISTERS_23_1_port, REGISTERS_23_0_port, 
      REGISTERS_24_31_port, REGISTERS_24_30_port, REGISTERS_24_29_port, 
      REGISTERS_24_28_port, REGISTERS_24_27_port, REGISTERS_24_26_port, 
      REGISTERS_24_25_port, REGISTERS_24_24_port, REGISTERS_24_23_port, 
      REGISTERS_24_22_port, REGISTERS_24_21_port, REGISTERS_24_20_port, 
      REGISTERS_24_19_port, REGISTERS_24_18_port, REGISTERS_24_17_port, 
      REGISTERS_24_16_port, REGISTERS_24_15_port, REGISTERS_24_14_port, 
      REGISTERS_24_13_port, REGISTERS_24_12_port, REGISTERS_24_11_port, 
      REGISTERS_24_10_port, REGISTERS_24_9_port, REGISTERS_24_8_port, 
      REGISTERS_24_7_port, REGISTERS_24_6_port, REGISTERS_24_5_port, 
      REGISTERS_24_4_port, REGISTERS_24_3_port, REGISTERS_24_2_port, 
      REGISTERS_24_1_port, REGISTERS_24_0_port, REGISTERS_25_31_port, 
      REGISTERS_25_30_port, REGISTERS_25_29_port, REGISTERS_25_28_port, 
      REGISTERS_25_27_port, REGISTERS_25_26_port, REGISTERS_25_25_port, 
      REGISTERS_25_24_port, REGISTERS_25_23_port, REGISTERS_25_22_port, 
      REGISTERS_25_21_port, REGISTERS_25_20_port, REGISTERS_25_19_port, 
      REGISTERS_25_18_port, REGISTERS_25_17_port, REGISTERS_25_16_port, 
      REGISTERS_25_15_port, REGISTERS_25_14_port, REGISTERS_25_13_port, 
      REGISTERS_25_12_port, REGISTERS_25_11_port, REGISTERS_25_10_port, 
      REGISTERS_25_9_port, REGISTERS_25_8_port, REGISTERS_25_7_port, 
      REGISTERS_25_6_port, REGISTERS_25_5_port, REGISTERS_25_4_port, 
      REGISTERS_25_3_port, REGISTERS_25_2_port, REGISTERS_25_1_port, 
      REGISTERS_25_0_port, REGISTERS_26_31_port, REGISTERS_26_30_port, 
      REGISTERS_26_29_port, REGISTERS_26_28_port, REGISTERS_26_27_port, 
      REGISTERS_26_26_port, REGISTERS_26_25_port, REGISTERS_26_24_port, 
      REGISTERS_26_23_port, REGISTERS_26_22_port, REGISTERS_26_21_port, 
      REGISTERS_26_20_port, REGISTERS_26_19_port, REGISTERS_26_18_port, 
      REGISTERS_26_17_port, REGISTERS_26_16_port, REGISTERS_26_15_port, 
      REGISTERS_26_14_port, REGISTERS_26_13_port, REGISTERS_26_12_port, 
      REGISTERS_26_11_port, REGISTERS_26_10_port, REGISTERS_26_9_port, 
      REGISTERS_26_8_port, REGISTERS_26_7_port, REGISTERS_26_6_port, 
      REGISTERS_26_5_port, REGISTERS_26_4_port, REGISTERS_26_3_port, 
      REGISTERS_26_2_port, REGISTERS_26_1_port, REGISTERS_26_0_port, 
      REGISTERS_27_31_port, REGISTERS_27_30_port, REGISTERS_27_29_port, 
      REGISTERS_27_28_port, REGISTERS_27_27_port, REGISTERS_27_26_port, 
      REGISTERS_27_25_port, REGISTERS_27_24_port, REGISTERS_27_23_port, 
      REGISTERS_27_22_port, REGISTERS_27_21_port, REGISTERS_27_20_port, 
      REGISTERS_27_19_port, REGISTERS_27_18_port, REGISTERS_27_17_port, 
      REGISTERS_27_16_port, REGISTERS_27_15_port, REGISTERS_27_14_port, 
      REGISTERS_27_13_port, REGISTERS_27_12_port, REGISTERS_27_11_port, 
      REGISTERS_27_10_port, REGISTERS_27_9_port, REGISTERS_27_8_port, 
      REGISTERS_27_7_port, REGISTERS_27_6_port, REGISTERS_27_5_port, 
      REGISTERS_27_4_port, REGISTERS_27_3_port, REGISTERS_27_2_port, 
      REGISTERS_27_1_port, REGISTERS_27_0_port, REGISTERS_28_31_port, 
      REGISTERS_28_30_port, REGISTERS_28_29_port, REGISTERS_28_28_port, 
      REGISTERS_28_27_port, REGISTERS_28_26_port, REGISTERS_28_25_port, 
      REGISTERS_28_24_port, REGISTERS_28_23_port, REGISTERS_28_22_port, 
      REGISTERS_28_21_port, REGISTERS_28_20_port, REGISTERS_28_19_port, 
      REGISTERS_28_18_port, REGISTERS_28_17_port, REGISTERS_28_16_port, 
      REGISTERS_28_15_port, REGISTERS_28_14_port, REGISTERS_28_13_port, 
      REGISTERS_28_12_port, REGISTERS_28_11_port, REGISTERS_28_10_port, 
      REGISTERS_28_9_port, REGISTERS_28_8_port, REGISTERS_28_7_port, 
      REGISTERS_28_6_port, REGISTERS_28_5_port, REGISTERS_28_4_port, 
      REGISTERS_28_3_port, REGISTERS_28_2_port, REGISTERS_28_1_port, 
      REGISTERS_28_0_port, REGISTERS_29_31_port, REGISTERS_29_30_port, 
      REGISTERS_29_29_port, REGISTERS_29_28_port, REGISTERS_29_27_port, 
      REGISTERS_29_26_port, REGISTERS_29_25_port, REGISTERS_29_24_port, 
      REGISTERS_29_23_port, REGISTERS_29_22_port, REGISTERS_29_21_port, 
      REGISTERS_29_20_port, REGISTERS_29_19_port, REGISTERS_29_18_port, 
      REGISTERS_29_17_port, REGISTERS_29_16_port, REGISTERS_29_15_port, 
      REGISTERS_29_14_port, REGISTERS_29_13_port, REGISTERS_29_12_port, 
      REGISTERS_29_11_port, REGISTERS_29_10_port, REGISTERS_29_9_port, 
      REGISTERS_29_8_port, REGISTERS_29_7_port, REGISTERS_29_6_port, 
      REGISTERS_29_5_port, REGISTERS_29_4_port, REGISTERS_29_3_port, 
      REGISTERS_29_2_port, REGISTERS_29_1_port, REGISTERS_29_0_port, 
      REGISTERS_30_31_port, REGISTERS_30_30_port, REGISTERS_30_29_port, 
      REGISTERS_30_28_port, REGISTERS_30_27_port, REGISTERS_30_26_port, 
      REGISTERS_30_25_port, REGISTERS_30_24_port, REGISTERS_30_23_port, 
      REGISTERS_30_22_port, REGISTERS_30_21_port, REGISTERS_30_20_port, 
      REGISTERS_30_19_port, REGISTERS_30_18_port, REGISTERS_30_17_port, 
      REGISTERS_30_16_port, REGISTERS_30_15_port, REGISTERS_30_14_port, 
      REGISTERS_30_13_port, REGISTERS_30_12_port, REGISTERS_30_11_port, 
      REGISTERS_30_10_port, REGISTERS_30_9_port, REGISTERS_30_8_port, 
      REGISTERS_30_7_port, REGISTERS_30_6_port, REGISTERS_30_5_port, 
      REGISTERS_30_4_port, REGISTERS_30_3_port, REGISTERS_30_2_port, 
      REGISTERS_30_1_port, REGISTERS_30_0_port, REGISTERS_31_31_port, 
      REGISTERS_31_30_port, REGISTERS_31_29_port, REGISTERS_31_28_port, 
      REGISTERS_31_27_port, REGISTERS_31_26_port, REGISTERS_31_25_port, 
      REGISTERS_31_24_port, REGISTERS_31_23_port, REGISTERS_31_22_port, 
      REGISTERS_31_21_port, REGISTERS_31_20_port, REGISTERS_31_19_port, 
      REGISTERS_31_18_port, REGISTERS_31_17_port, REGISTERS_31_16_port, 
      REGISTERS_31_15_port, REGISTERS_31_14_port, REGISTERS_31_13_port, 
      REGISTERS_31_12_port, REGISTERS_31_11_port, REGISTERS_31_10_port, 
      REGISTERS_31_9_port, REGISTERS_31_8_port, REGISTERS_31_7_port, 
      REGISTERS_31_6_port, REGISTERS_31_5_port, REGISTERS_31_4_port, 
      REGISTERS_31_3_port, REGISTERS_31_2_port, REGISTERS_31_1_port, 
      REGISTERS_31_0_port, N156, N157, N158, N159, N160, N161, N162, N163, N164
      , N165, N166, N167, N168, N169, N170, N171, N172, N173, N174, N175, N176,
      N177, N178, N179, N180, N181, N182, N183, N184, N185, N186, N187, N189, 
      N190, N191, N192, N193, N194, N195, N196, N197, N198, N199, N200, N201, 
      N202, N203, N204, N205, N206, N207, N208, N209, N210, N211, N212, N213, 
      N214, N215, N216, N217, N218, N219, N220, n1399, n1401, n1403, n1405, 
      n1407, n1409, n1411, n1413, n1415, n1417, n1419, n1421, n1423, n1425, 
      n1427, n1429, n1431, n1433, n1435, n1437, n1439, n1441, n1443, n1445, 
      n1447, n1449, n1451, n1453, n1455, n1457, n1459, n1461, n1463, n1464, 
      n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, 
      n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, 
      n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, 
      n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, 
      n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, 
      n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, 
      n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, 
      n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, 
      n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, 
      n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, 
      n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, 
      n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, 
      n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, 
      n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, 
      n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, 
      n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, 
      n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, 
      n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, 
      n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, 
      n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, 
      n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, 
      n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, 
      n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, 
      n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, 
      n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, 
      n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, 
      n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, 
      n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, 
      n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, 
      n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, 
      n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, 
      n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, 
      n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, 
      n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, 
      n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, 
      n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, 
      n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, 
      n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, 
      n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, 
      n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, 
      n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, 
      n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, 
      n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, 
      n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, 
      n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, 
      n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, 
      n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, 
      n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, 
      n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, 
      n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, 
      n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, 
      n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, 
      n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, 
      n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, 
      n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, 
      n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, 
      n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, 
      n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, 
      n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, 
      n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, 
      n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, 
      n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, 
      n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, 
      n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, 
      n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, 
      n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, 
      n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, 
      n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, 
      n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, 
      n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, 
      n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, 
      n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, 
      n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, 
      n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, 
      n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, 
      n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, 
      n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, 
      n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, 
      n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, 
      n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, 
      n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, 
      n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, 
      n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, 
      n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, 
      n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, 
      n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, 
      n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, 
      n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, 
      n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, 
      n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, 
      n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, 
      n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, 
      n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, 
      n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, 
      n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, 
      n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, 
      n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, 
      n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, 
      n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, 
      n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, 
      n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, 
      n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, 
      n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, 
      n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, 
      n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, 
      n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, 
      n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, 
      n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, 
      n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, 
      n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, 
      n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, 
      n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n1, n2, n3, n4, 
      n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20
      , n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, 
      n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49
      , n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, 
      n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78
      , n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, 
      n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, 
      n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, 
      n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, 
      n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, 
      n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, 
      n154, n155, n156_port, n157_port, n158_port, n159_port, n160_port, 
      n161_port, n162_port, n163_port, n164_port, n165_port, n166_port, 
      n167_port, n168_port, n169_port, n170_port, n171_port, n172_port, 
      n173_port, n174_port, n175_port, n176_port, n177_port, n178_port, 
      n179_port, n180_port, n181_port, n182_port, n183_port, n184_port, 
      n185_port, n186_port, n187_port, n188, n189_port, n190_port, n191_port, 
      n192_port, n193_port, n194_port, n195_port, n196_port, n197_port, 
      n198_port, n199_port, n200_port, n201_port, n202_port, n203_port, 
      n204_port, n205_port, n206_port, n207_port, n208_port, n209_port, 
      n210_port, n211_port, n212_port, n213_port, n214_port, n215_port, 
      n216_port, n217_port, n218_port, n219_port, n220_port, n221, n222, n223, 
      n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, 
      n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, 
      n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, 
      n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, 
      n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, 
      n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, 
      n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, 
      n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, 
      n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, 
      n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, 
      n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, 
      n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, 
      n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, 
      n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, 
      n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, 
      n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, 
      n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, 
      n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, 
      n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, 
      n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, 
      n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, 
      n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, 
      n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, 
      n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, 
      n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, 
      n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, 
      n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, 
      n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, 
      n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, 
      n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, 
      n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, 
      n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, 
      n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, 
      n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, 
      n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, 
      n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, 
      n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, 
      n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, 
      n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, 
      n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, 
      n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, 
      n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, 
      n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, 
      n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, 
      n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, 
      n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, 
      n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, 
      n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, 
      n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, 
      n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, 
      n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, 
      n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, 
      n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, 
      n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, 
      n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, 
      n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, 
      n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, 
      n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, 
      n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, 
      n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, 
      n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, 
      n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, 
      n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, 
      n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, 
      n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, 
      n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, 
      n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, 
      n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, 
      n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, 
      n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, 
      n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, 
      n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, 
      n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, 
      n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, 
      n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, 
      n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, 
      n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, 
      n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, 
      n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, 
      n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, 
      n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, 
      n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, 
      n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, 
      n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, 
      n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, 
      n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, 
      n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, 
      n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, 
      n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, 
      n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, 
      n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, 
      n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, 
      n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, 
      n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, 
      n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, 
      n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, 
      n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, 
      n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, 
      n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, 
      n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, 
      n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, 
      n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, 
      n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, 
      n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, 
      n1393, n1394, n1395, n1396, n1397, n1398, n1400, n1402, n1404, n1406, 
      n1408, n1410, n1412, n1414, n1416, n1418, n1420, n1422, n1424, n1426, 
      n1428, n1430, n1432, n1434, n1436, n1438, n1440, n1442, n1444, n1446, 
      n1448, n1450, n1452, n1454, n1456, n1458, n1460, n1462, n1495, n1496, 
      n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, 
      n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, 
      n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, 
      n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, 
      n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, 
      n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, 
      n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, 
      n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, 
      n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, 
      n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, 
      n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, 
      n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, 
      n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, 
      n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, 
      n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, 
      n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, 
      n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, 
      n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, 
      n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, 
      n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, 
      n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, 
      n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, 
      n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, 
      n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, 
      n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, 
      n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, 
      n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, 
      n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, 
      n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, 
      n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, 
      n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, 
      n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, 
      n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, 
      n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, 
      n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, 
      n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, 
      n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, 
      n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, 
      n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, 
      n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, 
      n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, 
      n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, 
      n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, 
      n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, 
      n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, 
      n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, 
      n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, 
      n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, 
      n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, 
      n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, 
      n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, 
      n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, 
      n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, 
      n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, 
      n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, 
      n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, 
      n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, 
      n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, 
      n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, 
      n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, 
      n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, 
      n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, 
      n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, 
      n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, 
      n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, 
      n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, 
      n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, 
      n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, 
      n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, 
      n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, 
      n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, 
      n3295, n3296, n3297, n3298, n3299, n3300, n_1000, n_1001, n_1002, n_1003,
      n_1004, n_1005, n_1006, n_1007, n_1008, n_1009, n_1010, n_1011, n_1012, 
      n_1013, n_1014, n_1015, n_1016, n_1017, n_1018, n_1019, n_1020, n_1021, 
      n_1022, n_1023, n_1024, n_1025, n_1026, n_1027, n_1028, n_1029, n_1030, 
      n_1031, n_1032, n_1033, n_1034, n_1035, n_1036, n_1037, n_1038, n_1039, 
      n_1040, n_1041, n_1042, n_1043, n_1044, n_1045, n_1046, n_1047, n_1048, 
      n_1049, n_1050, n_1051, n_1052, n_1053, n_1054, n_1055, n_1056, n_1057, 
      n_1058, n_1059, n_1060, n_1061, n_1062, n_1063, n_1064, n_1065, n_1066, 
      n_1067, n_1068, n_1069, n_1070, n_1071, n_1072, n_1073, n_1074, n_1075, 
      n_1076, n_1077, n_1078, n_1079, n_1080, n_1081, n_1082, n_1083, n_1084, 
      n_1085, n_1086, n_1087, n_1088, n_1089, n_1090, n_1091, n_1092, n_1093, 
      n_1094, n_1095, n_1096, n_1097, n_1098, n_1099, n_1100, n_1101, n_1102, 
      n_1103, n_1104, n_1105, n_1106, n_1107, n_1108, n_1109, n_1110, n_1111, 
      n_1112, n_1113, n_1114, n_1115, n_1116, n_1117, n_1118, n_1119, n_1120, 
      n_1121, n_1122, n_1123, n_1124, n_1125, n_1126, n_1127, n_1128, n_1129, 
      n_1130, n_1131, n_1132, n_1133, n_1134, n_1135, n_1136, n_1137, n_1138, 
      n_1139, n_1140, n_1141, n_1142, n_1143, n_1144, n_1145, n_1146, n_1147, 
      n_1148, n_1149, n_1150, n_1151, n_1152, n_1153, n_1154, n_1155, n_1156, 
      n_1157, n_1158, n_1159, n_1160, n_1161, n_1162, n_1163, n_1164, n_1165, 
      n_1166, n_1167, n_1168, n_1169, n_1170, n_1171, n_1172, n_1173, n_1174, 
      n_1175, n_1176, n_1177, n_1178, n_1179, n_1180, n_1181, n_1182, n_1183, 
      n_1184, n_1185, n_1186, n_1187, n_1188, n_1189, n_1190, n_1191, n_1192, 
      n_1193, n_1194, n_1195, n_1196, n_1197, n_1198, n_1199, n_1200, n_1201, 
      n_1202, n_1203, n_1204, n_1205, n_1206, n_1207, n_1208, n_1209, n_1210, 
      n_1211, n_1212, n_1213, n_1214, n_1215, n_1216, n_1217, n_1218, n_1219, 
      n_1220, n_1221, n_1222, n_1223, n_1224, n_1225, n_1226, n_1227, n_1228, 
      n_1229, n_1230, n_1231, n_1232, n_1233, n_1234, n_1235, n_1236, n_1237, 
      n_1238, n_1239, n_1240, n_1241, n_1242, n_1243, n_1244, n_1245, n_1246, 
      n_1247, n_1248, n_1249, n_1250, n_1251, n_1252, n_1253, n_1254, n_1255, 
      n_1256, n_1257, n_1258, n_1259, n_1260, n_1261, n_1262, n_1263, n_1264, 
      n_1265, n_1266, n_1267, n_1268, n_1269, n_1270, n_1271, n_1272, n_1273, 
      n_1274, n_1275, n_1276, n_1277, n_1278, n_1279, n_1280, n_1281, n_1282, 
      n_1283, n_1284, n_1285, n_1286, n_1287, n_1288, n_1289, n_1290, n_1291, 
      n_1292, n_1293, n_1294, n_1295, n_1296, n_1297, n_1298, n_1299, n_1300, 
      n_1301, n_1302, n_1303, n_1304, n_1305, n_1306, n_1307, n_1308, n_1309, 
      n_1310, n_1311, n_1312, n_1313, n_1314, n_1315, n_1316, n_1317, n_1318, 
      n_1319, n_1320, n_1321, n_1322, n_1323, n_1324, n_1325, n_1326, n_1327, 
      n_1328, n_1329, n_1330, n_1331, n_1332, n_1333, n_1334, n_1335, n_1336, 
      n_1337, n_1338, n_1339, n_1340, n_1341, n_1342, n_1343, n_1344, n_1345, 
      n_1346, n_1347, n_1348, n_1349, n_1350, n_1351, n_1352, n_1353, n_1354, 
      n_1355, n_1356, n_1357, n_1358, n_1359, n_1360, n_1361, n_1362, n_1363, 
      n_1364, n_1365, n_1366, n_1367, n_1368, n_1369, n_1370, n_1371, n_1372, 
      n_1373, n_1374, n_1375, n_1376, n_1377, n_1378, n_1379, n_1380, n_1381, 
      n_1382, n_1383, n_1384, n_1385, n_1386, n_1387, n_1388, n_1389, n_1390, 
      n_1391, n_1392, n_1393, n_1394, n_1395, n_1396, n_1397, n_1398, n_1399, 
      n_1400, n_1401, n_1402, n_1403, n_1404, n_1405, n_1406, n_1407, n_1408, 
      n_1409, n_1410, n_1411, n_1412, n_1413, n_1414, n_1415, n_1416, n_1417, 
      n_1418, n_1419, n_1420, n_1421, n_1422, n_1423, n_1424, n_1425, n_1426, 
      n_1427, n_1428, n_1429, n_1430, n_1431, n_1432, n_1433, n_1434, n_1435, 
      n_1436, n_1437, n_1438, n_1439, n_1440, n_1441, n_1442, n_1443, n_1444, 
      n_1445, n_1446, n_1447, n_1448, n_1449, n_1450, n_1451, n_1452, n_1453, 
      n_1454, n_1455, n_1456, n_1457, n_1458, n_1459, n_1460, n_1461, n_1462, 
      n_1463, n_1464, n_1465, n_1466, n_1467, n_1468, n_1469, n_1470, n_1471, 
      n_1472, n_1473, n_1474, n_1475, n_1476, n_1477, n_1478, n_1479, n_1480, 
      n_1481, n_1482, n_1483, n_1484, n_1485, n_1486, n_1487, n_1488, n_1489, 
      n_1490, n_1491, n_1492, n_1493, n_1494, n_1495, n_1496, n_1497, n_1498, 
      n_1499, n_1500, n_1501, n_1502, n_1503, n_1504, n_1505, n_1506, n_1507, 
      n_1508, n_1509, n_1510, n_1511, n_1512, n_1513, n_1514, n_1515, n_1516, 
      n_1517, n_1518, n_1519, n_1520, n_1521, n_1522, n_1523, n_1524, n_1525, 
      n_1526, n_1527, n_1528, n_1529, n_1530, n_1531, n_1532, n_1533, n_1534, 
      n_1535, n_1536, n_1537, n_1538, n_1539, n_1540, n_1541, n_1542, n_1543, 
      n_1544, n_1545, n_1546, n_1547, n_1548, n_1549, n_1550, n_1551, n_1552, 
      n_1553, n_1554, n_1555, n_1556, n_1557, n_1558, n_1559, n_1560, n_1561, 
      n_1562, n_1563, n_1564, n_1565, n_1566, n_1567, n_1568, n_1569, n_1570, 
      n_1571, n_1572, n_1573, n_1574, n_1575, n_1576, n_1577, n_1578, n_1579, 
      n_1580, n_1581, n_1582, n_1583, n_1584, n_1585, n_1586, n_1587, n_1588, 
      n_1589, n_1590, n_1591, n_1592, n_1593, n_1594, n_1595, n_1596, n_1597, 
      n_1598, n_1599, n_1600, n_1601, n_1602, n_1603, n_1604, n_1605, n_1606, 
      n_1607, n_1608, n_1609, n_1610, n_1611, n_1612, n_1613, n_1614, n_1615, 
      n_1616, n_1617, n_1618, n_1619, n_1620, n_1621, n_1622, n_1623, n_1624, 
      n_1625, n_1626, n_1627, n_1628, n_1629, n_1630, n_1631, n_1632, n_1633, 
      n_1634, n_1635, n_1636, n_1637, n_1638, n_1639, n_1640, n_1641, n_1642, 
      n_1643, n_1644, n_1645, n_1646, n_1647, n_1648, n_1649, n_1650, n_1651, 
      n_1652, n_1653, n_1654, n_1655, n_1656, n_1657, n_1658, n_1659, n_1660, 
      n_1661, n_1662, n_1663, n_1664, n_1665, n_1666, n_1667, n_1668, n_1669, 
      n_1670, n_1671, n_1672, n_1673, n_1674, n_1675, n_1676, n_1677, n_1678, 
      n_1679, n_1680, n_1681, n_1682, n_1683, n_1684, n_1685, n_1686, n_1687, 
      n_1688, n_1689, n_1690, n_1691, n_1692, n_1693, n_1694, n_1695, n_1696, 
      n_1697, n_1698, n_1699, n_1700, n_1701, n_1702, n_1703, n_1704, n_1705, 
      n_1706, n_1707, n_1708, n_1709, n_1710, n_1711, n_1712, n_1713, n_1714, 
      n_1715, n_1716, n_1717, n_1718, n_1719, n_1720, n_1721, n_1722, n_1723, 
      n_1724, n_1725, n_1726, n_1727, n_1728, n_1729, n_1730, n_1731, n_1732, 
      n_1733, n_1734, n_1735, n_1736, n_1737, n_1738, n_1739, n_1740, n_1741, 
      n_1742, n_1743, n_1744, n_1745, n_1746, n_1747, n_1748, n_1749, n_1750, 
      n_1751, n_1752, n_1753, n_1754, n_1755, n_1756, n_1757, n_1758, n_1759, 
      n_1760, n_1761, n_1762, n_1763, n_1764, n_1765, n_1766, n_1767, n_1768, 
      n_1769, n_1770, n_1771, n_1772, n_1773, n_1774, n_1775, n_1776, n_1777, 
      n_1778, n_1779, n_1780, n_1781, n_1782, n_1783, n_1784, n_1785, n_1786, 
      n_1787, n_1788, n_1789, n_1790, n_1791, n_1792, n_1793, n_1794, n_1795, 
      n_1796, n_1797, n_1798, n_1799, n_1800, n_1801, n_1802, n_1803, n_1804, 
      n_1805, n_1806, n_1807, n_1808, n_1809, n_1810, n_1811, n_1812, n_1813, 
      n_1814, n_1815, n_1816, n_1817, n_1818, n_1819, n_1820, n_1821, n_1822, 
      n_1823, n_1824, n_1825, n_1826, n_1827, n_1828, n_1829, n_1830, n_1831, 
      n_1832, n_1833, n_1834, n_1835, n_1836, n_1837, n_1838, n_1839, n_1840, 
      n_1841, n_1842, n_1843, n_1844, n_1845, n_1846, n_1847, n_1848, n_1849, 
      n_1850, n_1851, n_1852, n_1853, n_1854, n_1855, n_1856, n_1857, n_1858, 
      n_1859, n_1860, n_1861, n_1862, n_1863, n_1864, n_1865, n_1866, n_1867, 
      n_1868, n_1869, n_1870, n_1871, n_1872, n_1873, n_1874, n_1875, n_1876, 
      n_1877, n_1878, n_1879, n_1880, n_1881, n_1882, n_1883, n_1884, n_1885, 
      n_1886, n_1887, n_1888, n_1889, n_1890, n_1891, n_1892, n_1893, n_1894, 
      n_1895, n_1896, n_1897, n_1898, n_1899, n_1900, n_1901, n_1902, n_1903, 
      n_1904, n_1905, n_1906, n_1907, n_1908, n_1909, n_1910, n_1911, n_1912, 
      n_1913, n_1914, n_1915, n_1916, n_1917, n_1918, n_1919, n_1920, n_1921, 
      n_1922, n_1923, n_1924, n_1925, n_1926, n_1927, n_1928, n_1929, n_1930, 
      n_1931, n_1932, n_1933, n_1934, n_1935, n_1936, n_1937, n_1938, n_1939, 
      n_1940, n_1941, n_1942, n_1943, n_1944, n_1945, n_1946, n_1947, n_1948, 
      n_1949, n_1950, n_1951, n_1952, n_1953, n_1954, n_1955, n_1956, n_1957, 
      n_1958, n_1959, n_1960, n_1961, n_1962, n_1963, n_1964, n_1965, n_1966, 
      n_1967, n_1968, n_1969, n_1970, n_1971, n_1972, n_1973, n_1974, n_1975, 
      n_1976, n_1977, n_1978, n_1979, n_1980, n_1981, n_1982, n_1983, n_1984, 
      n_1985, n_1986, n_1987, n_1988, n_1989, n_1990, n_1991, n_1992, n_1993, 
      n_1994, n_1995, n_1996, n_1997, n_1998, n_1999, n_2000, n_2001, n_2002, 
      n_2003, n_2004, n_2005, n_2006, n_2007, n_2008, n_2009, n_2010, n_2011, 
      n_2012, n_2013, n_2014, n_2015, n_2016, n_2017, n_2018, n_2019, n_2020, 
      n_2021, n_2022, n_2023, n_2024, n_2025, n_2026, n_2027, n_2028, n_2029, 
      n_2030, n_2031, n_2032, n_2033, n_2034, n_2035, n_2036, n_2037, n_2038, 
      n_2039, n_2040, n_2041, n_2042, n_2043, n_2044, n_2045, n_2046, n_2047, 
      n_2048, n_2049, n_2050, n_2051, n_2052, n_2053, n_2054, n_2055, n_2056, 
      n_2057, n_2058, n_2059, n_2060, n_2061, n_2062, n_2063, n_2064, n_2065, 
      n_2066, n_2067, n_2068, n_2069, n_2070, n_2071, n_2072, n_2073, n_2074, 
      n_2075, n_2076, n_2077, n_2078, n_2079, n_2080, n_2081, n_2082, n_2083, 
      n_2084, n_2085, n_2086, n_2087 : std_logic;

begin
   
   OUT1_reg_31_inst : DFF_X1 port map( D => n1399, CK => n415, Q => n3173, QN 
                           => n_1000);
   OUT1_tri_enable_reg_31_inst : DFF_X1 port map( D => n2614, CK => n513, Q => 
                           n3174, QN => n17);
   OUT1_reg_30_inst : DFF_X1 port map( D => n1401, CK => n415, Q => n3175, QN 
                           => n_1001);
   OUT1_tri_enable_reg_30_inst : DFF_X1 port map( D => n2613, CK => n514, Q => 
                           n3176, QN => n18);
   OUT1_reg_29_inst : DFF_X1 port map( D => n1403, CK => n415, Q => n3177, QN 
                           => n_1002);
   OUT1_tri_enable_reg_29_inst : DFF_X1 port map( D => n2612, CK => n514, Q => 
                           n3178, QN => n19);
   OUT1_reg_28_inst : DFF_X1 port map( D => n1405, CK => n415, Q => n3179, QN 
                           => n_1003);
   OUT1_tri_enable_reg_28_inst : DFF_X1 port map( D => n2611, CK => n514, Q => 
                           n3180, QN => n20);
   OUT1_reg_27_inst : DFF_X1 port map( D => n1407, CK => n415, Q => n3181, QN 
                           => n_1004);
   OUT1_tri_enable_reg_27_inst : DFF_X1 port map( D => n2610, CK => n514, Q => 
                           n3182, QN => n21);
   OUT1_reg_26_inst : DFF_X1 port map( D => n1409, CK => n415, Q => n3183, QN 
                           => n_1005);
   OUT1_tri_enable_reg_26_inst : DFF_X1 port map( D => n2609, CK => n514, Q => 
                           n3184, QN => n22);
   OUT1_reg_25_inst : DFF_X1 port map( D => n1411, CK => n415, Q => n3185, QN 
                           => n_1006);
   OUT1_tri_enable_reg_25_inst : DFF_X1 port map( D => n2608, CK => n514, Q => 
                           n3186, QN => n23);
   OUT1_reg_24_inst : DFF_X1 port map( D => n1413, CK => n415, Q => n3187, QN 
                           => n_1007);
   OUT1_tri_enable_reg_24_inst : DFF_X1 port map( D => n2607, CK => n514, Q => 
                           n3188, QN => n24);
   OUT1_reg_23_inst : DFF_X1 port map( D => n1415, CK => n415, Q => n3189, QN 
                           => n_1008);
   OUT1_tri_enable_reg_23_inst : DFF_X1 port map( D => n2606, CK => n514, Q => 
                           n3190, QN => n25);
   OUT1_reg_22_inst : DFF_X1 port map( D => n1417, CK => n415, Q => n3191, QN 
                           => n_1009);
   OUT1_tri_enable_reg_22_inst : DFF_X1 port map( D => n2605, CK => n514, Q => 
                           n3192, QN => n26);
   OUT1_reg_21_inst : DFF_X1 port map( D => n1419, CK => n415, Q => n3193, QN 
                           => n_1010);
   OUT1_tri_enable_reg_21_inst : DFF_X1 port map( D => n2604, CK => n514, Q => 
                           n3194, QN => n27);
   OUT1_reg_20_inst : DFF_X1 port map( D => n1421, CK => n416, Q => n3195, QN 
                           => n_1011);
   OUT1_tri_enable_reg_20_inst : DFF_X1 port map( D => n2603, CK => n514, Q => 
                           n3196, QN => n28);
   OUT1_reg_19_inst : DFF_X1 port map( D => n1423, CK => n416, Q => n3197, QN 
                           => n_1012);
   OUT1_tri_enable_reg_19_inst : DFF_X1 port map( D => n2602, CK => n515, Q => 
                           n3198, QN => n29);
   OUT1_reg_18_inst : DFF_X1 port map( D => n1425, CK => n416, Q => n3199, QN 
                           => n_1013);
   OUT1_tri_enable_reg_18_inst : DFF_X1 port map( D => n2601, CK => n515, Q => 
                           n3200, QN => n30);
   OUT1_reg_17_inst : DFF_X1 port map( D => n1427, CK => n416, Q => n3201, QN 
                           => n_1014);
   OUT1_tri_enable_reg_17_inst : DFF_X1 port map( D => n2600, CK => n515, Q => 
                           n3202, QN => n31);
   OUT1_reg_16_inst : DFF_X1 port map( D => n1429, CK => n416, Q => n3203, QN 
                           => n_1015);
   OUT1_tri_enable_reg_16_inst : DFF_X1 port map( D => n2599, CK => n515, Q => 
                           n3204, QN => n32);
   OUT1_reg_15_inst : DFF_X1 port map( D => n1431, CK => n416, Q => n3205, QN 
                           => n_1016);
   OUT1_tri_enable_reg_15_inst : DFF_X1 port map( D => n2598, CK => n515, Q => 
                           n3206, QN => n33);
   OUT1_reg_14_inst : DFF_X1 port map( D => n1433, CK => n416, Q => n3207, QN 
                           => n_1017);
   OUT1_tri_enable_reg_14_inst : DFF_X1 port map( D => n2597, CK => n515, Q => 
                           n3208, QN => n34);
   OUT1_reg_13_inst : DFF_X1 port map( D => n1435, CK => n416, Q => n3209, QN 
                           => n_1018);
   OUT1_tri_enable_reg_13_inst : DFF_X1 port map( D => n2596, CK => n515, Q => 
                           n3210, QN => n35);
   OUT1_reg_12_inst : DFF_X1 port map( D => n1437, CK => n416, Q => n3211, QN 
                           => n_1019);
   OUT1_tri_enable_reg_12_inst : DFF_X1 port map( D => n2595, CK => n515, Q => 
                           n3212, QN => n36);
   OUT1_reg_11_inst : DFF_X1 port map( D => n1439, CK => n416, Q => n3213, QN 
                           => n_1020);
   OUT1_tri_enable_reg_11_inst : DFF_X1 port map( D => n2594, CK => n515, Q => 
                           n3214, QN => n37);
   OUT1_reg_10_inst : DFF_X1 port map( D => n1441, CK => n416, Q => n3215, QN 
                           => n_1021);
   OUT1_tri_enable_reg_10_inst : DFF_X1 port map( D => n2593, CK => n515, Q => 
                           n3216, QN => n38);
   OUT1_reg_9_inst : DFF_X1 port map( D => n1443, CK => n417, Q => n3217, QN =>
                           n_1022);
   OUT1_tri_enable_reg_9_inst : DFF_X1 port map( D => n2592, CK => n515, Q => 
                           n3218, QN => n39);
   OUT1_reg_8_inst : DFF_X1 port map( D => n1445, CK => n417, Q => n3219, QN =>
                           n_1023);
   OUT1_tri_enable_reg_8_inst : DFF_X1 port map( D => n2591, CK => n516, Q => 
                           n3220, QN => n40);
   OUT1_reg_7_inst : DFF_X1 port map( D => n1447, CK => n417, Q => n3221, QN =>
                           n_1024);
   OUT1_tri_enable_reg_7_inst : DFF_X1 port map( D => n2590, CK => n516, Q => 
                           n3222, QN => n41);
   OUT1_reg_6_inst : DFF_X1 port map( D => n1449, CK => n417, Q => n3223, QN =>
                           n_1025);
   OUT1_tri_enable_reg_6_inst : DFF_X1 port map( D => n2589, CK => n516, Q => 
                           n3224, QN => n42);
   OUT1_reg_5_inst : DFF_X1 port map( D => n1451, CK => n417, Q => n3225, QN =>
                           n_1026);
   OUT1_tri_enable_reg_5_inst : DFF_X1 port map( D => n2588, CK => n516, Q => 
                           n3226, QN => n43);
   OUT1_reg_4_inst : DFF_X1 port map( D => n1453, CK => n417, Q => n3227, QN =>
                           n_1027);
   OUT1_tri_enable_reg_4_inst : DFF_X1 port map( D => n2587, CK => n516, Q => 
                           n3228, QN => n44);
   OUT1_reg_3_inst : DFF_X1 port map( D => n1455, CK => n417, Q => n3229, QN =>
                           n_1028);
   OUT1_tri_enable_reg_3_inst : DFF_X1 port map( D => n2586, CK => n516, Q => 
                           n3230, QN => n45);
   OUT1_reg_2_inst : DFF_X1 port map( D => n1457, CK => n417, Q => n3231, QN =>
                           n_1029);
   OUT1_tri_enable_reg_2_inst : DFF_X1 port map( D => n2585, CK => n516, Q => 
                           n3232, QN => n46);
   OUT1_reg_1_inst : DFF_X1 port map( D => n1459, CK => n417, Q => n3233, QN =>
                           n_1030);
   OUT1_tri_enable_reg_1_inst : DFF_X1 port map( D => n2584, CK => n516, Q => 
                           n3234, QN => n47);
   OUT1_reg_0_inst : DFF_X1 port map( D => n1461, CK => n417, Q => n3235, QN =>
                           n_1031);
   OUT1_tri_enable_reg_0_inst : DFF_X1 port map( D => n2583, CK => n516, Q => 
                           n3236, QN => n48);
   REGISTERS_reg_0_31_inst : DFF_X1 port map( D => n2582, CK => n467, Q => 
                           REGISTERS_0_31_port, QN => n_1032);
   REGISTERS_reg_0_30_inst : DFF_X1 port map( D => n2581, CK => n467, Q => 
                           REGISTERS_0_30_port, QN => n_1033);
   REGISTERS_reg_0_29_inst : DFF_X1 port map( D => n2580, CK => n467, Q => 
                           REGISTERS_0_29_port, QN => n_1034);
   REGISTERS_reg_0_28_inst : DFF_X1 port map( D => n2579, CK => n467, Q => 
                           REGISTERS_0_28_port, QN => n_1035);
   REGISTERS_reg_0_27_inst : DFF_X1 port map( D => n2578, CK => n467, Q => 
                           REGISTERS_0_27_port, QN => n_1036);
   REGISTERS_reg_0_26_inst : DFF_X1 port map( D => n2577, CK => n467, Q => 
                           REGISTERS_0_26_port, QN => n_1037);
   REGISTERS_reg_0_25_inst : DFF_X1 port map( D => n2576, CK => n467, Q => 
                           REGISTERS_0_25_port, QN => n_1038);
   REGISTERS_reg_0_24_inst : DFF_X1 port map( D => n2575, CK => n468, Q => 
                           REGISTERS_0_24_port, QN => n_1039);
   REGISTERS_reg_0_23_inst : DFF_X1 port map( D => n2574, CK => n468, Q => 
                           REGISTERS_0_23_port, QN => n_1040);
   REGISTERS_reg_0_22_inst : DFF_X1 port map( D => n2573, CK => n468, Q => 
                           REGISTERS_0_22_port, QN => n_1041);
   REGISTERS_reg_0_21_inst : DFF_X1 port map( D => n2572, CK => n468, Q => 
                           REGISTERS_0_21_port, QN => n_1042);
   REGISTERS_reg_0_20_inst : DFF_X1 port map( D => n2571, CK => n468, Q => 
                           REGISTERS_0_20_port, QN => n_1043);
   REGISTERS_reg_0_19_inst : DFF_X1 port map( D => n2570, CK => n468, Q => 
                           REGISTERS_0_19_port, QN => n_1044);
   REGISTERS_reg_0_18_inst : DFF_X1 port map( D => n2569, CK => n468, Q => 
                           REGISTERS_0_18_port, QN => n_1045);
   REGISTERS_reg_0_17_inst : DFF_X1 port map( D => n2568, CK => n468, Q => 
                           REGISTERS_0_17_port, QN => n_1046);
   REGISTERS_reg_0_16_inst : DFF_X1 port map( D => n2567, CK => n468, Q => 
                           REGISTERS_0_16_port, QN => n_1047);
   REGISTERS_reg_0_15_inst : DFF_X1 port map( D => n2566, CK => n468, Q => 
                           REGISTERS_0_15_port, QN => n_1048);
   REGISTERS_reg_0_14_inst : DFF_X1 port map( D => n2565, CK => n468, Q => 
                           REGISTERS_0_14_port, QN => n_1049);
   REGISTERS_reg_0_13_inst : DFF_X1 port map( D => n2564, CK => n469, Q => 
                           REGISTERS_0_13_port, QN => n_1050);
   REGISTERS_reg_0_12_inst : DFF_X1 port map( D => n2563, CK => n469, Q => 
                           REGISTERS_0_12_port, QN => n_1051);
   REGISTERS_reg_0_11_inst : DFF_X1 port map( D => n2562, CK => n469, Q => 
                           REGISTERS_0_11_port, QN => n_1052);
   REGISTERS_reg_0_10_inst : DFF_X1 port map( D => n2561, CK => n469, Q => 
                           REGISTERS_0_10_port, QN => n_1053);
   REGISTERS_reg_0_9_inst : DFF_X1 port map( D => n2560, CK => n469, Q => 
                           REGISTERS_0_9_port, QN => n_1054);
   REGISTERS_reg_0_8_inst : DFF_X1 port map( D => n2559, CK => n469, Q => 
                           REGISTERS_0_8_port, QN => n_1055);
   REGISTERS_reg_0_7_inst : DFF_X1 port map( D => n2558, CK => n469, Q => 
                           REGISTERS_0_7_port, QN => n_1056);
   REGISTERS_reg_0_6_inst : DFF_X1 port map( D => n2557, CK => n469, Q => 
                           REGISTERS_0_6_port, QN => n_1057);
   REGISTERS_reg_0_5_inst : DFF_X1 port map( D => n2556, CK => n469, Q => 
                           REGISTERS_0_5_port, QN => n_1058);
   REGISTERS_reg_0_4_inst : DFF_X1 port map( D => n2555, CK => n469, Q => 
                           REGISTERS_0_4_port, QN => n_1059);
   REGISTERS_reg_0_3_inst : DFF_X1 port map( D => n2554, CK => n469, Q => 
                           REGISTERS_0_3_port, QN => n_1060);
   REGISTERS_reg_0_2_inst : DFF_X1 port map( D => n2553, CK => n470, Q => 
                           REGISTERS_0_2_port, QN => n_1061);
   REGISTERS_reg_0_1_inst : DFF_X1 port map( D => n2552, CK => n470, Q => 
                           REGISTERS_0_1_port, QN => n_1062);
   REGISTERS_reg_0_0_inst : DFF_X1 port map( D => n2551, CK => n470, Q => 
                           REGISTERS_0_0_port, QN => n_1063);
   REGISTERS_reg_1_31_inst : DFF_X1 port map( D => n2550, CK => n470, Q => 
                           REGISTERS_1_31_port, QN => n_1064);
   REGISTERS_reg_1_30_inst : DFF_X1 port map( D => n2549, CK => n470, Q => 
                           REGISTERS_1_30_port, QN => n_1065);
   REGISTERS_reg_1_29_inst : DFF_X1 port map( D => n2548, CK => n470, Q => 
                           REGISTERS_1_29_port, QN => n_1066);
   REGISTERS_reg_1_28_inst : DFF_X1 port map( D => n2547, CK => n470, Q => 
                           REGISTERS_1_28_port, QN => n_1067);
   REGISTERS_reg_1_27_inst : DFF_X1 port map( D => n2546, CK => n470, Q => 
                           REGISTERS_1_27_port, QN => n_1068);
   REGISTERS_reg_1_26_inst : DFF_X1 port map( D => n2545, CK => n470, Q => 
                           REGISTERS_1_26_port, QN => n_1069);
   REGISTERS_reg_1_25_inst : DFF_X1 port map( D => n2544, CK => n470, Q => 
                           REGISTERS_1_25_port, QN => n_1070);
   REGISTERS_reg_1_24_inst : DFF_X1 port map( D => n2543, CK => n470, Q => 
                           REGISTERS_1_24_port, QN => n_1071);
   REGISTERS_reg_1_23_inst : DFF_X1 port map( D => n2542, CK => n471, Q => 
                           REGISTERS_1_23_port, QN => n_1072);
   REGISTERS_reg_1_22_inst : DFF_X1 port map( D => n2541, CK => n471, Q => 
                           REGISTERS_1_22_port, QN => n_1073);
   REGISTERS_reg_1_21_inst : DFF_X1 port map( D => n2540, CK => n471, Q => 
                           REGISTERS_1_21_port, QN => n_1074);
   REGISTERS_reg_1_20_inst : DFF_X1 port map( D => n2539, CK => n471, Q => 
                           REGISTERS_1_20_port, QN => n_1075);
   REGISTERS_reg_1_19_inst : DFF_X1 port map( D => n2538, CK => n471, Q => 
                           REGISTERS_1_19_port, QN => n_1076);
   REGISTERS_reg_1_18_inst : DFF_X1 port map( D => n2537, CK => n471, Q => 
                           REGISTERS_1_18_port, QN => n_1077);
   REGISTERS_reg_1_17_inst : DFF_X1 port map( D => n2536, CK => n471, Q => 
                           REGISTERS_1_17_port, QN => n_1078);
   REGISTERS_reg_1_16_inst : DFF_X1 port map( D => n2535, CK => n471, Q => 
                           REGISTERS_1_16_port, QN => n_1079);
   REGISTERS_reg_1_15_inst : DFF_X1 port map( D => n2534, CK => n471, Q => 
                           REGISTERS_1_15_port, QN => n_1080);
   REGISTERS_reg_1_14_inst : DFF_X1 port map( D => n2533, CK => n471, Q => 
                           REGISTERS_1_14_port, QN => n_1081);
   REGISTERS_reg_1_13_inst : DFF_X1 port map( D => n2532, CK => n471, Q => 
                           REGISTERS_1_13_port, QN => n_1082);
   REGISTERS_reg_1_12_inst : DFF_X1 port map( D => n2531, CK => n472, Q => 
                           REGISTERS_1_12_port, QN => n_1083);
   REGISTERS_reg_1_11_inst : DFF_X1 port map( D => n2530, CK => n472, Q => 
                           REGISTERS_1_11_port, QN => n_1084);
   REGISTERS_reg_1_10_inst : DFF_X1 port map( D => n2529, CK => n472, Q => 
                           REGISTERS_1_10_port, QN => n_1085);
   REGISTERS_reg_1_9_inst : DFF_X1 port map( D => n2528, CK => n472, Q => 
                           REGISTERS_1_9_port, QN => n_1086);
   REGISTERS_reg_1_8_inst : DFF_X1 port map( D => n2527, CK => n472, Q => 
                           REGISTERS_1_8_port, QN => n_1087);
   REGISTERS_reg_1_7_inst : DFF_X1 port map( D => n2526, CK => n472, Q => 
                           REGISTERS_1_7_port, QN => n_1088);
   REGISTERS_reg_1_6_inst : DFF_X1 port map( D => n2525, CK => n472, Q => 
                           REGISTERS_1_6_port, QN => n_1089);
   REGISTERS_reg_1_5_inst : DFF_X1 port map( D => n2524, CK => n472, Q => 
                           REGISTERS_1_5_port, QN => n_1090);
   REGISTERS_reg_1_4_inst : DFF_X1 port map( D => n2523, CK => n472, Q => 
                           REGISTERS_1_4_port, QN => n_1091);
   REGISTERS_reg_1_3_inst : DFF_X1 port map( D => n2522, CK => n472, Q => 
                           REGISTERS_1_3_port, QN => n_1092);
   REGISTERS_reg_1_2_inst : DFF_X1 port map( D => n2521, CK => n472, Q => 
                           REGISTERS_1_2_port, QN => n_1093);
   REGISTERS_reg_1_1_inst : DFF_X1 port map( D => n2520, CK => n473, Q => 
                           REGISTERS_1_1_port, QN => n_1094);
   REGISTERS_reg_1_0_inst : DFF_X1 port map( D => n2519, CK => n473, Q => 
                           REGISTERS_1_0_port, QN => n_1095);
   REGISTERS_reg_2_31_inst : DFF_X1 port map( D => n2518, CK => n473, Q => 
                           REGISTERS_2_31_port, QN => n_1096);
   REGISTERS_reg_2_30_inst : DFF_X1 port map( D => n2517, CK => n473, Q => 
                           REGISTERS_2_30_port, QN => n_1097);
   REGISTERS_reg_2_29_inst : DFF_X1 port map( D => n2516, CK => n473, Q => 
                           REGISTERS_2_29_port, QN => n_1098);
   REGISTERS_reg_2_28_inst : DFF_X1 port map( D => n2515, CK => n473, Q => 
                           REGISTERS_2_28_port, QN => n_1099);
   REGISTERS_reg_2_27_inst : DFF_X1 port map( D => n2514, CK => n473, Q => 
                           REGISTERS_2_27_port, QN => n_1100);
   REGISTERS_reg_2_26_inst : DFF_X1 port map( D => n2513, CK => n473, Q => 
                           REGISTERS_2_26_port, QN => n_1101);
   REGISTERS_reg_2_25_inst : DFF_X1 port map( D => n2512, CK => n473, Q => 
                           REGISTERS_2_25_port, QN => n_1102);
   REGISTERS_reg_2_24_inst : DFF_X1 port map( D => n2511, CK => n473, Q => 
                           REGISTERS_2_24_port, QN => n_1103);
   REGISTERS_reg_2_23_inst : DFF_X1 port map( D => n2510, CK => n473, Q => 
                           REGISTERS_2_23_port, QN => n_1104);
   REGISTERS_reg_2_22_inst : DFF_X1 port map( D => n2509, CK => n474, Q => 
                           REGISTERS_2_22_port, QN => n_1105);
   REGISTERS_reg_2_21_inst : DFF_X1 port map( D => n2508, CK => n474, Q => 
                           REGISTERS_2_21_port, QN => n_1106);
   REGISTERS_reg_2_20_inst : DFF_X1 port map( D => n2507, CK => n474, Q => 
                           REGISTERS_2_20_port, QN => n_1107);
   REGISTERS_reg_2_19_inst : DFF_X1 port map( D => n2506, CK => n474, Q => 
                           REGISTERS_2_19_port, QN => n_1108);
   REGISTERS_reg_2_18_inst : DFF_X1 port map( D => n2505, CK => n474, Q => 
                           REGISTERS_2_18_port, QN => n_1109);
   REGISTERS_reg_2_17_inst : DFF_X1 port map( D => n2504, CK => n474, Q => 
                           REGISTERS_2_17_port, QN => n_1110);
   REGISTERS_reg_2_16_inst : DFF_X1 port map( D => n2503, CK => n474, Q => 
                           REGISTERS_2_16_port, QN => n_1111);
   REGISTERS_reg_2_15_inst : DFF_X1 port map( D => n2502, CK => n474, Q => 
                           REGISTERS_2_15_port, QN => n_1112);
   REGISTERS_reg_2_14_inst : DFF_X1 port map( D => n2501, CK => n474, Q => 
                           REGISTERS_2_14_port, QN => n_1113);
   REGISTERS_reg_2_13_inst : DFF_X1 port map( D => n2500, CK => n474, Q => 
                           REGISTERS_2_13_port, QN => n_1114);
   REGISTERS_reg_2_12_inst : DFF_X1 port map( D => n2499, CK => n474, Q => 
                           REGISTERS_2_12_port, QN => n_1115);
   REGISTERS_reg_2_11_inst : DFF_X1 port map( D => n2498, CK => n475, Q => 
                           REGISTERS_2_11_port, QN => n_1116);
   REGISTERS_reg_2_10_inst : DFF_X1 port map( D => n2497, CK => n475, Q => 
                           REGISTERS_2_10_port, QN => n_1117);
   REGISTERS_reg_2_9_inst : DFF_X1 port map( D => n2496, CK => n475, Q => 
                           REGISTERS_2_9_port, QN => n_1118);
   REGISTERS_reg_2_8_inst : DFF_X1 port map( D => n2495, CK => n475, Q => 
                           REGISTERS_2_8_port, QN => n_1119);
   REGISTERS_reg_2_7_inst : DFF_X1 port map( D => n2494, CK => n475, Q => 
                           REGISTERS_2_7_port, QN => n_1120);
   REGISTERS_reg_2_6_inst : DFF_X1 port map( D => n2493, CK => n475, Q => 
                           REGISTERS_2_6_port, QN => n_1121);
   REGISTERS_reg_2_5_inst : DFF_X1 port map( D => n2492, CK => n475, Q => 
                           REGISTERS_2_5_port, QN => n_1122);
   REGISTERS_reg_2_4_inst : DFF_X1 port map( D => n2491, CK => n475, Q => 
                           REGISTERS_2_4_port, QN => n_1123);
   REGISTERS_reg_2_3_inst : DFF_X1 port map( D => n2490, CK => n475, Q => 
                           REGISTERS_2_3_port, QN => n_1124);
   REGISTERS_reg_2_2_inst : DFF_X1 port map( D => n2489, CK => n475, Q => 
                           REGISTERS_2_2_port, QN => n_1125);
   REGISTERS_reg_2_1_inst : DFF_X1 port map( D => n2488, CK => n475, Q => 
                           REGISTERS_2_1_port, QN => n_1126);
   REGISTERS_reg_2_0_inst : DFF_X1 port map( D => n2487, CK => n476, Q => 
                           REGISTERS_2_0_port, QN => n_1127);
   REGISTERS_reg_3_31_inst : DFF_X1 port map( D => n2486, CK => n476, Q => 
                           REGISTERS_3_31_port, QN => n_1128);
   REGISTERS_reg_3_30_inst : DFF_X1 port map( D => n2485, CK => n476, Q => 
                           REGISTERS_3_30_port, QN => n_1129);
   REGISTERS_reg_3_29_inst : DFF_X1 port map( D => n2484, CK => n476, Q => 
                           REGISTERS_3_29_port, QN => n_1130);
   REGISTERS_reg_3_28_inst : DFF_X1 port map( D => n2483, CK => n476, Q => 
                           REGISTERS_3_28_port, QN => n_1131);
   REGISTERS_reg_3_27_inst : DFF_X1 port map( D => n2482, CK => n476, Q => 
                           REGISTERS_3_27_port, QN => n_1132);
   REGISTERS_reg_3_26_inst : DFF_X1 port map( D => n2481, CK => n476, Q => 
                           REGISTERS_3_26_port, QN => n_1133);
   REGISTERS_reg_3_25_inst : DFF_X1 port map( D => n2480, CK => n476, Q => 
                           REGISTERS_3_25_port, QN => n_1134);
   REGISTERS_reg_3_24_inst : DFF_X1 port map( D => n2479, CK => n476, Q => 
                           REGISTERS_3_24_port, QN => n_1135);
   REGISTERS_reg_3_23_inst : DFF_X1 port map( D => n2478, CK => n476, Q => 
                           REGISTERS_3_23_port, QN => n_1136);
   REGISTERS_reg_3_22_inst : DFF_X1 port map( D => n2477, CK => n476, Q => 
                           REGISTERS_3_22_port, QN => n_1137);
   REGISTERS_reg_3_21_inst : DFF_X1 port map( D => n2476, CK => n477, Q => 
                           REGISTERS_3_21_port, QN => n_1138);
   REGISTERS_reg_3_20_inst : DFF_X1 port map( D => n2475, CK => n477, Q => 
                           REGISTERS_3_20_port, QN => n_1139);
   REGISTERS_reg_3_19_inst : DFF_X1 port map( D => n2474, CK => n477, Q => 
                           REGISTERS_3_19_port, QN => n_1140);
   REGISTERS_reg_3_18_inst : DFF_X1 port map( D => n2473, CK => n477, Q => 
                           REGISTERS_3_18_port, QN => n_1141);
   REGISTERS_reg_3_17_inst : DFF_X1 port map( D => n2472, CK => n477, Q => 
                           REGISTERS_3_17_port, QN => n_1142);
   REGISTERS_reg_3_16_inst : DFF_X1 port map( D => n2471, CK => n477, Q => 
                           REGISTERS_3_16_port, QN => n_1143);
   REGISTERS_reg_3_15_inst : DFF_X1 port map( D => n2470, CK => n477, Q => 
                           REGISTERS_3_15_port, QN => n_1144);
   REGISTERS_reg_3_14_inst : DFF_X1 port map( D => n2469, CK => n477, Q => 
                           REGISTERS_3_14_port, QN => n_1145);
   REGISTERS_reg_3_13_inst : DFF_X1 port map( D => n2468, CK => n477, Q => 
                           REGISTERS_3_13_port, QN => n_1146);
   REGISTERS_reg_3_12_inst : DFF_X1 port map( D => n2467, CK => n477, Q => 
                           REGISTERS_3_12_port, QN => n_1147);
   REGISTERS_reg_3_11_inst : DFF_X1 port map( D => n2466, CK => n477, Q => 
                           REGISTERS_3_11_port, QN => n_1148);
   REGISTERS_reg_3_10_inst : DFF_X1 port map( D => n2465, CK => n478, Q => 
                           REGISTERS_3_10_port, QN => n_1149);
   REGISTERS_reg_3_9_inst : DFF_X1 port map( D => n2464, CK => n478, Q => 
                           REGISTERS_3_9_port, QN => n_1150);
   REGISTERS_reg_3_8_inst : DFF_X1 port map( D => n2463, CK => n478, Q => 
                           REGISTERS_3_8_port, QN => n_1151);
   REGISTERS_reg_3_7_inst : DFF_X1 port map( D => n2462, CK => n478, Q => 
                           REGISTERS_3_7_port, QN => n_1152);
   REGISTERS_reg_3_6_inst : DFF_X1 port map( D => n2461, CK => n478, Q => 
                           REGISTERS_3_6_port, QN => n_1153);
   REGISTERS_reg_3_5_inst : DFF_X1 port map( D => n2460, CK => n478, Q => 
                           REGISTERS_3_5_port, QN => n_1154);
   REGISTERS_reg_3_4_inst : DFF_X1 port map( D => n2459, CK => n478, Q => 
                           REGISTERS_3_4_port, QN => n_1155);
   REGISTERS_reg_3_3_inst : DFF_X1 port map( D => n2458, CK => n478, Q => 
                           REGISTERS_3_3_port, QN => n_1156);
   REGISTERS_reg_3_2_inst : DFF_X1 port map( D => n2457, CK => n478, Q => 
                           REGISTERS_3_2_port, QN => n_1157);
   REGISTERS_reg_3_1_inst : DFF_X1 port map( D => n2456, CK => n478, Q => 
                           REGISTERS_3_1_port, QN => n_1158);
   REGISTERS_reg_3_0_inst : DFF_X1 port map( D => n2455, CK => n478, Q => 
                           REGISTERS_3_0_port, QN => n_1159);
   REGISTERS_reg_4_31_inst : DFF_X1 port map( D => n2454, CK => n479, Q => 
                           REGISTERS_4_31_port, QN => n_1160);
   REGISTERS_reg_4_30_inst : DFF_X1 port map( D => n2453, CK => n479, Q => 
                           REGISTERS_4_30_port, QN => n_1161);
   REGISTERS_reg_4_29_inst : DFF_X1 port map( D => n2452, CK => n479, Q => 
                           REGISTERS_4_29_port, QN => n_1162);
   REGISTERS_reg_4_28_inst : DFF_X1 port map( D => n2451, CK => n479, Q => 
                           REGISTERS_4_28_port, QN => n_1163);
   REGISTERS_reg_4_27_inst : DFF_X1 port map( D => n2450, CK => n479, Q => 
                           REGISTERS_4_27_port, QN => n_1164);
   REGISTERS_reg_4_26_inst : DFF_X1 port map( D => n2449, CK => n479, Q => 
                           REGISTERS_4_26_port, QN => n_1165);
   REGISTERS_reg_4_25_inst : DFF_X1 port map( D => n2448, CK => n479, Q => 
                           REGISTERS_4_25_port, QN => n_1166);
   REGISTERS_reg_4_24_inst : DFF_X1 port map( D => n2447, CK => n479, Q => 
                           REGISTERS_4_24_port, QN => n_1167);
   REGISTERS_reg_4_23_inst : DFF_X1 port map( D => n2446, CK => n479, Q => 
                           REGISTERS_4_23_port, QN => n_1168);
   REGISTERS_reg_4_22_inst : DFF_X1 port map( D => n2445, CK => n479, Q => 
                           REGISTERS_4_22_port, QN => n_1169);
   REGISTERS_reg_4_21_inst : DFF_X1 port map( D => n2444, CK => n479, Q => 
                           REGISTERS_4_21_port, QN => n_1170);
   REGISTERS_reg_4_20_inst : DFF_X1 port map( D => n2443, CK => n480, Q => 
                           REGISTERS_4_20_port, QN => n_1171);
   REGISTERS_reg_4_19_inst : DFF_X1 port map( D => n2442, CK => n480, Q => 
                           REGISTERS_4_19_port, QN => n_1172);
   REGISTERS_reg_4_18_inst : DFF_X1 port map( D => n2441, CK => n480, Q => 
                           REGISTERS_4_18_port, QN => n_1173);
   REGISTERS_reg_4_17_inst : DFF_X1 port map( D => n2440, CK => n480, Q => 
                           REGISTERS_4_17_port, QN => n_1174);
   REGISTERS_reg_4_16_inst : DFF_X1 port map( D => n2439, CK => n480, Q => 
                           REGISTERS_4_16_port, QN => n_1175);
   REGISTERS_reg_4_15_inst : DFF_X1 port map( D => n2438, CK => n480, Q => 
                           REGISTERS_4_15_port, QN => n_1176);
   REGISTERS_reg_4_14_inst : DFF_X1 port map( D => n2437, CK => n480, Q => 
                           REGISTERS_4_14_port, QN => n_1177);
   REGISTERS_reg_4_13_inst : DFF_X1 port map( D => n2436, CK => n480, Q => 
                           REGISTERS_4_13_port, QN => n_1178);
   REGISTERS_reg_4_12_inst : DFF_X1 port map( D => n2435, CK => n480, Q => 
                           REGISTERS_4_12_port, QN => n_1179);
   REGISTERS_reg_4_11_inst : DFF_X1 port map( D => n2434, CK => n480, Q => 
                           REGISTERS_4_11_port, QN => n_1180);
   REGISTERS_reg_4_10_inst : DFF_X1 port map( D => n2433, CK => n480, Q => 
                           REGISTERS_4_10_port, QN => n_1181);
   REGISTERS_reg_4_9_inst : DFF_X1 port map( D => n2432, CK => n481, Q => 
                           REGISTERS_4_9_port, QN => n_1182);
   REGISTERS_reg_4_8_inst : DFF_X1 port map( D => n2431, CK => n481, Q => 
                           REGISTERS_4_8_port, QN => n_1183);
   REGISTERS_reg_4_7_inst : DFF_X1 port map( D => n2430, CK => n481, Q => 
                           REGISTERS_4_7_port, QN => n_1184);
   REGISTERS_reg_4_6_inst : DFF_X1 port map( D => n2429, CK => n481, Q => 
                           REGISTERS_4_6_port, QN => n_1185);
   REGISTERS_reg_4_5_inst : DFF_X1 port map( D => n2428, CK => n481, Q => 
                           REGISTERS_4_5_port, QN => n_1186);
   REGISTERS_reg_4_4_inst : DFF_X1 port map( D => n2427, CK => n481, Q => 
                           REGISTERS_4_4_port, QN => n_1187);
   REGISTERS_reg_4_3_inst : DFF_X1 port map( D => n2426, CK => n481, Q => 
                           REGISTERS_4_3_port, QN => n_1188);
   REGISTERS_reg_4_2_inst : DFF_X1 port map( D => n2425, CK => n481, Q => 
                           REGISTERS_4_2_port, QN => n_1189);
   REGISTERS_reg_4_1_inst : DFF_X1 port map( D => n2424, CK => n481, Q => 
                           REGISTERS_4_1_port, QN => n_1190);
   REGISTERS_reg_4_0_inst : DFF_X1 port map( D => n2423, CK => n481, Q => 
                           REGISTERS_4_0_port, QN => n_1191);
   REGISTERS_reg_5_31_inst : DFF_X1 port map( D => n2422, CK => n481, Q => 
                           REGISTERS_5_31_port, QN => n_1192);
   REGISTERS_reg_5_30_inst : DFF_X1 port map( D => n2421, CK => n482, Q => 
                           REGISTERS_5_30_port, QN => n_1193);
   REGISTERS_reg_5_29_inst : DFF_X1 port map( D => n2420, CK => n482, Q => 
                           REGISTERS_5_29_port, QN => n_1194);
   REGISTERS_reg_5_28_inst : DFF_X1 port map( D => n2419, CK => n482, Q => 
                           REGISTERS_5_28_port, QN => n_1195);
   REGISTERS_reg_5_27_inst : DFF_X1 port map( D => n2418, CK => n482, Q => 
                           REGISTERS_5_27_port, QN => n_1196);
   REGISTERS_reg_5_26_inst : DFF_X1 port map( D => n2417, CK => n482, Q => 
                           REGISTERS_5_26_port, QN => n_1197);
   REGISTERS_reg_5_25_inst : DFF_X1 port map( D => n2416, CK => n482, Q => 
                           REGISTERS_5_25_port, QN => n_1198);
   REGISTERS_reg_5_24_inst : DFF_X1 port map( D => n2415, CK => n482, Q => 
                           REGISTERS_5_24_port, QN => n_1199);
   REGISTERS_reg_5_23_inst : DFF_X1 port map( D => n2414, CK => n482, Q => 
                           REGISTERS_5_23_port, QN => n_1200);
   REGISTERS_reg_5_22_inst : DFF_X1 port map( D => n2413, CK => n482, Q => 
                           REGISTERS_5_22_port, QN => n_1201);
   REGISTERS_reg_5_21_inst : DFF_X1 port map( D => n2412, CK => n482, Q => 
                           REGISTERS_5_21_port, QN => n_1202);
   REGISTERS_reg_5_20_inst : DFF_X1 port map( D => n2411, CK => n482, Q => 
                           REGISTERS_5_20_port, QN => n_1203);
   REGISTERS_reg_5_19_inst : DFF_X1 port map( D => n2410, CK => n483, Q => 
                           REGISTERS_5_19_port, QN => n_1204);
   REGISTERS_reg_5_18_inst : DFF_X1 port map( D => n2409, CK => n483, Q => 
                           REGISTERS_5_18_port, QN => n_1205);
   REGISTERS_reg_5_17_inst : DFF_X1 port map( D => n2408, CK => n483, Q => 
                           REGISTERS_5_17_port, QN => n_1206);
   REGISTERS_reg_5_16_inst : DFF_X1 port map( D => n2407, CK => n483, Q => 
                           REGISTERS_5_16_port, QN => n_1207);
   REGISTERS_reg_5_15_inst : DFF_X1 port map( D => n2406, CK => n483, Q => 
                           REGISTERS_5_15_port, QN => n_1208);
   REGISTERS_reg_5_14_inst : DFF_X1 port map( D => n2405, CK => n483, Q => 
                           REGISTERS_5_14_port, QN => n_1209);
   REGISTERS_reg_5_13_inst : DFF_X1 port map( D => n2404, CK => n483, Q => 
                           REGISTERS_5_13_port, QN => n_1210);
   REGISTERS_reg_5_12_inst : DFF_X1 port map( D => n2403, CK => n483, Q => 
                           REGISTERS_5_12_port, QN => n_1211);
   REGISTERS_reg_5_11_inst : DFF_X1 port map( D => n2402, CK => n483, Q => 
                           REGISTERS_5_11_port, QN => n_1212);
   REGISTERS_reg_5_10_inst : DFF_X1 port map( D => n2401, CK => n483, Q => 
                           REGISTERS_5_10_port, QN => n_1213);
   REGISTERS_reg_5_9_inst : DFF_X1 port map( D => n2400, CK => n483, Q => 
                           REGISTERS_5_9_port, QN => n_1214);
   REGISTERS_reg_5_8_inst : DFF_X1 port map( D => n2399, CK => n484, Q => 
                           REGISTERS_5_8_port, QN => n_1215);
   REGISTERS_reg_5_7_inst : DFF_X1 port map( D => n2398, CK => n484, Q => 
                           REGISTERS_5_7_port, QN => n_1216);
   REGISTERS_reg_5_6_inst : DFF_X1 port map( D => n2397, CK => n484, Q => 
                           REGISTERS_5_6_port, QN => n_1217);
   REGISTERS_reg_5_5_inst : DFF_X1 port map( D => n2396, CK => n484, Q => 
                           REGISTERS_5_5_port, QN => n_1218);
   REGISTERS_reg_5_4_inst : DFF_X1 port map( D => n2395, CK => n484, Q => 
                           REGISTERS_5_4_port, QN => n_1219);
   REGISTERS_reg_5_3_inst : DFF_X1 port map( D => n2394, CK => n484, Q => 
                           REGISTERS_5_3_port, QN => n_1220);
   REGISTERS_reg_5_2_inst : DFF_X1 port map( D => n2393, CK => n484, Q => 
                           REGISTERS_5_2_port, QN => n_1221);
   REGISTERS_reg_5_1_inst : DFF_X1 port map( D => n2392, CK => n484, Q => 
                           REGISTERS_5_1_port, QN => n_1222);
   REGISTERS_reg_5_0_inst : DFF_X1 port map( D => n2391, CK => n484, Q => 
                           REGISTERS_5_0_port, QN => n_1223);
   REGISTERS_reg_6_31_inst : DFF_X1 port map( D => n2390, CK => n484, Q => 
                           REGISTERS_6_31_port, QN => n_1224);
   REGISTERS_reg_6_30_inst : DFF_X1 port map( D => n2389, CK => n484, Q => 
                           REGISTERS_6_30_port, QN => n_1225);
   REGISTERS_reg_6_29_inst : DFF_X1 port map( D => n2388, CK => n485, Q => 
                           REGISTERS_6_29_port, QN => n_1226);
   REGISTERS_reg_6_28_inst : DFF_X1 port map( D => n2387, CK => n485, Q => 
                           REGISTERS_6_28_port, QN => n_1227);
   REGISTERS_reg_6_27_inst : DFF_X1 port map( D => n2386, CK => n485, Q => 
                           REGISTERS_6_27_port, QN => n_1228);
   REGISTERS_reg_6_26_inst : DFF_X1 port map( D => n2385, CK => n485, Q => 
                           REGISTERS_6_26_port, QN => n_1229);
   REGISTERS_reg_6_25_inst : DFF_X1 port map( D => n2384, CK => n485, Q => 
                           REGISTERS_6_25_port, QN => n_1230);
   REGISTERS_reg_6_24_inst : DFF_X1 port map( D => n2383, CK => n485, Q => 
                           REGISTERS_6_24_port, QN => n_1231);
   REGISTERS_reg_6_23_inst : DFF_X1 port map( D => n2382, CK => n485, Q => 
                           REGISTERS_6_23_port, QN => n_1232);
   REGISTERS_reg_6_22_inst : DFF_X1 port map( D => n2381, CK => n485, Q => 
                           REGISTERS_6_22_port, QN => n_1233);
   REGISTERS_reg_6_21_inst : DFF_X1 port map( D => n2380, CK => n485, Q => 
                           REGISTERS_6_21_port, QN => n_1234);
   REGISTERS_reg_6_20_inst : DFF_X1 port map( D => n2379, CK => n485, Q => 
                           REGISTERS_6_20_port, QN => n_1235);
   REGISTERS_reg_6_19_inst : DFF_X1 port map( D => n2378, CK => n485, Q => 
                           REGISTERS_6_19_port, QN => n_1236);
   REGISTERS_reg_6_18_inst : DFF_X1 port map( D => n2377, CK => n486, Q => 
                           REGISTERS_6_18_port, QN => n_1237);
   REGISTERS_reg_6_17_inst : DFF_X1 port map( D => n2376, CK => n486, Q => 
                           REGISTERS_6_17_port, QN => n_1238);
   REGISTERS_reg_6_16_inst : DFF_X1 port map( D => n2375, CK => n486, Q => 
                           REGISTERS_6_16_port, QN => n_1239);
   REGISTERS_reg_6_15_inst : DFF_X1 port map( D => n2374, CK => n486, Q => 
                           REGISTERS_6_15_port, QN => n_1240);
   REGISTERS_reg_6_14_inst : DFF_X1 port map( D => n2373, CK => n486, Q => 
                           REGISTERS_6_14_port, QN => n_1241);
   REGISTERS_reg_6_13_inst : DFF_X1 port map( D => n2372, CK => n486, Q => 
                           REGISTERS_6_13_port, QN => n_1242);
   REGISTERS_reg_6_12_inst : DFF_X1 port map( D => n2371, CK => n486, Q => 
                           REGISTERS_6_12_port, QN => n_1243);
   REGISTERS_reg_6_11_inst : DFF_X1 port map( D => n2370, CK => n486, Q => 
                           REGISTERS_6_11_port, QN => n_1244);
   REGISTERS_reg_6_10_inst : DFF_X1 port map( D => n2369, CK => n486, Q => 
                           REGISTERS_6_10_port, QN => n_1245);
   REGISTERS_reg_6_9_inst : DFF_X1 port map( D => n2368, CK => n486, Q => 
                           REGISTERS_6_9_port, QN => n_1246);
   REGISTERS_reg_6_8_inst : DFF_X1 port map( D => n2367, CK => n486, Q => 
                           REGISTERS_6_8_port, QN => n_1247);
   REGISTERS_reg_6_7_inst : DFF_X1 port map( D => n2366, CK => n487, Q => 
                           REGISTERS_6_7_port, QN => n_1248);
   REGISTERS_reg_6_6_inst : DFF_X1 port map( D => n2365, CK => n487, Q => 
                           REGISTERS_6_6_port, QN => n_1249);
   REGISTERS_reg_6_5_inst : DFF_X1 port map( D => n2364, CK => n487, Q => 
                           REGISTERS_6_5_port, QN => n_1250);
   REGISTERS_reg_6_4_inst : DFF_X1 port map( D => n2363, CK => n487, Q => 
                           REGISTERS_6_4_port, QN => n_1251);
   REGISTERS_reg_6_3_inst : DFF_X1 port map( D => n2362, CK => n487, Q => 
                           REGISTERS_6_3_port, QN => n_1252);
   REGISTERS_reg_6_2_inst : DFF_X1 port map( D => n2361, CK => n487, Q => 
                           REGISTERS_6_2_port, QN => n_1253);
   REGISTERS_reg_6_1_inst : DFF_X1 port map( D => n2360, CK => n487, Q => 
                           REGISTERS_6_1_port, QN => n_1254);
   REGISTERS_reg_6_0_inst : DFF_X1 port map( D => n2359, CK => n487, Q => 
                           REGISTERS_6_0_port, QN => n_1255);
   REGISTERS_reg_7_31_inst : DFF_X1 port map( D => n2358, CK => n487, Q => 
                           REGISTERS_7_31_port, QN => n_1256);
   REGISTERS_reg_7_30_inst : DFF_X1 port map( D => n2357, CK => n487, Q => 
                           REGISTERS_7_30_port, QN => n_1257);
   REGISTERS_reg_7_29_inst : DFF_X1 port map( D => n2356, CK => n487, Q => 
                           REGISTERS_7_29_port, QN => n_1258);
   REGISTERS_reg_7_28_inst : DFF_X1 port map( D => n2355, CK => n488, Q => 
                           REGISTERS_7_28_port, QN => n_1259);
   REGISTERS_reg_7_27_inst : DFF_X1 port map( D => n2354, CK => n488, Q => 
                           REGISTERS_7_27_port, QN => n_1260);
   REGISTERS_reg_7_26_inst : DFF_X1 port map( D => n2353, CK => n488, Q => 
                           REGISTERS_7_26_port, QN => n_1261);
   REGISTERS_reg_7_25_inst : DFF_X1 port map( D => n2352, CK => n488, Q => 
                           REGISTERS_7_25_port, QN => n_1262);
   REGISTERS_reg_7_24_inst : DFF_X1 port map( D => n2351, CK => n488, Q => 
                           REGISTERS_7_24_port, QN => n_1263);
   REGISTERS_reg_7_23_inst : DFF_X1 port map( D => n2350, CK => n488, Q => 
                           REGISTERS_7_23_port, QN => n_1264);
   REGISTERS_reg_7_22_inst : DFF_X1 port map( D => n2349, CK => n488, Q => 
                           REGISTERS_7_22_port, QN => n_1265);
   REGISTERS_reg_7_21_inst : DFF_X1 port map( D => n2348, CK => n488, Q => 
                           REGISTERS_7_21_port, QN => n_1266);
   REGISTERS_reg_7_20_inst : DFF_X1 port map( D => n2347, CK => n488, Q => 
                           REGISTERS_7_20_port, QN => n_1267);
   REGISTERS_reg_7_19_inst : DFF_X1 port map( D => n2346, CK => n488, Q => 
                           REGISTERS_7_19_port, QN => n_1268);
   REGISTERS_reg_7_18_inst : DFF_X1 port map( D => n2345, CK => n488, Q => 
                           REGISTERS_7_18_port, QN => n_1269);
   REGISTERS_reg_7_17_inst : DFF_X1 port map( D => n2344, CK => n489, Q => 
                           REGISTERS_7_17_port, QN => n_1270);
   REGISTERS_reg_7_16_inst : DFF_X1 port map( D => n2343, CK => n489, Q => 
                           REGISTERS_7_16_port, QN => n_1271);
   REGISTERS_reg_7_15_inst : DFF_X1 port map( D => n2342, CK => n489, Q => 
                           REGISTERS_7_15_port, QN => n_1272);
   REGISTERS_reg_7_14_inst : DFF_X1 port map( D => n2341, CK => n489, Q => 
                           REGISTERS_7_14_port, QN => n_1273);
   REGISTERS_reg_7_13_inst : DFF_X1 port map( D => n2340, CK => n489, Q => 
                           REGISTERS_7_13_port, QN => n_1274);
   REGISTERS_reg_7_12_inst : DFF_X1 port map( D => n2339, CK => n489, Q => 
                           REGISTERS_7_12_port, QN => n_1275);
   REGISTERS_reg_7_11_inst : DFF_X1 port map( D => n2338, CK => n489, Q => 
                           REGISTERS_7_11_port, QN => n_1276);
   REGISTERS_reg_7_10_inst : DFF_X1 port map( D => n2337, CK => n489, Q => 
                           REGISTERS_7_10_port, QN => n_1277);
   REGISTERS_reg_7_9_inst : DFF_X1 port map( D => n2336, CK => n489, Q => 
                           REGISTERS_7_9_port, QN => n_1278);
   REGISTERS_reg_7_8_inst : DFF_X1 port map( D => n2335, CK => n489, Q => 
                           REGISTERS_7_8_port, QN => n_1279);
   REGISTERS_reg_7_7_inst : DFF_X1 port map( D => n2334, CK => n489, Q => 
                           REGISTERS_7_7_port, QN => n_1280);
   REGISTERS_reg_7_6_inst : DFF_X1 port map( D => n2333, CK => n490, Q => 
                           REGISTERS_7_6_port, QN => n_1281);
   REGISTERS_reg_7_5_inst : DFF_X1 port map( D => n2332, CK => n490, Q => 
                           REGISTERS_7_5_port, QN => n_1282);
   REGISTERS_reg_7_4_inst : DFF_X1 port map( D => n2331, CK => n490, Q => 
                           REGISTERS_7_4_port, QN => n_1283);
   REGISTERS_reg_7_3_inst : DFF_X1 port map( D => n2330, CK => n490, Q => 
                           REGISTERS_7_3_port, QN => n_1284);
   REGISTERS_reg_7_2_inst : DFF_X1 port map( D => n2329, CK => n490, Q => 
                           REGISTERS_7_2_port, QN => n_1285);
   REGISTERS_reg_7_1_inst : DFF_X1 port map( D => n2328, CK => n490, Q => 
                           REGISTERS_7_1_port, QN => n_1286);
   REGISTERS_reg_7_0_inst : DFF_X1 port map( D => n2327, CK => n490, Q => 
                           REGISTERS_7_0_port, QN => n_1287);
   REGISTERS_reg_8_31_inst : DFF_X1 port map( D => n2326, CK => n490, Q => 
                           REGISTERS_8_31_port, QN => n_1288);
   REGISTERS_reg_8_30_inst : DFF_X1 port map( D => n2325, CK => n490, Q => 
                           REGISTERS_8_30_port, QN => n_1289);
   REGISTERS_reg_8_29_inst : DFF_X1 port map( D => n2324, CK => n490, Q => 
                           REGISTERS_8_29_port, QN => n_1290);
   REGISTERS_reg_8_28_inst : DFF_X1 port map( D => n2323, CK => n490, Q => 
                           REGISTERS_8_28_port, QN => n_1291);
   REGISTERS_reg_8_27_inst : DFF_X1 port map( D => n2322, CK => n491, Q => 
                           REGISTERS_8_27_port, QN => n_1292);
   REGISTERS_reg_8_26_inst : DFF_X1 port map( D => n2321, CK => n491, Q => 
                           REGISTERS_8_26_port, QN => n_1293);
   REGISTERS_reg_8_25_inst : DFF_X1 port map( D => n2320, CK => n491, Q => 
                           REGISTERS_8_25_port, QN => n_1294);
   REGISTERS_reg_8_24_inst : DFF_X1 port map( D => n2319, CK => n491, Q => 
                           REGISTERS_8_24_port, QN => n_1295);
   REGISTERS_reg_8_23_inst : DFF_X1 port map( D => n2318, CK => n491, Q => 
                           REGISTERS_8_23_port, QN => n_1296);
   REGISTERS_reg_8_22_inst : DFF_X1 port map( D => n2317, CK => n491, Q => 
                           REGISTERS_8_22_port, QN => n_1297);
   REGISTERS_reg_8_21_inst : DFF_X1 port map( D => n2316, CK => n491, Q => 
                           REGISTERS_8_21_port, QN => n_1298);
   REGISTERS_reg_8_20_inst : DFF_X1 port map( D => n2315, CK => n491, Q => 
                           REGISTERS_8_20_port, QN => n_1299);
   REGISTERS_reg_8_19_inst : DFF_X1 port map( D => n2314, CK => n491, Q => 
                           REGISTERS_8_19_port, QN => n_1300);
   REGISTERS_reg_8_18_inst : DFF_X1 port map( D => n2313, CK => n491, Q => 
                           REGISTERS_8_18_port, QN => n_1301);
   REGISTERS_reg_8_17_inst : DFF_X1 port map( D => n2312, CK => n491, Q => 
                           REGISTERS_8_17_port, QN => n_1302);
   REGISTERS_reg_8_16_inst : DFF_X1 port map( D => n2311, CK => n492, Q => 
                           REGISTERS_8_16_port, QN => n_1303);
   REGISTERS_reg_8_15_inst : DFF_X1 port map( D => n2310, CK => n492, Q => 
                           REGISTERS_8_15_port, QN => n_1304);
   REGISTERS_reg_8_14_inst : DFF_X1 port map( D => n2309, CK => n492, Q => 
                           REGISTERS_8_14_port, QN => n_1305);
   REGISTERS_reg_8_13_inst : DFF_X1 port map( D => n2308, CK => n492, Q => 
                           REGISTERS_8_13_port, QN => n_1306);
   REGISTERS_reg_8_12_inst : DFF_X1 port map( D => n2307, CK => n492, Q => 
                           REGISTERS_8_12_port, QN => n_1307);
   REGISTERS_reg_8_11_inst : DFF_X1 port map( D => n2306, CK => n492, Q => 
                           REGISTERS_8_11_port, QN => n_1308);
   REGISTERS_reg_8_10_inst : DFF_X1 port map( D => n2305, CK => n492, Q => 
                           REGISTERS_8_10_port, QN => n_1309);
   REGISTERS_reg_8_9_inst : DFF_X1 port map( D => n2304, CK => n492, Q => 
                           REGISTERS_8_9_port, QN => n_1310);
   REGISTERS_reg_8_8_inst : DFF_X1 port map( D => n2303, CK => n492, Q => 
                           REGISTERS_8_8_port, QN => n_1311);
   REGISTERS_reg_8_7_inst : DFF_X1 port map( D => n2302, CK => n492, Q => 
                           REGISTERS_8_7_port, QN => n_1312);
   REGISTERS_reg_8_6_inst : DFF_X1 port map( D => n2301, CK => n492, Q => 
                           REGISTERS_8_6_port, QN => n_1313);
   REGISTERS_reg_8_5_inst : DFF_X1 port map( D => n2300, CK => n493, Q => 
                           REGISTERS_8_5_port, QN => n_1314);
   REGISTERS_reg_8_4_inst : DFF_X1 port map( D => n2299, CK => n493, Q => 
                           REGISTERS_8_4_port, QN => n_1315);
   REGISTERS_reg_8_3_inst : DFF_X1 port map( D => n2298, CK => n493, Q => 
                           REGISTERS_8_3_port, QN => n_1316);
   REGISTERS_reg_8_2_inst : DFF_X1 port map( D => n2297, CK => n493, Q => 
                           REGISTERS_8_2_port, QN => n_1317);
   REGISTERS_reg_8_1_inst : DFF_X1 port map( D => n2296, CK => n493, Q => 
                           REGISTERS_8_1_port, QN => n_1318);
   REGISTERS_reg_8_0_inst : DFF_X1 port map( D => n2295, CK => n493, Q => 
                           REGISTERS_8_0_port, QN => n_1319);
   REGISTERS_reg_9_31_inst : DFF_X1 port map( D => n2294, CK => n493, Q => 
                           REGISTERS_9_31_port, QN => n_1320);
   REGISTERS_reg_9_30_inst : DFF_X1 port map( D => n2293, CK => n493, Q => 
                           REGISTERS_9_30_port, QN => n_1321);
   REGISTERS_reg_9_29_inst : DFF_X1 port map( D => n2292, CK => n493, Q => 
                           REGISTERS_9_29_port, QN => n_1322);
   REGISTERS_reg_9_28_inst : DFF_X1 port map( D => n2291, CK => n493, Q => 
                           REGISTERS_9_28_port, QN => n_1323);
   REGISTERS_reg_9_27_inst : DFF_X1 port map( D => n2290, CK => n493, Q => 
                           REGISTERS_9_27_port, QN => n_1324);
   REGISTERS_reg_9_26_inst : DFF_X1 port map( D => n2289, CK => n494, Q => 
                           REGISTERS_9_26_port, QN => n_1325);
   REGISTERS_reg_9_25_inst : DFF_X1 port map( D => n2288, CK => n494, Q => 
                           REGISTERS_9_25_port, QN => n_1326);
   REGISTERS_reg_9_24_inst : DFF_X1 port map( D => n2287, CK => n494, Q => 
                           REGISTERS_9_24_port, QN => n_1327);
   REGISTERS_reg_9_23_inst : DFF_X1 port map( D => n2286, CK => n494, Q => 
                           REGISTERS_9_23_port, QN => n_1328);
   REGISTERS_reg_9_22_inst : DFF_X1 port map( D => n2285, CK => n494, Q => 
                           REGISTERS_9_22_port, QN => n_1329);
   REGISTERS_reg_9_21_inst : DFF_X1 port map( D => n2284, CK => n494, Q => 
                           REGISTERS_9_21_port, QN => n_1330);
   REGISTERS_reg_9_20_inst : DFF_X1 port map( D => n2283, CK => n494, Q => 
                           REGISTERS_9_20_port, QN => n_1331);
   REGISTERS_reg_9_19_inst : DFF_X1 port map( D => n2282, CK => n494, Q => 
                           REGISTERS_9_19_port, QN => n_1332);
   REGISTERS_reg_9_18_inst : DFF_X1 port map( D => n2281, CK => n494, Q => 
                           REGISTERS_9_18_port, QN => n_1333);
   REGISTERS_reg_9_17_inst : DFF_X1 port map( D => n2280, CK => n494, Q => 
                           REGISTERS_9_17_port, QN => n_1334);
   REGISTERS_reg_9_16_inst : DFF_X1 port map( D => n2279, CK => n494, Q => 
                           REGISTERS_9_16_port, QN => n_1335);
   REGISTERS_reg_9_15_inst : DFF_X1 port map( D => n2278, CK => n495, Q => 
                           REGISTERS_9_15_port, QN => n_1336);
   REGISTERS_reg_9_14_inst : DFF_X1 port map( D => n2277, CK => n495, Q => 
                           REGISTERS_9_14_port, QN => n_1337);
   REGISTERS_reg_9_13_inst : DFF_X1 port map( D => n2276, CK => n495, Q => 
                           REGISTERS_9_13_port, QN => n_1338);
   REGISTERS_reg_9_12_inst : DFF_X1 port map( D => n2275, CK => n495, Q => 
                           REGISTERS_9_12_port, QN => n_1339);
   REGISTERS_reg_9_11_inst : DFF_X1 port map( D => n2274, CK => n495, Q => 
                           REGISTERS_9_11_port, QN => n_1340);
   REGISTERS_reg_9_10_inst : DFF_X1 port map( D => n2273, CK => n495, Q => 
                           REGISTERS_9_10_port, QN => n_1341);
   REGISTERS_reg_9_9_inst : DFF_X1 port map( D => n2272, CK => n495, Q => 
                           REGISTERS_9_9_port, QN => n_1342);
   REGISTERS_reg_9_8_inst : DFF_X1 port map( D => n2271, CK => n495, Q => 
                           REGISTERS_9_8_port, QN => n_1343);
   REGISTERS_reg_9_7_inst : DFF_X1 port map( D => n2270, CK => n495, Q => 
                           REGISTERS_9_7_port, QN => n_1344);
   REGISTERS_reg_9_6_inst : DFF_X1 port map( D => n2269, CK => n495, Q => 
                           REGISTERS_9_6_port, QN => n_1345);
   REGISTERS_reg_9_5_inst : DFF_X1 port map( D => n2268, CK => n495, Q => 
                           REGISTERS_9_5_port, QN => n_1346);
   REGISTERS_reg_9_4_inst : DFF_X1 port map( D => n2267, CK => n496, Q => 
                           REGISTERS_9_4_port, QN => n_1347);
   REGISTERS_reg_9_3_inst : DFF_X1 port map( D => n2266, CK => n496, Q => 
                           REGISTERS_9_3_port, QN => n_1348);
   REGISTERS_reg_9_2_inst : DFF_X1 port map( D => n2265, CK => n496, Q => 
                           REGISTERS_9_2_port, QN => n_1349);
   REGISTERS_reg_9_1_inst : DFF_X1 port map( D => n2264, CK => n496, Q => 
                           REGISTERS_9_1_port, QN => n_1350);
   REGISTERS_reg_9_0_inst : DFF_X1 port map( D => n2263, CK => n496, Q => 
                           REGISTERS_9_0_port, QN => n_1351);
   REGISTERS_reg_10_31_inst : DFF_X1 port map( D => n2262, CK => n496, Q => 
                           REGISTERS_10_31_port, QN => n_1352);
   REGISTERS_reg_10_30_inst : DFF_X1 port map( D => n2261, CK => n496, Q => 
                           REGISTERS_10_30_port, QN => n_1353);
   REGISTERS_reg_10_29_inst : DFF_X1 port map( D => n2260, CK => n496, Q => 
                           REGISTERS_10_29_port, QN => n_1354);
   REGISTERS_reg_10_28_inst : DFF_X1 port map( D => n2259, CK => n496, Q => 
                           REGISTERS_10_28_port, QN => n_1355);
   REGISTERS_reg_10_27_inst : DFF_X1 port map( D => n2258, CK => n496, Q => 
                           REGISTERS_10_27_port, QN => n_1356);
   REGISTERS_reg_10_26_inst : DFF_X1 port map( D => n2257, CK => n496, Q => 
                           REGISTERS_10_26_port, QN => n_1357);
   REGISTERS_reg_10_25_inst : DFF_X1 port map( D => n2256, CK => n497, Q => 
                           REGISTERS_10_25_port, QN => n_1358);
   REGISTERS_reg_10_24_inst : DFF_X1 port map( D => n2255, CK => n497, Q => 
                           REGISTERS_10_24_port, QN => n_1359);
   REGISTERS_reg_10_23_inst : DFF_X1 port map( D => n2254, CK => n497, Q => 
                           REGISTERS_10_23_port, QN => n_1360);
   REGISTERS_reg_10_22_inst : DFF_X1 port map( D => n2253, CK => n497, Q => 
                           REGISTERS_10_22_port, QN => n_1361);
   REGISTERS_reg_10_21_inst : DFF_X1 port map( D => n2252, CK => n497, Q => 
                           REGISTERS_10_21_port, QN => n_1362);
   REGISTERS_reg_10_20_inst : DFF_X1 port map( D => n2251, CK => n497, Q => 
                           REGISTERS_10_20_port, QN => n_1363);
   REGISTERS_reg_10_19_inst : DFF_X1 port map( D => n2250, CK => n497, Q => 
                           REGISTERS_10_19_port, QN => n_1364);
   REGISTERS_reg_10_18_inst : DFF_X1 port map( D => n2249, CK => n497, Q => 
                           REGISTERS_10_18_port, QN => n_1365);
   REGISTERS_reg_10_17_inst : DFF_X1 port map( D => n2248, CK => n497, Q => 
                           REGISTERS_10_17_port, QN => n_1366);
   REGISTERS_reg_10_16_inst : DFF_X1 port map( D => n2247, CK => n497, Q => 
                           REGISTERS_10_16_port, QN => n_1367);
   REGISTERS_reg_10_15_inst : DFF_X1 port map( D => n2246, CK => n497, Q => 
                           REGISTERS_10_15_port, QN => n_1368);
   REGISTERS_reg_10_14_inst : DFF_X1 port map( D => n2245, CK => n498, Q => 
                           REGISTERS_10_14_port, QN => n_1369);
   REGISTERS_reg_10_13_inst : DFF_X1 port map( D => n2244, CK => n498, Q => 
                           REGISTERS_10_13_port, QN => n_1370);
   REGISTERS_reg_10_12_inst : DFF_X1 port map( D => n2243, CK => n498, Q => 
                           REGISTERS_10_12_port, QN => n_1371);
   REGISTERS_reg_10_11_inst : DFF_X1 port map( D => n2242, CK => n498, Q => 
                           REGISTERS_10_11_port, QN => n_1372);
   REGISTERS_reg_10_10_inst : DFF_X1 port map( D => n2241, CK => n498, Q => 
                           REGISTERS_10_10_port, QN => n_1373);
   REGISTERS_reg_10_9_inst : DFF_X1 port map( D => n2240, CK => n498, Q => 
                           REGISTERS_10_9_port, QN => n_1374);
   REGISTERS_reg_10_8_inst : DFF_X1 port map( D => n2239, CK => n498, Q => 
                           REGISTERS_10_8_port, QN => n_1375);
   REGISTERS_reg_10_7_inst : DFF_X1 port map( D => n2238, CK => n498, Q => 
                           REGISTERS_10_7_port, QN => n_1376);
   REGISTERS_reg_10_6_inst : DFF_X1 port map( D => n2237, CK => n498, Q => 
                           REGISTERS_10_6_port, QN => n_1377);
   REGISTERS_reg_10_5_inst : DFF_X1 port map( D => n2236, CK => n498, Q => 
                           REGISTERS_10_5_port, QN => n_1378);
   REGISTERS_reg_10_4_inst : DFF_X1 port map( D => n2235, CK => n498, Q => 
                           REGISTERS_10_4_port, QN => n_1379);
   REGISTERS_reg_10_3_inst : DFF_X1 port map( D => n2234, CK => n499, Q => 
                           REGISTERS_10_3_port, QN => n_1380);
   REGISTERS_reg_10_2_inst : DFF_X1 port map( D => n2233, CK => n499, Q => 
                           REGISTERS_10_2_port, QN => n_1381);
   REGISTERS_reg_10_1_inst : DFF_X1 port map( D => n2232, CK => n499, Q => 
                           REGISTERS_10_1_port, QN => n_1382);
   REGISTERS_reg_10_0_inst : DFF_X1 port map( D => n2231, CK => n499, Q => 
                           REGISTERS_10_0_port, QN => n_1383);
   REGISTERS_reg_11_31_inst : DFF_X1 port map( D => n2230, CK => n499, Q => 
                           REGISTERS_11_31_port, QN => n_1384);
   REGISTERS_reg_11_30_inst : DFF_X1 port map( D => n2229, CK => n499, Q => 
                           REGISTERS_11_30_port, QN => n_1385);
   REGISTERS_reg_11_29_inst : DFF_X1 port map( D => n2228, CK => n499, Q => 
                           REGISTERS_11_29_port, QN => n_1386);
   REGISTERS_reg_11_28_inst : DFF_X1 port map( D => n2227, CK => n499, Q => 
                           REGISTERS_11_28_port, QN => n_1387);
   REGISTERS_reg_11_27_inst : DFF_X1 port map( D => n2226, CK => n499, Q => 
                           REGISTERS_11_27_port, QN => n_1388);
   REGISTERS_reg_11_26_inst : DFF_X1 port map( D => n2225, CK => n499, Q => 
                           REGISTERS_11_26_port, QN => n_1389);
   REGISTERS_reg_11_25_inst : DFF_X1 port map( D => n2224, CK => n499, Q => 
                           REGISTERS_11_25_port, QN => n_1390);
   REGISTERS_reg_11_24_inst : DFF_X1 port map( D => n2223, CK => n500, Q => 
                           REGISTERS_11_24_port, QN => n_1391);
   REGISTERS_reg_11_23_inst : DFF_X1 port map( D => n2222, CK => n500, Q => 
                           REGISTERS_11_23_port, QN => n_1392);
   REGISTERS_reg_11_22_inst : DFF_X1 port map( D => n2221, CK => n500, Q => 
                           REGISTERS_11_22_port, QN => n_1393);
   REGISTERS_reg_11_21_inst : DFF_X1 port map( D => n2220, CK => n500, Q => 
                           REGISTERS_11_21_port, QN => n_1394);
   REGISTERS_reg_11_20_inst : DFF_X1 port map( D => n2219, CK => n500, Q => 
                           REGISTERS_11_20_port, QN => n_1395);
   REGISTERS_reg_11_19_inst : DFF_X1 port map( D => n2218, CK => n500, Q => 
                           REGISTERS_11_19_port, QN => n_1396);
   REGISTERS_reg_11_18_inst : DFF_X1 port map( D => n2217, CK => n500, Q => 
                           REGISTERS_11_18_port, QN => n_1397);
   REGISTERS_reg_11_17_inst : DFF_X1 port map( D => n2216, CK => n500, Q => 
                           REGISTERS_11_17_port, QN => n_1398);
   REGISTERS_reg_11_16_inst : DFF_X1 port map( D => n2215, CK => n500, Q => 
                           REGISTERS_11_16_port, QN => n_1399);
   REGISTERS_reg_11_15_inst : DFF_X1 port map( D => n2214, CK => n500, Q => 
                           REGISTERS_11_15_port, QN => n_1400);
   REGISTERS_reg_11_14_inst : DFF_X1 port map( D => n2213, CK => n500, Q => 
                           REGISTERS_11_14_port, QN => n_1401);
   REGISTERS_reg_11_13_inst : DFF_X1 port map( D => n2212, CK => n501, Q => 
                           REGISTERS_11_13_port, QN => n_1402);
   REGISTERS_reg_11_12_inst : DFF_X1 port map( D => n2211, CK => n501, Q => 
                           REGISTERS_11_12_port, QN => n_1403);
   REGISTERS_reg_11_11_inst : DFF_X1 port map( D => n2210, CK => n501, Q => 
                           REGISTERS_11_11_port, QN => n_1404);
   REGISTERS_reg_11_10_inst : DFF_X1 port map( D => n2209, CK => n501, Q => 
                           REGISTERS_11_10_port, QN => n_1405);
   REGISTERS_reg_11_9_inst : DFF_X1 port map( D => n2208, CK => n501, Q => 
                           REGISTERS_11_9_port, QN => n_1406);
   REGISTERS_reg_11_8_inst : DFF_X1 port map( D => n2207, CK => n501, Q => 
                           REGISTERS_11_8_port, QN => n_1407);
   REGISTERS_reg_11_7_inst : DFF_X1 port map( D => n2206, CK => n501, Q => 
                           REGISTERS_11_7_port, QN => n_1408);
   REGISTERS_reg_11_6_inst : DFF_X1 port map( D => n2205, CK => n501, Q => 
                           REGISTERS_11_6_port, QN => n_1409);
   REGISTERS_reg_11_5_inst : DFF_X1 port map( D => n2204, CK => n501, Q => 
                           REGISTERS_11_5_port, QN => n_1410);
   REGISTERS_reg_11_4_inst : DFF_X1 port map( D => n2203, CK => n501, Q => 
                           REGISTERS_11_4_port, QN => n_1411);
   REGISTERS_reg_11_3_inst : DFF_X1 port map( D => n2202, CK => n501, Q => 
                           REGISTERS_11_3_port, QN => n_1412);
   REGISTERS_reg_11_2_inst : DFF_X1 port map( D => n2201, CK => n502, Q => 
                           REGISTERS_11_2_port, QN => n_1413);
   REGISTERS_reg_11_1_inst : DFF_X1 port map( D => n2200, CK => n502, Q => 
                           REGISTERS_11_1_port, QN => n_1414);
   REGISTERS_reg_11_0_inst : DFF_X1 port map( D => n2199, CK => n502, Q => 
                           REGISTERS_11_0_port, QN => n_1415);
   REGISTERS_reg_12_31_inst : DFF_X1 port map( D => n2198, CK => n502, Q => 
                           REGISTERS_12_31_port, QN => n_1416);
   REGISTERS_reg_12_30_inst : DFF_X1 port map( D => n2197, CK => n502, Q => 
                           REGISTERS_12_30_port, QN => n_1417);
   REGISTERS_reg_12_29_inst : DFF_X1 port map( D => n2196, CK => n502, Q => 
                           REGISTERS_12_29_port, QN => n_1418);
   REGISTERS_reg_12_28_inst : DFF_X1 port map( D => n2195, CK => n502, Q => 
                           REGISTERS_12_28_port, QN => n_1419);
   REGISTERS_reg_12_27_inst : DFF_X1 port map( D => n2194, CK => n502, Q => 
                           REGISTERS_12_27_port, QN => n_1420);
   REGISTERS_reg_12_26_inst : DFF_X1 port map( D => n2193, CK => n502, Q => 
                           REGISTERS_12_26_port, QN => n_1421);
   REGISTERS_reg_12_25_inst : DFF_X1 port map( D => n2192, CK => n502, Q => 
                           REGISTERS_12_25_port, QN => n_1422);
   REGISTERS_reg_12_24_inst : DFF_X1 port map( D => n2191, CK => n502, Q => 
                           REGISTERS_12_24_port, QN => n_1423);
   REGISTERS_reg_12_23_inst : DFF_X1 port map( D => n2190, CK => n503, Q => 
                           REGISTERS_12_23_port, QN => n_1424);
   REGISTERS_reg_12_22_inst : DFF_X1 port map( D => n2189, CK => n503, Q => 
                           REGISTERS_12_22_port, QN => n_1425);
   REGISTERS_reg_12_21_inst : DFF_X1 port map( D => n2188, CK => n503, Q => 
                           REGISTERS_12_21_port, QN => n_1426);
   REGISTERS_reg_12_20_inst : DFF_X1 port map( D => n2187, CK => n503, Q => 
                           REGISTERS_12_20_port, QN => n_1427);
   REGISTERS_reg_12_19_inst : DFF_X1 port map( D => n2186, CK => n503, Q => 
                           REGISTERS_12_19_port, QN => n_1428);
   REGISTERS_reg_12_18_inst : DFF_X1 port map( D => n2185, CK => n503, Q => 
                           REGISTERS_12_18_port, QN => n_1429);
   REGISTERS_reg_12_17_inst : DFF_X1 port map( D => n2184, CK => n503, Q => 
                           REGISTERS_12_17_port, QN => n_1430);
   REGISTERS_reg_12_16_inst : DFF_X1 port map( D => n2183, CK => n503, Q => 
                           REGISTERS_12_16_port, QN => n_1431);
   REGISTERS_reg_12_15_inst : DFF_X1 port map( D => n2182, CK => n503, Q => 
                           REGISTERS_12_15_port, QN => n_1432);
   REGISTERS_reg_12_14_inst : DFF_X1 port map( D => n2181, CK => n503, Q => 
                           REGISTERS_12_14_port, QN => n_1433);
   REGISTERS_reg_12_13_inst : DFF_X1 port map( D => n2180, CK => n503, Q => 
                           REGISTERS_12_13_port, QN => n_1434);
   REGISTERS_reg_12_12_inst : DFF_X1 port map( D => n2179, CK => n504, Q => 
                           REGISTERS_12_12_port, QN => n_1435);
   REGISTERS_reg_12_11_inst : DFF_X1 port map( D => n2178, CK => n504, Q => 
                           REGISTERS_12_11_port, QN => n_1436);
   REGISTERS_reg_12_10_inst : DFF_X1 port map( D => n2177, CK => n504, Q => 
                           REGISTERS_12_10_port, QN => n_1437);
   REGISTERS_reg_12_9_inst : DFF_X1 port map( D => n2176, CK => n504, Q => 
                           REGISTERS_12_9_port, QN => n_1438);
   REGISTERS_reg_12_8_inst : DFF_X1 port map( D => n2175, CK => n504, Q => 
                           REGISTERS_12_8_port, QN => n_1439);
   REGISTERS_reg_12_7_inst : DFF_X1 port map( D => n2174, CK => n504, Q => 
                           REGISTERS_12_7_port, QN => n_1440);
   REGISTERS_reg_12_6_inst : DFF_X1 port map( D => n2173, CK => n504, Q => 
                           REGISTERS_12_6_port, QN => n_1441);
   REGISTERS_reg_12_5_inst : DFF_X1 port map( D => n2172, CK => n504, Q => 
                           REGISTERS_12_5_port, QN => n_1442);
   REGISTERS_reg_12_4_inst : DFF_X1 port map( D => n2171, CK => n504, Q => 
                           REGISTERS_12_4_port, QN => n_1443);
   REGISTERS_reg_12_3_inst : DFF_X1 port map( D => n2170, CK => n504, Q => 
                           REGISTERS_12_3_port, QN => n_1444);
   REGISTERS_reg_12_2_inst : DFF_X1 port map( D => n2169, CK => n504, Q => 
                           REGISTERS_12_2_port, QN => n_1445);
   REGISTERS_reg_12_1_inst : DFF_X1 port map( D => n2168, CK => n505, Q => 
                           REGISTERS_12_1_port, QN => n_1446);
   REGISTERS_reg_12_0_inst : DFF_X1 port map( D => n2167, CK => n505, Q => 
                           REGISTERS_12_0_port, QN => n_1447);
   REGISTERS_reg_13_31_inst : DFF_X1 port map( D => n2166, CK => n505, Q => 
                           REGISTERS_13_31_port, QN => n_1448);
   REGISTERS_reg_13_30_inst : DFF_X1 port map( D => n2165, CK => n505, Q => 
                           REGISTERS_13_30_port, QN => n_1449);
   REGISTERS_reg_13_29_inst : DFF_X1 port map( D => n2164, CK => n505, Q => 
                           REGISTERS_13_29_port, QN => n_1450);
   REGISTERS_reg_13_28_inst : DFF_X1 port map( D => n2163, CK => n505, Q => 
                           REGISTERS_13_28_port, QN => n_1451);
   REGISTERS_reg_13_27_inst : DFF_X1 port map( D => n2162, CK => n505, Q => 
                           REGISTERS_13_27_port, QN => n_1452);
   REGISTERS_reg_13_26_inst : DFF_X1 port map( D => n2161, CK => n505, Q => 
                           REGISTERS_13_26_port, QN => n_1453);
   REGISTERS_reg_13_25_inst : DFF_X1 port map( D => n2160, CK => n505, Q => 
                           REGISTERS_13_25_port, QN => n_1454);
   REGISTERS_reg_13_24_inst : DFF_X1 port map( D => n2159, CK => n505, Q => 
                           REGISTERS_13_24_port, QN => n_1455);
   REGISTERS_reg_13_23_inst : DFF_X1 port map( D => n2158, CK => n505, Q => 
                           REGISTERS_13_23_port, QN => n_1456);
   REGISTERS_reg_13_22_inst : DFF_X1 port map( D => n2157, CK => n506, Q => 
                           REGISTERS_13_22_port, QN => n_1457);
   REGISTERS_reg_13_21_inst : DFF_X1 port map( D => n2156, CK => n506, Q => 
                           REGISTERS_13_21_port, QN => n_1458);
   REGISTERS_reg_13_20_inst : DFF_X1 port map( D => n2155, CK => n506, Q => 
                           REGISTERS_13_20_port, QN => n_1459);
   REGISTERS_reg_13_19_inst : DFF_X1 port map( D => n2154, CK => n506, Q => 
                           REGISTERS_13_19_port, QN => n_1460);
   REGISTERS_reg_13_18_inst : DFF_X1 port map( D => n2153, CK => n506, Q => 
                           REGISTERS_13_18_port, QN => n_1461);
   REGISTERS_reg_13_17_inst : DFF_X1 port map( D => n2152, CK => n506, Q => 
                           REGISTERS_13_17_port, QN => n_1462);
   REGISTERS_reg_13_16_inst : DFF_X1 port map( D => n2151, CK => n506, Q => 
                           REGISTERS_13_16_port, QN => n_1463);
   REGISTERS_reg_13_15_inst : DFF_X1 port map( D => n2150, CK => n506, Q => 
                           REGISTERS_13_15_port, QN => n_1464);
   REGISTERS_reg_13_14_inst : DFF_X1 port map( D => n2149, CK => n506, Q => 
                           REGISTERS_13_14_port, QN => n_1465);
   REGISTERS_reg_13_13_inst : DFF_X1 port map( D => n2148, CK => n506, Q => 
                           REGISTERS_13_13_port, QN => n_1466);
   REGISTERS_reg_13_12_inst : DFF_X1 port map( D => n2147, CK => n506, Q => 
                           REGISTERS_13_12_port, QN => n_1467);
   REGISTERS_reg_13_11_inst : DFF_X1 port map( D => n2146, CK => n507, Q => 
                           REGISTERS_13_11_port, QN => n_1468);
   REGISTERS_reg_13_10_inst : DFF_X1 port map( D => n2145, CK => n507, Q => 
                           REGISTERS_13_10_port, QN => n_1469);
   REGISTERS_reg_13_9_inst : DFF_X1 port map( D => n2144, CK => n507, Q => 
                           REGISTERS_13_9_port, QN => n_1470);
   REGISTERS_reg_13_8_inst : DFF_X1 port map( D => n2143, CK => n507, Q => 
                           REGISTERS_13_8_port, QN => n_1471);
   REGISTERS_reg_13_7_inst : DFF_X1 port map( D => n2142, CK => n507, Q => 
                           REGISTERS_13_7_port, QN => n_1472);
   REGISTERS_reg_13_6_inst : DFF_X1 port map( D => n2141, CK => n507, Q => 
                           REGISTERS_13_6_port, QN => n_1473);
   REGISTERS_reg_13_5_inst : DFF_X1 port map( D => n2140, CK => n507, Q => 
                           REGISTERS_13_5_port, QN => n_1474);
   REGISTERS_reg_13_4_inst : DFF_X1 port map( D => n2139, CK => n507, Q => 
                           REGISTERS_13_4_port, QN => n_1475);
   REGISTERS_reg_13_3_inst : DFF_X1 port map( D => n2138, CK => n507, Q => 
                           REGISTERS_13_3_port, QN => n_1476);
   REGISTERS_reg_13_2_inst : DFF_X1 port map( D => n2137, CK => n507, Q => 
                           REGISTERS_13_2_port, QN => n_1477);
   REGISTERS_reg_13_1_inst : DFF_X1 port map( D => n2136, CK => n507, Q => 
                           REGISTERS_13_1_port, QN => n_1478);
   REGISTERS_reg_13_0_inst : DFF_X1 port map( D => n2135, CK => n508, Q => 
                           REGISTERS_13_0_port, QN => n_1479);
   REGISTERS_reg_14_31_inst : DFF_X1 port map( D => n2134, CK => n508, Q => 
                           REGISTERS_14_31_port, QN => n_1480);
   REGISTERS_reg_14_30_inst : DFF_X1 port map( D => n2133, CK => n508, Q => 
                           REGISTERS_14_30_port, QN => n_1481);
   REGISTERS_reg_14_29_inst : DFF_X1 port map( D => n2132, CK => n508, Q => 
                           REGISTERS_14_29_port, QN => n_1482);
   REGISTERS_reg_14_28_inst : DFF_X1 port map( D => n2131, CK => n508, Q => 
                           REGISTERS_14_28_port, QN => n_1483);
   REGISTERS_reg_14_27_inst : DFF_X1 port map( D => n2130, CK => n508, Q => 
                           REGISTERS_14_27_port, QN => n_1484);
   REGISTERS_reg_14_26_inst : DFF_X1 port map( D => n2129, CK => n508, Q => 
                           REGISTERS_14_26_port, QN => n_1485);
   REGISTERS_reg_14_25_inst : DFF_X1 port map( D => n2128, CK => n508, Q => 
                           REGISTERS_14_25_port, QN => n_1486);
   REGISTERS_reg_14_24_inst : DFF_X1 port map( D => n2127, CK => n508, Q => 
                           REGISTERS_14_24_port, QN => n_1487);
   REGISTERS_reg_14_23_inst : DFF_X1 port map( D => n2126, CK => n508, Q => 
                           REGISTERS_14_23_port, QN => n_1488);
   REGISTERS_reg_14_22_inst : DFF_X1 port map( D => n2125, CK => n508, Q => 
                           REGISTERS_14_22_port, QN => n_1489);
   REGISTERS_reg_14_21_inst : DFF_X1 port map( D => n2124, CK => n509, Q => 
                           REGISTERS_14_21_port, QN => n_1490);
   REGISTERS_reg_14_20_inst : DFF_X1 port map( D => n2123, CK => n509, Q => 
                           REGISTERS_14_20_port, QN => n_1491);
   REGISTERS_reg_14_19_inst : DFF_X1 port map( D => n2122, CK => n509, Q => 
                           REGISTERS_14_19_port, QN => n_1492);
   REGISTERS_reg_14_18_inst : DFF_X1 port map( D => n2121, CK => n509, Q => 
                           REGISTERS_14_18_port, QN => n_1493);
   REGISTERS_reg_14_17_inst : DFF_X1 port map( D => n2120, CK => n509, Q => 
                           REGISTERS_14_17_port, QN => n_1494);
   REGISTERS_reg_14_16_inst : DFF_X1 port map( D => n2119, CK => n509, Q => 
                           REGISTERS_14_16_port, QN => n_1495);
   REGISTERS_reg_14_15_inst : DFF_X1 port map( D => n2118, CK => n509, Q => 
                           REGISTERS_14_15_port, QN => n_1496);
   REGISTERS_reg_14_14_inst : DFF_X1 port map( D => n2117, CK => n509, Q => 
                           REGISTERS_14_14_port, QN => n_1497);
   REGISTERS_reg_14_13_inst : DFF_X1 port map( D => n2116, CK => n509, Q => 
                           REGISTERS_14_13_port, QN => n_1498);
   REGISTERS_reg_14_12_inst : DFF_X1 port map( D => n2115, CK => n509, Q => 
                           REGISTERS_14_12_port, QN => n_1499);
   REGISTERS_reg_14_11_inst : DFF_X1 port map( D => n2114, CK => n509, Q => 
                           REGISTERS_14_11_port, QN => n_1500);
   REGISTERS_reg_14_10_inst : DFF_X1 port map( D => n2113, CK => n510, Q => 
                           REGISTERS_14_10_port, QN => n_1501);
   REGISTERS_reg_14_9_inst : DFF_X1 port map( D => n2112, CK => n510, Q => 
                           REGISTERS_14_9_port, QN => n_1502);
   REGISTERS_reg_14_8_inst : DFF_X1 port map( D => n2111, CK => n510, Q => 
                           REGISTERS_14_8_port, QN => n_1503);
   REGISTERS_reg_14_7_inst : DFF_X1 port map( D => n2110, CK => n510, Q => 
                           REGISTERS_14_7_port, QN => n_1504);
   REGISTERS_reg_14_6_inst : DFF_X1 port map( D => n2109, CK => n510, Q => 
                           REGISTERS_14_6_port, QN => n_1505);
   REGISTERS_reg_14_5_inst : DFF_X1 port map( D => n2108, CK => n510, Q => 
                           REGISTERS_14_5_port, QN => n_1506);
   REGISTERS_reg_14_4_inst : DFF_X1 port map( D => n2107, CK => n510, Q => 
                           REGISTERS_14_4_port, QN => n_1507);
   REGISTERS_reg_14_3_inst : DFF_X1 port map( D => n2106, CK => n510, Q => 
                           REGISTERS_14_3_port, QN => n_1508);
   REGISTERS_reg_14_2_inst : DFF_X1 port map( D => n2105, CK => n510, Q => 
                           REGISTERS_14_2_port, QN => n_1509);
   REGISTERS_reg_14_1_inst : DFF_X1 port map( D => n2104, CK => n510, Q => 
                           REGISTERS_14_1_port, QN => n_1510);
   REGISTERS_reg_14_0_inst : DFF_X1 port map( D => n2103, CK => n510, Q => 
                           REGISTERS_14_0_port, QN => n_1511);
   REGISTERS_reg_15_31_inst : DFF_X1 port map( D => n2102, CK => n511, Q => 
                           REGISTERS_15_31_port, QN => n_1512);
   REGISTERS_reg_15_30_inst : DFF_X1 port map( D => n2101, CK => n511, Q => 
                           REGISTERS_15_30_port, QN => n_1513);
   REGISTERS_reg_15_29_inst : DFF_X1 port map( D => n2100, CK => n511, Q => 
                           REGISTERS_15_29_port, QN => n_1514);
   REGISTERS_reg_15_28_inst : DFF_X1 port map( D => n2099, CK => n511, Q => 
                           REGISTERS_15_28_port, QN => n_1515);
   REGISTERS_reg_15_27_inst : DFF_X1 port map( D => n2098, CK => n511, Q => 
                           REGISTERS_15_27_port, QN => n_1516);
   REGISTERS_reg_15_26_inst : DFF_X1 port map( D => n2097, CK => n511, Q => 
                           REGISTERS_15_26_port, QN => n_1517);
   REGISTERS_reg_15_25_inst : DFF_X1 port map( D => n2096, CK => n511, Q => 
                           REGISTERS_15_25_port, QN => n_1518);
   REGISTERS_reg_15_24_inst : DFF_X1 port map( D => n2095, CK => n511, Q => 
                           REGISTERS_15_24_port, QN => n_1519);
   REGISTERS_reg_15_23_inst : DFF_X1 port map( D => n2094, CK => n511, Q => 
                           REGISTERS_15_23_port, QN => n_1520);
   REGISTERS_reg_15_22_inst : DFF_X1 port map( D => n2093, CK => n511, Q => 
                           REGISTERS_15_22_port, QN => n_1521);
   REGISTERS_reg_15_21_inst : DFF_X1 port map( D => n2092, CK => n511, Q => 
                           REGISTERS_15_21_port, QN => n_1522);
   REGISTERS_reg_15_20_inst : DFF_X1 port map( D => n2091, CK => n512, Q => 
                           REGISTERS_15_20_port, QN => n_1523);
   REGISTERS_reg_15_19_inst : DFF_X1 port map( D => n2090, CK => n512, Q => 
                           REGISTERS_15_19_port, QN => n_1524);
   REGISTERS_reg_15_18_inst : DFF_X1 port map( D => n2089, CK => n512, Q => 
                           REGISTERS_15_18_port, QN => n_1525);
   REGISTERS_reg_15_17_inst : DFF_X1 port map( D => n2088, CK => n512, Q => 
                           REGISTERS_15_17_port, QN => n_1526);
   REGISTERS_reg_15_16_inst : DFF_X1 port map( D => n2087, CK => n512, Q => 
                           REGISTERS_15_16_port, QN => n_1527);
   REGISTERS_reg_15_15_inst : DFF_X1 port map( D => n2086, CK => n512, Q => 
                           REGISTERS_15_15_port, QN => n_1528);
   REGISTERS_reg_15_14_inst : DFF_X1 port map( D => n2085, CK => n512, Q => 
                           REGISTERS_15_14_port, QN => n_1529);
   REGISTERS_reg_15_13_inst : DFF_X1 port map( D => n2084, CK => n512, Q => 
                           REGISTERS_15_13_port, QN => n_1530);
   REGISTERS_reg_15_12_inst : DFF_X1 port map( D => n2083, CK => n512, Q => 
                           REGISTERS_15_12_port, QN => n_1531);
   REGISTERS_reg_15_11_inst : DFF_X1 port map( D => n2082, CK => n512, Q => 
                           REGISTERS_15_11_port, QN => n_1532);
   REGISTERS_reg_15_10_inst : DFF_X1 port map( D => n2081, CK => n512, Q => 
                           REGISTERS_15_10_port, QN => n_1533);
   REGISTERS_reg_15_9_inst : DFF_X1 port map( D => n2080, CK => n513, Q => 
                           REGISTERS_15_9_port, QN => n_1534);
   REGISTERS_reg_15_8_inst : DFF_X1 port map( D => n2079, CK => n513, Q => 
                           REGISTERS_15_8_port, QN => n_1535);
   REGISTERS_reg_15_7_inst : DFF_X1 port map( D => n2078, CK => n513, Q => 
                           REGISTERS_15_7_port, QN => n_1536);
   REGISTERS_reg_15_6_inst : DFF_X1 port map( D => n2077, CK => n513, Q => 
                           REGISTERS_15_6_port, QN => n_1537);
   REGISTERS_reg_15_5_inst : DFF_X1 port map( D => n2076, CK => n513, Q => 
                           REGISTERS_15_5_port, QN => n_1538);
   REGISTERS_reg_15_4_inst : DFF_X1 port map( D => n2075, CK => n513, Q => 
                           REGISTERS_15_4_port, QN => n_1539);
   REGISTERS_reg_15_3_inst : DFF_X1 port map( D => n2074, CK => n513, Q => 
                           REGISTERS_15_3_port, QN => n_1540);
   REGISTERS_reg_15_2_inst : DFF_X1 port map( D => n2073, CK => n513, Q => 
                           REGISTERS_15_2_port, QN => n_1541);
   REGISTERS_reg_15_1_inst : DFF_X1 port map( D => n2072, CK => n513, Q => 
                           REGISTERS_15_1_port, QN => n_1542);
   REGISTERS_reg_15_0_inst : DFF_X1 port map( D => n2071, CK => n513, Q => 
                           REGISTERS_15_0_port, QN => n_1543);
   REGISTERS_reg_16_31_inst : DFF_X1 port map( D => n2070, CK => n444, Q => 
                           REGISTERS_16_31_port, QN => n_1544);
   REGISTERS_reg_16_30_inst : DFF_X1 port map( D => n2069, CK => n444, Q => 
                           REGISTERS_16_30_port, QN => n_1545);
   REGISTERS_reg_16_29_inst : DFF_X1 port map( D => n2068, CK => n444, Q => 
                           REGISTERS_16_29_port, QN => n_1546);
   REGISTERS_reg_16_28_inst : DFF_X1 port map( D => n2067, CK => n444, Q => 
                           REGISTERS_16_28_port, QN => n_1547);
   REGISTERS_reg_16_27_inst : DFF_X1 port map( D => n2066, CK => n444, Q => 
                           REGISTERS_16_27_port, QN => n_1548);
   REGISTERS_reg_16_26_inst : DFF_X1 port map( D => n2065, CK => n444, Q => 
                           REGISTERS_16_26_port, QN => n_1549);
   REGISTERS_reg_16_25_inst : DFF_X1 port map( D => n2064, CK => n444, Q => 
                           REGISTERS_16_25_port, QN => n_1550);
   REGISTERS_reg_16_24_inst : DFF_X1 port map( D => n2063, CK => n444, Q => 
                           REGISTERS_16_24_port, QN => n_1551);
   REGISTERS_reg_16_23_inst : DFF_X1 port map( D => n2062, CK => n444, Q => 
                           REGISTERS_16_23_port, QN => n_1552);
   REGISTERS_reg_16_22_inst : DFF_X1 port map( D => n2061, CK => n444, Q => 
                           REGISTERS_16_22_port, QN => n_1553);
   REGISTERS_reg_16_21_inst : DFF_X1 port map( D => n2060, CK => n445, Q => 
                           REGISTERS_16_21_port, QN => n_1554);
   REGISTERS_reg_16_20_inst : DFF_X1 port map( D => n2059, CK => n445, Q => 
                           REGISTERS_16_20_port, QN => n_1555);
   REGISTERS_reg_16_19_inst : DFF_X1 port map( D => n2058, CK => n445, Q => 
                           REGISTERS_16_19_port, QN => n_1556);
   REGISTERS_reg_16_18_inst : DFF_X1 port map( D => n2057, CK => n445, Q => 
                           REGISTERS_16_18_port, QN => n_1557);
   REGISTERS_reg_16_17_inst : DFF_X1 port map( D => n2056, CK => n445, Q => 
                           REGISTERS_16_17_port, QN => n_1558);
   REGISTERS_reg_16_16_inst : DFF_X1 port map( D => n2055, CK => n445, Q => 
                           REGISTERS_16_16_port, QN => n_1559);
   REGISTERS_reg_16_15_inst : DFF_X1 port map( D => n2054, CK => n445, Q => 
                           REGISTERS_16_15_port, QN => n_1560);
   REGISTERS_reg_16_14_inst : DFF_X1 port map( D => n2053, CK => n445, Q => 
                           REGISTERS_16_14_port, QN => n_1561);
   REGISTERS_reg_16_13_inst : DFF_X1 port map( D => n2052, CK => n445, Q => 
                           REGISTERS_16_13_port, QN => n_1562);
   REGISTERS_reg_16_12_inst : DFF_X1 port map( D => n2051, CK => n445, Q => 
                           REGISTERS_16_12_port, QN => n_1563);
   REGISTERS_reg_16_11_inst : DFF_X1 port map( D => n2050, CK => n445, Q => 
                           REGISTERS_16_11_port, QN => n_1564);
   REGISTERS_reg_16_10_inst : DFF_X1 port map( D => n2049, CK => n446, Q => 
                           REGISTERS_16_10_port, QN => n_1565);
   REGISTERS_reg_16_9_inst : DFF_X1 port map( D => n2048, CK => n446, Q => 
                           REGISTERS_16_9_port, QN => n_1566);
   REGISTERS_reg_16_8_inst : DFF_X1 port map( D => n2047, CK => n446, Q => 
                           REGISTERS_16_8_port, QN => n_1567);
   REGISTERS_reg_16_7_inst : DFF_X1 port map( D => n2046, CK => n446, Q => 
                           REGISTERS_16_7_port, QN => n_1568);
   REGISTERS_reg_16_6_inst : DFF_X1 port map( D => n2045, CK => n446, Q => 
                           REGISTERS_16_6_port, QN => n_1569);
   REGISTERS_reg_16_5_inst : DFF_X1 port map( D => n2044, CK => n446, Q => 
                           REGISTERS_16_5_port, QN => n_1570);
   REGISTERS_reg_16_4_inst : DFF_X1 port map( D => n2043, CK => n446, Q => 
                           REGISTERS_16_4_port, QN => n_1571);
   REGISTERS_reg_16_3_inst : DFF_X1 port map( D => n2042, CK => n446, Q => 
                           REGISTERS_16_3_port, QN => n_1572);
   REGISTERS_reg_16_2_inst : DFF_X1 port map( D => n2041, CK => n446, Q => 
                           REGISTERS_16_2_port, QN => n_1573);
   REGISTERS_reg_16_1_inst : DFF_X1 port map( D => n2040, CK => n446, Q => 
                           REGISTERS_16_1_port, QN => n_1574);
   REGISTERS_reg_16_0_inst : DFF_X1 port map( D => n2039, CK => n446, Q => 
                           REGISTERS_16_0_port, QN => n_1575);
   REGISTERS_reg_17_31_inst : DFF_X1 port map( D => n2038, CK => n447, Q => 
                           REGISTERS_17_31_port, QN => n_1576);
   REGISTERS_reg_17_30_inst : DFF_X1 port map( D => n2037, CK => n447, Q => 
                           REGISTERS_17_30_port, QN => n_1577);
   REGISTERS_reg_17_29_inst : DFF_X1 port map( D => n2036, CK => n447, Q => 
                           REGISTERS_17_29_port, QN => n_1578);
   REGISTERS_reg_17_28_inst : DFF_X1 port map( D => n2035, CK => n447, Q => 
                           REGISTERS_17_28_port, QN => n_1579);
   REGISTERS_reg_17_27_inst : DFF_X1 port map( D => n2034, CK => n447, Q => 
                           REGISTERS_17_27_port, QN => n_1580);
   REGISTERS_reg_17_26_inst : DFF_X1 port map( D => n2033, CK => n447, Q => 
                           REGISTERS_17_26_port, QN => n_1581);
   REGISTERS_reg_17_25_inst : DFF_X1 port map( D => n2032, CK => n447, Q => 
                           REGISTERS_17_25_port, QN => n_1582);
   REGISTERS_reg_17_24_inst : DFF_X1 port map( D => n2031, CK => n447, Q => 
                           REGISTERS_17_24_port, QN => n_1583);
   REGISTERS_reg_17_23_inst : DFF_X1 port map( D => n2030, CK => n447, Q => 
                           REGISTERS_17_23_port, QN => n_1584);
   REGISTERS_reg_17_22_inst : DFF_X1 port map( D => n2029, CK => n447, Q => 
                           REGISTERS_17_22_port, QN => n_1585);
   REGISTERS_reg_17_21_inst : DFF_X1 port map( D => n2028, CK => n447, Q => 
                           REGISTERS_17_21_port, QN => n_1586);
   REGISTERS_reg_17_20_inst : DFF_X1 port map( D => n2027, CK => n448, Q => 
                           REGISTERS_17_20_port, QN => n_1587);
   REGISTERS_reg_17_19_inst : DFF_X1 port map( D => n2026, CK => n448, Q => 
                           REGISTERS_17_19_port, QN => n_1588);
   REGISTERS_reg_17_18_inst : DFF_X1 port map( D => n2025, CK => n448, Q => 
                           REGISTERS_17_18_port, QN => n_1589);
   REGISTERS_reg_17_17_inst : DFF_X1 port map( D => n2024, CK => n448, Q => 
                           REGISTERS_17_17_port, QN => n_1590);
   REGISTERS_reg_17_16_inst : DFF_X1 port map( D => n2023, CK => n448, Q => 
                           REGISTERS_17_16_port, QN => n_1591);
   REGISTERS_reg_17_15_inst : DFF_X1 port map( D => n2022, CK => n448, Q => 
                           REGISTERS_17_15_port, QN => n_1592);
   REGISTERS_reg_17_14_inst : DFF_X1 port map( D => n2021, CK => n448, Q => 
                           REGISTERS_17_14_port, QN => n_1593);
   REGISTERS_reg_17_13_inst : DFF_X1 port map( D => n2020, CK => n448, Q => 
                           REGISTERS_17_13_port, QN => n_1594);
   REGISTERS_reg_17_12_inst : DFF_X1 port map( D => n2019, CK => n448, Q => 
                           REGISTERS_17_12_port, QN => n_1595);
   REGISTERS_reg_17_11_inst : DFF_X1 port map( D => n2018, CK => n448, Q => 
                           REGISTERS_17_11_port, QN => n_1596);
   REGISTERS_reg_17_10_inst : DFF_X1 port map( D => n2017, CK => n448, Q => 
                           REGISTERS_17_10_port, QN => n_1597);
   REGISTERS_reg_17_9_inst : DFF_X1 port map( D => n2016, CK => n449, Q => 
                           REGISTERS_17_9_port, QN => n_1598);
   REGISTERS_reg_17_8_inst : DFF_X1 port map( D => n2015, CK => n449, Q => 
                           REGISTERS_17_8_port, QN => n_1599);
   REGISTERS_reg_17_7_inst : DFF_X1 port map( D => n2014, CK => n449, Q => 
                           REGISTERS_17_7_port, QN => n_1600);
   REGISTERS_reg_17_6_inst : DFF_X1 port map( D => n2013, CK => n449, Q => 
                           REGISTERS_17_6_port, QN => n_1601);
   REGISTERS_reg_17_5_inst : DFF_X1 port map( D => n2012, CK => n449, Q => 
                           REGISTERS_17_5_port, QN => n_1602);
   REGISTERS_reg_17_4_inst : DFF_X1 port map( D => n2011, CK => n449, Q => 
                           REGISTERS_17_4_port, QN => n_1603);
   REGISTERS_reg_17_3_inst : DFF_X1 port map( D => n2010, CK => n449, Q => 
                           REGISTERS_17_3_port, QN => n_1604);
   REGISTERS_reg_17_2_inst : DFF_X1 port map( D => n2009, CK => n449, Q => 
                           REGISTERS_17_2_port, QN => n_1605);
   REGISTERS_reg_17_1_inst : DFF_X1 port map( D => n2008, CK => n449, Q => 
                           REGISTERS_17_1_port, QN => n_1606);
   REGISTERS_reg_17_0_inst : DFF_X1 port map( D => n2007, CK => n449, Q => 
                           REGISTERS_17_0_port, QN => n_1607);
   REGISTERS_reg_18_31_inst : DFF_X1 port map( D => n2006, CK => n449, Q => 
                           REGISTERS_18_31_port, QN => n_1608);
   REGISTERS_reg_18_30_inst : DFF_X1 port map( D => n2005, CK => n450, Q => 
                           REGISTERS_18_30_port, QN => n_1609);
   REGISTERS_reg_18_29_inst : DFF_X1 port map( D => n2004, CK => n450, Q => 
                           REGISTERS_18_29_port, QN => n_1610);
   REGISTERS_reg_18_28_inst : DFF_X1 port map( D => n2003, CK => n450, Q => 
                           REGISTERS_18_28_port, QN => n_1611);
   REGISTERS_reg_18_27_inst : DFF_X1 port map( D => n2002, CK => n450, Q => 
                           REGISTERS_18_27_port, QN => n_1612);
   REGISTERS_reg_18_26_inst : DFF_X1 port map( D => n2001, CK => n450, Q => 
                           REGISTERS_18_26_port, QN => n_1613);
   REGISTERS_reg_18_25_inst : DFF_X1 port map( D => n2000, CK => n450, Q => 
                           REGISTERS_18_25_port, QN => n_1614);
   REGISTERS_reg_18_24_inst : DFF_X1 port map( D => n1999, CK => n450, Q => 
                           REGISTERS_18_24_port, QN => n_1615);
   REGISTERS_reg_18_23_inst : DFF_X1 port map( D => n1998, CK => n450, Q => 
                           REGISTERS_18_23_port, QN => n_1616);
   REGISTERS_reg_18_22_inst : DFF_X1 port map( D => n1997, CK => n450, Q => 
                           REGISTERS_18_22_port, QN => n_1617);
   REGISTERS_reg_18_21_inst : DFF_X1 port map( D => n1996, CK => n450, Q => 
                           REGISTERS_18_21_port, QN => n_1618);
   REGISTERS_reg_18_20_inst : DFF_X1 port map( D => n1995, CK => n450, Q => 
                           REGISTERS_18_20_port, QN => n_1619);
   REGISTERS_reg_18_19_inst : DFF_X1 port map( D => n1994, CK => n451, Q => 
                           REGISTERS_18_19_port, QN => n_1620);
   REGISTERS_reg_18_18_inst : DFF_X1 port map( D => n1993, CK => n451, Q => 
                           REGISTERS_18_18_port, QN => n_1621);
   REGISTERS_reg_18_17_inst : DFF_X1 port map( D => n1992, CK => n451, Q => 
                           REGISTERS_18_17_port, QN => n_1622);
   REGISTERS_reg_18_16_inst : DFF_X1 port map( D => n1991, CK => n451, Q => 
                           REGISTERS_18_16_port, QN => n_1623);
   REGISTERS_reg_18_15_inst : DFF_X1 port map( D => n1990, CK => n451, Q => 
                           REGISTERS_18_15_port, QN => n_1624);
   REGISTERS_reg_18_14_inst : DFF_X1 port map( D => n1989, CK => n451, Q => 
                           REGISTERS_18_14_port, QN => n_1625);
   REGISTERS_reg_18_13_inst : DFF_X1 port map( D => n1988, CK => n451, Q => 
                           REGISTERS_18_13_port, QN => n_1626);
   REGISTERS_reg_18_12_inst : DFF_X1 port map( D => n1987, CK => n451, Q => 
                           REGISTERS_18_12_port, QN => n_1627);
   REGISTERS_reg_18_11_inst : DFF_X1 port map( D => n1986, CK => n451, Q => 
                           REGISTERS_18_11_port, QN => n_1628);
   REGISTERS_reg_18_10_inst : DFF_X1 port map( D => n1985, CK => n451, Q => 
                           REGISTERS_18_10_port, QN => n_1629);
   REGISTERS_reg_18_9_inst : DFF_X1 port map( D => n1984, CK => n451, Q => 
                           REGISTERS_18_9_port, QN => n_1630);
   REGISTERS_reg_18_8_inst : DFF_X1 port map( D => n1983, CK => n452, Q => 
                           REGISTERS_18_8_port, QN => n_1631);
   REGISTERS_reg_18_7_inst : DFF_X1 port map( D => n1982, CK => n452, Q => 
                           REGISTERS_18_7_port, QN => n_1632);
   REGISTERS_reg_18_6_inst : DFF_X1 port map( D => n1981, CK => n452, Q => 
                           REGISTERS_18_6_port, QN => n_1633);
   REGISTERS_reg_18_5_inst : DFF_X1 port map( D => n1980, CK => n452, Q => 
                           REGISTERS_18_5_port, QN => n_1634);
   REGISTERS_reg_18_4_inst : DFF_X1 port map( D => n1979, CK => n452, Q => 
                           REGISTERS_18_4_port, QN => n_1635);
   REGISTERS_reg_18_3_inst : DFF_X1 port map( D => n1978, CK => n452, Q => 
                           REGISTERS_18_3_port, QN => n_1636);
   REGISTERS_reg_18_2_inst : DFF_X1 port map( D => n1977, CK => n452, Q => 
                           REGISTERS_18_2_port, QN => n_1637);
   REGISTERS_reg_18_1_inst : DFF_X1 port map( D => n1976, CK => n452, Q => 
                           REGISTERS_18_1_port, QN => n_1638);
   REGISTERS_reg_18_0_inst : DFF_X1 port map( D => n1975, CK => n452, Q => 
                           REGISTERS_18_0_port, QN => n_1639);
   REGISTERS_reg_19_31_inst : DFF_X1 port map( D => n1974, CK => n452, Q => 
                           REGISTERS_19_31_port, QN => n_1640);
   REGISTERS_reg_19_30_inst : DFF_X1 port map( D => n1973, CK => n452, Q => 
                           REGISTERS_19_30_port, QN => n_1641);
   REGISTERS_reg_19_29_inst : DFF_X1 port map( D => n1972, CK => n453, Q => 
                           REGISTERS_19_29_port, QN => n_1642);
   REGISTERS_reg_19_28_inst : DFF_X1 port map( D => n1971, CK => n453, Q => 
                           REGISTERS_19_28_port, QN => n_1643);
   REGISTERS_reg_19_27_inst : DFF_X1 port map( D => n1970, CK => n453, Q => 
                           REGISTERS_19_27_port, QN => n_1644);
   REGISTERS_reg_19_26_inst : DFF_X1 port map( D => n1969, CK => n453, Q => 
                           REGISTERS_19_26_port, QN => n_1645);
   REGISTERS_reg_19_25_inst : DFF_X1 port map( D => n1968, CK => n453, Q => 
                           REGISTERS_19_25_port, QN => n_1646);
   REGISTERS_reg_19_24_inst : DFF_X1 port map( D => n1967, CK => n453, Q => 
                           REGISTERS_19_24_port, QN => n_1647);
   REGISTERS_reg_19_23_inst : DFF_X1 port map( D => n1966, CK => n453, Q => 
                           REGISTERS_19_23_port, QN => n_1648);
   REGISTERS_reg_19_22_inst : DFF_X1 port map( D => n1965, CK => n453, Q => 
                           REGISTERS_19_22_port, QN => n_1649);
   REGISTERS_reg_19_21_inst : DFF_X1 port map( D => n1964, CK => n453, Q => 
                           REGISTERS_19_21_port, QN => n_1650);
   REGISTERS_reg_19_20_inst : DFF_X1 port map( D => n1963, CK => n453, Q => 
                           REGISTERS_19_20_port, QN => n_1651);
   REGISTERS_reg_19_19_inst : DFF_X1 port map( D => n1962, CK => n453, Q => 
                           REGISTERS_19_19_port, QN => n_1652);
   REGISTERS_reg_19_18_inst : DFF_X1 port map( D => n1961, CK => n454, Q => 
                           REGISTERS_19_18_port, QN => n_1653);
   REGISTERS_reg_19_17_inst : DFF_X1 port map( D => n1960, CK => n454, Q => 
                           REGISTERS_19_17_port, QN => n_1654);
   REGISTERS_reg_19_16_inst : DFF_X1 port map( D => n1959, CK => n454, Q => 
                           REGISTERS_19_16_port, QN => n_1655);
   REGISTERS_reg_19_15_inst : DFF_X1 port map( D => n1958, CK => n454, Q => 
                           REGISTERS_19_15_port, QN => n_1656);
   REGISTERS_reg_19_14_inst : DFF_X1 port map( D => n1957, CK => n454, Q => 
                           REGISTERS_19_14_port, QN => n_1657);
   REGISTERS_reg_19_13_inst : DFF_X1 port map( D => n1956, CK => n454, Q => 
                           REGISTERS_19_13_port, QN => n_1658);
   REGISTERS_reg_19_12_inst : DFF_X1 port map( D => n1955, CK => n454, Q => 
                           REGISTERS_19_12_port, QN => n_1659);
   REGISTERS_reg_19_11_inst : DFF_X1 port map( D => n1954, CK => n454, Q => 
                           REGISTERS_19_11_port, QN => n_1660);
   REGISTERS_reg_19_10_inst : DFF_X1 port map( D => n1953, CK => n454, Q => 
                           REGISTERS_19_10_port, QN => n_1661);
   REGISTERS_reg_19_9_inst : DFF_X1 port map( D => n1952, CK => n454, Q => 
                           REGISTERS_19_9_port, QN => n_1662);
   REGISTERS_reg_19_8_inst : DFF_X1 port map( D => n1951, CK => n454, Q => 
                           REGISTERS_19_8_port, QN => n_1663);
   REGISTERS_reg_19_7_inst : DFF_X1 port map( D => n1950, CK => n455, Q => 
                           REGISTERS_19_7_port, QN => n_1664);
   REGISTERS_reg_19_6_inst : DFF_X1 port map( D => n1949, CK => n455, Q => 
                           REGISTERS_19_6_port, QN => n_1665);
   REGISTERS_reg_19_5_inst : DFF_X1 port map( D => n1948, CK => n455, Q => 
                           REGISTERS_19_5_port, QN => n_1666);
   REGISTERS_reg_19_4_inst : DFF_X1 port map( D => n1947, CK => n455, Q => 
                           REGISTERS_19_4_port, QN => n_1667);
   REGISTERS_reg_19_3_inst : DFF_X1 port map( D => n1946, CK => n455, Q => 
                           REGISTERS_19_3_port, QN => n_1668);
   REGISTERS_reg_19_2_inst : DFF_X1 port map( D => n1945, CK => n455, Q => 
                           REGISTERS_19_2_port, QN => n_1669);
   REGISTERS_reg_19_1_inst : DFF_X1 port map( D => n1944, CK => n455, Q => 
                           REGISTERS_19_1_port, QN => n_1670);
   REGISTERS_reg_19_0_inst : DFF_X1 port map( D => n1943, CK => n455, Q => 
                           REGISTERS_19_0_port, QN => n_1671);
   REGISTERS_reg_20_31_inst : DFF_X1 port map( D => n1942, CK => n455, Q => 
                           REGISTERS_20_31_port, QN => n_1672);
   REGISTERS_reg_20_30_inst : DFF_X1 port map( D => n1941, CK => n455, Q => 
                           REGISTERS_20_30_port, QN => n_1673);
   REGISTERS_reg_20_29_inst : DFF_X1 port map( D => n1940, CK => n455, Q => 
                           REGISTERS_20_29_port, QN => n_1674);
   REGISTERS_reg_20_28_inst : DFF_X1 port map( D => n1939, CK => n456, Q => 
                           REGISTERS_20_28_port, QN => n_1675);
   REGISTERS_reg_20_27_inst : DFF_X1 port map( D => n1938, CK => n456, Q => 
                           REGISTERS_20_27_port, QN => n_1676);
   REGISTERS_reg_20_26_inst : DFF_X1 port map( D => n1937, CK => n456, Q => 
                           REGISTERS_20_26_port, QN => n_1677);
   REGISTERS_reg_20_25_inst : DFF_X1 port map( D => n1936, CK => n456, Q => 
                           REGISTERS_20_25_port, QN => n_1678);
   REGISTERS_reg_20_24_inst : DFF_X1 port map( D => n1935, CK => n456, Q => 
                           REGISTERS_20_24_port, QN => n_1679);
   REGISTERS_reg_20_23_inst : DFF_X1 port map( D => n1934, CK => n456, Q => 
                           REGISTERS_20_23_port, QN => n_1680);
   REGISTERS_reg_20_22_inst : DFF_X1 port map( D => n1933, CK => n456, Q => 
                           REGISTERS_20_22_port, QN => n_1681);
   REGISTERS_reg_20_21_inst : DFF_X1 port map( D => n1932, CK => n456, Q => 
                           REGISTERS_20_21_port, QN => n_1682);
   REGISTERS_reg_20_20_inst : DFF_X1 port map( D => n1931, CK => n456, Q => 
                           REGISTERS_20_20_port, QN => n_1683);
   REGISTERS_reg_20_19_inst : DFF_X1 port map( D => n1930, CK => n456, Q => 
                           REGISTERS_20_19_port, QN => n_1684);
   REGISTERS_reg_20_18_inst : DFF_X1 port map( D => n1929, CK => n456, Q => 
                           REGISTERS_20_18_port, QN => n_1685);
   REGISTERS_reg_20_17_inst : DFF_X1 port map( D => n1928, CK => n457, Q => 
                           REGISTERS_20_17_port, QN => n_1686);
   REGISTERS_reg_20_16_inst : DFF_X1 port map( D => n1927, CK => n457, Q => 
                           REGISTERS_20_16_port, QN => n_1687);
   REGISTERS_reg_20_15_inst : DFF_X1 port map( D => n1926, CK => n457, Q => 
                           REGISTERS_20_15_port, QN => n_1688);
   REGISTERS_reg_20_14_inst : DFF_X1 port map( D => n1925, CK => n457, Q => 
                           REGISTERS_20_14_port, QN => n_1689);
   REGISTERS_reg_20_13_inst : DFF_X1 port map( D => n1924, CK => n457, Q => 
                           REGISTERS_20_13_port, QN => n_1690);
   REGISTERS_reg_20_12_inst : DFF_X1 port map( D => n1923, CK => n457, Q => 
                           REGISTERS_20_12_port, QN => n_1691);
   REGISTERS_reg_20_11_inst : DFF_X1 port map( D => n1922, CK => n457, Q => 
                           REGISTERS_20_11_port, QN => n_1692);
   REGISTERS_reg_20_10_inst : DFF_X1 port map( D => n1921, CK => n457, Q => 
                           REGISTERS_20_10_port, QN => n_1693);
   REGISTERS_reg_20_9_inst : DFF_X1 port map( D => n1920, CK => n457, Q => 
                           REGISTERS_20_9_port, QN => n_1694);
   REGISTERS_reg_20_8_inst : DFF_X1 port map( D => n1919, CK => n457, Q => 
                           REGISTERS_20_8_port, QN => n_1695);
   REGISTERS_reg_20_7_inst : DFF_X1 port map( D => n1918, CK => n457, Q => 
                           REGISTERS_20_7_port, QN => n_1696);
   REGISTERS_reg_20_6_inst : DFF_X1 port map( D => n1917, CK => n458, Q => 
                           REGISTERS_20_6_port, QN => n_1697);
   REGISTERS_reg_20_5_inst : DFF_X1 port map( D => n1916, CK => n458, Q => 
                           REGISTERS_20_5_port, QN => n_1698);
   REGISTERS_reg_20_4_inst : DFF_X1 port map( D => n1915, CK => n458, Q => 
                           REGISTERS_20_4_port, QN => n_1699);
   REGISTERS_reg_20_3_inst : DFF_X1 port map( D => n1914, CK => n458, Q => 
                           REGISTERS_20_3_port, QN => n_1700);
   REGISTERS_reg_20_2_inst : DFF_X1 port map( D => n1913, CK => n458, Q => 
                           REGISTERS_20_2_port, QN => n_1701);
   REGISTERS_reg_20_1_inst : DFF_X1 port map( D => n1912, CK => n458, Q => 
                           REGISTERS_20_1_port, QN => n_1702);
   REGISTERS_reg_20_0_inst : DFF_X1 port map( D => n1911, CK => n458, Q => 
                           REGISTERS_20_0_port, QN => n_1703);
   REGISTERS_reg_21_31_inst : DFF_X1 port map( D => n1910, CK => n458, Q => 
                           REGISTERS_21_31_port, QN => n_1704);
   REGISTERS_reg_21_30_inst : DFF_X1 port map( D => n1909, CK => n458, Q => 
                           REGISTERS_21_30_port, QN => n_1705);
   REGISTERS_reg_21_29_inst : DFF_X1 port map( D => n1908, CK => n458, Q => 
                           REGISTERS_21_29_port, QN => n_1706);
   REGISTERS_reg_21_28_inst : DFF_X1 port map( D => n1907, CK => n458, Q => 
                           REGISTERS_21_28_port, QN => n_1707);
   REGISTERS_reg_21_27_inst : DFF_X1 port map( D => n1906, CK => n459, Q => 
                           REGISTERS_21_27_port, QN => n_1708);
   REGISTERS_reg_21_26_inst : DFF_X1 port map( D => n1905, CK => n459, Q => 
                           REGISTERS_21_26_port, QN => n_1709);
   REGISTERS_reg_21_25_inst : DFF_X1 port map( D => n1904, CK => n459, Q => 
                           REGISTERS_21_25_port, QN => n_1710);
   REGISTERS_reg_21_24_inst : DFF_X1 port map( D => n1903, CK => n459, Q => 
                           REGISTERS_21_24_port, QN => n_1711);
   REGISTERS_reg_21_23_inst : DFF_X1 port map( D => n1902, CK => n459, Q => 
                           REGISTERS_21_23_port, QN => n_1712);
   REGISTERS_reg_21_22_inst : DFF_X1 port map( D => n1901, CK => n459, Q => 
                           REGISTERS_21_22_port, QN => n_1713);
   REGISTERS_reg_21_21_inst : DFF_X1 port map( D => n1900, CK => n459, Q => 
                           REGISTERS_21_21_port, QN => n_1714);
   REGISTERS_reg_21_20_inst : DFF_X1 port map( D => n1899, CK => n459, Q => 
                           REGISTERS_21_20_port, QN => n_1715);
   REGISTERS_reg_21_19_inst : DFF_X1 port map( D => n1898, CK => n459, Q => 
                           REGISTERS_21_19_port, QN => n_1716);
   REGISTERS_reg_21_18_inst : DFF_X1 port map( D => n1897, CK => n459, Q => 
                           REGISTERS_21_18_port, QN => n_1717);
   REGISTERS_reg_21_17_inst : DFF_X1 port map( D => n1896, CK => n459, Q => 
                           REGISTERS_21_17_port, QN => n_1718);
   REGISTERS_reg_21_16_inst : DFF_X1 port map( D => n1895, CK => n460, Q => 
                           REGISTERS_21_16_port, QN => n_1719);
   REGISTERS_reg_21_15_inst : DFF_X1 port map( D => n1894, CK => n460, Q => 
                           REGISTERS_21_15_port, QN => n_1720);
   REGISTERS_reg_21_14_inst : DFF_X1 port map( D => n1893, CK => n460, Q => 
                           REGISTERS_21_14_port, QN => n_1721);
   REGISTERS_reg_21_13_inst : DFF_X1 port map( D => n1892, CK => n460, Q => 
                           REGISTERS_21_13_port, QN => n_1722);
   REGISTERS_reg_21_12_inst : DFF_X1 port map( D => n1891, CK => n460, Q => 
                           REGISTERS_21_12_port, QN => n_1723);
   REGISTERS_reg_21_11_inst : DFF_X1 port map( D => n1890, CK => n460, Q => 
                           REGISTERS_21_11_port, QN => n_1724);
   REGISTERS_reg_21_10_inst : DFF_X1 port map( D => n1889, CK => n460, Q => 
                           REGISTERS_21_10_port, QN => n_1725);
   REGISTERS_reg_21_9_inst : DFF_X1 port map( D => n1888, CK => n460, Q => 
                           REGISTERS_21_9_port, QN => n_1726);
   REGISTERS_reg_21_8_inst : DFF_X1 port map( D => n1887, CK => n460, Q => 
                           REGISTERS_21_8_port, QN => n_1727);
   REGISTERS_reg_21_7_inst : DFF_X1 port map( D => n1886, CK => n460, Q => 
                           REGISTERS_21_7_port, QN => n_1728);
   REGISTERS_reg_21_6_inst : DFF_X1 port map( D => n1885, CK => n460, Q => 
                           REGISTERS_21_6_port, QN => n_1729);
   REGISTERS_reg_21_5_inst : DFF_X1 port map( D => n1884, CK => n461, Q => 
                           REGISTERS_21_5_port, QN => n_1730);
   REGISTERS_reg_21_4_inst : DFF_X1 port map( D => n1883, CK => n461, Q => 
                           REGISTERS_21_4_port, QN => n_1731);
   REGISTERS_reg_21_3_inst : DFF_X1 port map( D => n1882, CK => n461, Q => 
                           REGISTERS_21_3_port, QN => n_1732);
   REGISTERS_reg_21_2_inst : DFF_X1 port map( D => n1881, CK => n461, Q => 
                           REGISTERS_21_2_port, QN => n_1733);
   REGISTERS_reg_21_1_inst : DFF_X1 port map( D => n1880, CK => n461, Q => 
                           REGISTERS_21_1_port, QN => n_1734);
   REGISTERS_reg_21_0_inst : DFF_X1 port map( D => n1879, CK => n461, Q => 
                           REGISTERS_21_0_port, QN => n_1735);
   REGISTERS_reg_22_31_inst : DFF_X1 port map( D => n1878, CK => n461, Q => 
                           REGISTERS_22_31_port, QN => n_1736);
   REGISTERS_reg_22_30_inst : DFF_X1 port map( D => n1877, CK => n461, Q => 
                           REGISTERS_22_30_port, QN => n_1737);
   REGISTERS_reg_22_29_inst : DFF_X1 port map( D => n1876, CK => n461, Q => 
                           REGISTERS_22_29_port, QN => n_1738);
   REGISTERS_reg_22_28_inst : DFF_X1 port map( D => n1875, CK => n461, Q => 
                           REGISTERS_22_28_port, QN => n_1739);
   REGISTERS_reg_22_27_inst : DFF_X1 port map( D => n1874, CK => n461, Q => 
                           REGISTERS_22_27_port, QN => n_1740);
   REGISTERS_reg_22_26_inst : DFF_X1 port map( D => n1873, CK => n462, Q => 
                           REGISTERS_22_26_port, QN => n_1741);
   REGISTERS_reg_22_25_inst : DFF_X1 port map( D => n1872, CK => n462, Q => 
                           REGISTERS_22_25_port, QN => n_1742);
   REGISTERS_reg_22_24_inst : DFF_X1 port map( D => n1871, CK => n462, Q => 
                           REGISTERS_22_24_port, QN => n_1743);
   REGISTERS_reg_22_23_inst : DFF_X1 port map( D => n1870, CK => n462, Q => 
                           REGISTERS_22_23_port, QN => n_1744);
   REGISTERS_reg_22_22_inst : DFF_X1 port map( D => n1869, CK => n462, Q => 
                           REGISTERS_22_22_port, QN => n_1745);
   REGISTERS_reg_22_21_inst : DFF_X1 port map( D => n1868, CK => n462, Q => 
                           REGISTERS_22_21_port, QN => n_1746);
   REGISTERS_reg_22_20_inst : DFF_X1 port map( D => n1867, CK => n462, Q => 
                           REGISTERS_22_20_port, QN => n_1747);
   REGISTERS_reg_22_19_inst : DFF_X1 port map( D => n1866, CK => n462, Q => 
                           REGISTERS_22_19_port, QN => n_1748);
   REGISTERS_reg_22_18_inst : DFF_X1 port map( D => n1865, CK => n462, Q => 
                           REGISTERS_22_18_port, QN => n_1749);
   REGISTERS_reg_22_17_inst : DFF_X1 port map( D => n1864, CK => n462, Q => 
                           REGISTERS_22_17_port, QN => n_1750);
   REGISTERS_reg_22_16_inst : DFF_X1 port map( D => n1863, CK => n462, Q => 
                           REGISTERS_22_16_port, QN => n_1751);
   REGISTERS_reg_22_15_inst : DFF_X1 port map( D => n1862, CK => n463, Q => 
                           REGISTERS_22_15_port, QN => n_1752);
   REGISTERS_reg_22_14_inst : DFF_X1 port map( D => n1861, CK => n463, Q => 
                           REGISTERS_22_14_port, QN => n_1753);
   REGISTERS_reg_22_13_inst : DFF_X1 port map( D => n1860, CK => n463, Q => 
                           REGISTERS_22_13_port, QN => n_1754);
   REGISTERS_reg_22_12_inst : DFF_X1 port map( D => n1859, CK => n463, Q => 
                           REGISTERS_22_12_port, QN => n_1755);
   REGISTERS_reg_22_11_inst : DFF_X1 port map( D => n1858, CK => n463, Q => 
                           REGISTERS_22_11_port, QN => n_1756);
   REGISTERS_reg_22_10_inst : DFF_X1 port map( D => n1857, CK => n463, Q => 
                           REGISTERS_22_10_port, QN => n_1757);
   REGISTERS_reg_22_9_inst : DFF_X1 port map( D => n1856, CK => n463, Q => 
                           REGISTERS_22_9_port, QN => n_1758);
   REGISTERS_reg_22_8_inst : DFF_X1 port map( D => n1855, CK => n463, Q => 
                           REGISTERS_22_8_port, QN => n_1759);
   REGISTERS_reg_22_7_inst : DFF_X1 port map( D => n1854, CK => n463, Q => 
                           REGISTERS_22_7_port, QN => n_1760);
   REGISTERS_reg_22_6_inst : DFF_X1 port map( D => n1853, CK => n463, Q => 
                           REGISTERS_22_6_port, QN => n_1761);
   REGISTERS_reg_22_5_inst : DFF_X1 port map( D => n1852, CK => n463, Q => 
                           REGISTERS_22_5_port, QN => n_1762);
   REGISTERS_reg_22_4_inst : DFF_X1 port map( D => n1851, CK => n464, Q => 
                           REGISTERS_22_4_port, QN => n_1763);
   REGISTERS_reg_22_3_inst : DFF_X1 port map( D => n1850, CK => n464, Q => 
                           REGISTERS_22_3_port, QN => n_1764);
   REGISTERS_reg_22_2_inst : DFF_X1 port map( D => n1849, CK => n464, Q => 
                           REGISTERS_22_2_port, QN => n_1765);
   REGISTERS_reg_22_1_inst : DFF_X1 port map( D => n1848, CK => n464, Q => 
                           REGISTERS_22_1_port, QN => n_1766);
   REGISTERS_reg_22_0_inst : DFF_X1 port map( D => n1847, CK => n464, Q => 
                           REGISTERS_22_0_port, QN => n_1767);
   REGISTERS_reg_23_31_inst : DFF_X1 port map( D => n1846, CK => n464, Q => 
                           REGISTERS_23_31_port, QN => n_1768);
   REGISTERS_reg_23_30_inst : DFF_X1 port map( D => n1845, CK => n464, Q => 
                           REGISTERS_23_30_port, QN => n_1769);
   REGISTERS_reg_23_29_inst : DFF_X1 port map( D => n1844, CK => n464, Q => 
                           REGISTERS_23_29_port, QN => n_1770);
   REGISTERS_reg_23_28_inst : DFF_X1 port map( D => n1843, CK => n464, Q => 
                           REGISTERS_23_28_port, QN => n_1771);
   REGISTERS_reg_23_27_inst : DFF_X1 port map( D => n1842, CK => n464, Q => 
                           REGISTERS_23_27_port, QN => n_1772);
   REGISTERS_reg_23_26_inst : DFF_X1 port map( D => n1841, CK => n464, Q => 
                           REGISTERS_23_26_port, QN => n_1773);
   REGISTERS_reg_23_25_inst : DFF_X1 port map( D => n1840, CK => n465, Q => 
                           REGISTERS_23_25_port, QN => n_1774);
   REGISTERS_reg_23_24_inst : DFF_X1 port map( D => n1839, CK => n465, Q => 
                           REGISTERS_23_24_port, QN => n_1775);
   REGISTERS_reg_23_23_inst : DFF_X1 port map( D => n1838, CK => n465, Q => 
                           REGISTERS_23_23_port, QN => n_1776);
   REGISTERS_reg_23_22_inst : DFF_X1 port map( D => n1837, CK => n465, Q => 
                           REGISTERS_23_22_port, QN => n_1777);
   REGISTERS_reg_23_21_inst : DFF_X1 port map( D => n1836, CK => n465, Q => 
                           REGISTERS_23_21_port, QN => n_1778);
   REGISTERS_reg_23_20_inst : DFF_X1 port map( D => n1835, CK => n465, Q => 
                           REGISTERS_23_20_port, QN => n_1779);
   REGISTERS_reg_23_19_inst : DFF_X1 port map( D => n1834, CK => n465, Q => 
                           REGISTERS_23_19_port, QN => n_1780);
   REGISTERS_reg_23_18_inst : DFF_X1 port map( D => n1833, CK => n465, Q => 
                           REGISTERS_23_18_port, QN => n_1781);
   REGISTERS_reg_23_17_inst : DFF_X1 port map( D => n1832, CK => n465, Q => 
                           REGISTERS_23_17_port, QN => n_1782);
   REGISTERS_reg_23_16_inst : DFF_X1 port map( D => n1831, CK => n465, Q => 
                           REGISTERS_23_16_port, QN => n_1783);
   REGISTERS_reg_23_15_inst : DFF_X1 port map( D => n1830, CK => n465, Q => 
                           REGISTERS_23_15_port, QN => n_1784);
   REGISTERS_reg_23_14_inst : DFF_X1 port map( D => n1829, CK => n466, Q => 
                           REGISTERS_23_14_port, QN => n_1785);
   REGISTERS_reg_23_13_inst : DFF_X1 port map( D => n1828, CK => n466, Q => 
                           REGISTERS_23_13_port, QN => n_1786);
   REGISTERS_reg_23_12_inst : DFF_X1 port map( D => n1827, CK => n466, Q => 
                           REGISTERS_23_12_port, QN => n_1787);
   REGISTERS_reg_23_11_inst : DFF_X1 port map( D => n1826, CK => n466, Q => 
                           REGISTERS_23_11_port, QN => n_1788);
   REGISTERS_reg_23_10_inst : DFF_X1 port map( D => n1825, CK => n466, Q => 
                           REGISTERS_23_10_port, QN => n_1789);
   REGISTERS_reg_23_9_inst : DFF_X1 port map( D => n1824, CK => n466, Q => 
                           REGISTERS_23_9_port, QN => n_1790);
   REGISTERS_reg_23_8_inst : DFF_X1 port map( D => n1823, CK => n466, Q => 
                           REGISTERS_23_8_port, QN => n_1791);
   REGISTERS_reg_23_7_inst : DFF_X1 port map( D => n1822, CK => n466, Q => 
                           REGISTERS_23_7_port, QN => n_1792);
   REGISTERS_reg_23_6_inst : DFF_X1 port map( D => n1821, CK => n466, Q => 
                           REGISTERS_23_6_port, QN => n_1793);
   REGISTERS_reg_23_5_inst : DFF_X1 port map( D => n1820, CK => n466, Q => 
                           REGISTERS_23_5_port, QN => n_1794);
   REGISTERS_reg_23_4_inst : DFF_X1 port map( D => n1819, CK => n466, Q => 
                           REGISTERS_23_4_port, QN => n_1795);
   REGISTERS_reg_23_3_inst : DFF_X1 port map( D => n1818, CK => n467, Q => 
                           REGISTERS_23_3_port, QN => n_1796);
   REGISTERS_reg_23_2_inst : DFF_X1 port map( D => n1817, CK => n467, Q => 
                           REGISTERS_23_2_port, QN => n_1797);
   REGISTERS_reg_23_1_inst : DFF_X1 port map( D => n1816, CK => n467, Q => 
                           REGISTERS_23_1_port, QN => n_1798);
   REGISTERS_reg_23_0_inst : DFF_X1 port map( D => n1815, CK => n467, Q => 
                           REGISTERS_23_0_port, QN => n_1799);
   REGISTERS_reg_24_31_inst : DFF_X1 port map( D => n1814, CK => n418, Q => 
                           REGISTERS_24_31_port, QN => n_1800);
   REGISTERS_reg_24_30_inst : DFF_X1 port map( D => n1813, CK => n418, Q => 
                           REGISTERS_24_30_port, QN => n_1801);
   REGISTERS_reg_24_29_inst : DFF_X1 port map( D => n1812, CK => n418, Q => 
                           REGISTERS_24_29_port, QN => n_1802);
   REGISTERS_reg_24_28_inst : DFF_X1 port map( D => n1811, CK => n418, Q => 
                           REGISTERS_24_28_port, QN => n_1803);
   REGISTERS_reg_24_27_inst : DFF_X1 port map( D => n1810, CK => n418, Q => 
                           REGISTERS_24_27_port, QN => n_1804);
   REGISTERS_reg_24_26_inst : DFF_X1 port map( D => n1809, CK => n418, Q => 
                           REGISTERS_24_26_port, QN => n_1805);
   REGISTERS_reg_24_25_inst : DFF_X1 port map( D => n1808, CK => n419, Q => 
                           REGISTERS_24_25_port, QN => n_1806);
   REGISTERS_reg_24_24_inst : DFF_X1 port map( D => n1807, CK => n419, Q => 
                           REGISTERS_24_24_port, QN => n_1807);
   REGISTERS_reg_24_23_inst : DFF_X1 port map( D => n1806, CK => n419, Q => 
                           REGISTERS_24_23_port, QN => n_1808);
   REGISTERS_reg_24_22_inst : DFF_X1 port map( D => n1805, CK => n419, Q => 
                           REGISTERS_24_22_port, QN => n_1809);
   REGISTERS_reg_24_21_inst : DFF_X1 port map( D => n1804, CK => n419, Q => 
                           REGISTERS_24_21_port, QN => n_1810);
   REGISTERS_reg_24_20_inst : DFF_X1 port map( D => n1803, CK => n420, Q => 
                           REGISTERS_24_20_port, QN => n_1811);
   REGISTERS_reg_24_19_inst : DFF_X1 port map( D => n1802, CK => n420, Q => 
                           REGISTERS_24_19_port, QN => n_1812);
   REGISTERS_reg_24_18_inst : DFF_X1 port map( D => n1801, CK => n420, Q => 
                           REGISTERS_24_18_port, QN => n_1813);
   REGISTERS_reg_24_17_inst : DFF_X1 port map( D => n1800, CK => n420, Q => 
                           REGISTERS_24_17_port, QN => n_1814);
   REGISTERS_reg_24_16_inst : DFF_X1 port map( D => n1799, CK => n420, Q => 
                           REGISTERS_24_16_port, QN => n_1815);
   REGISTERS_reg_24_15_inst : DFF_X1 port map( D => n1798, CK => n420, Q => 
                           REGISTERS_24_15_port, QN => n_1816);
   REGISTERS_reg_24_14_inst : DFF_X1 port map( D => n1797, CK => n421, Q => 
                           REGISTERS_24_14_port, QN => n_1817);
   REGISTERS_reg_24_13_inst : DFF_X1 port map( D => n1796, CK => n421, Q => 
                           REGISTERS_24_13_port, QN => n_1818);
   REGISTERS_reg_24_12_inst : DFF_X1 port map( D => n1795, CK => n421, Q => 
                           REGISTERS_24_12_port, QN => n_1819);
   REGISTERS_reg_24_11_inst : DFF_X1 port map( D => n1794, CK => n421, Q => 
                           REGISTERS_24_11_port, QN => n_1820);
   REGISTERS_reg_24_10_inst : DFF_X1 port map( D => n1793, CK => n421, Q => 
                           REGISTERS_24_10_port, QN => n_1821);
   REGISTERS_reg_24_9_inst : DFF_X1 port map( D => n1792, CK => n422, Q => 
                           REGISTERS_24_9_port, QN => n_1822);
   REGISTERS_reg_24_8_inst : DFF_X1 port map( D => n1791, CK => n422, Q => 
                           REGISTERS_24_8_port, QN => n_1823);
   REGISTERS_reg_24_7_inst : DFF_X1 port map( D => n1790, CK => n422, Q => 
                           REGISTERS_24_7_port, QN => n_1824);
   REGISTERS_reg_24_6_inst : DFF_X1 port map( D => n1789, CK => n422, Q => 
                           REGISTERS_24_6_port, QN => n_1825);
   REGISTERS_reg_24_5_inst : DFF_X1 port map( D => n1788, CK => n422, Q => 
                           REGISTERS_24_5_port, QN => n_1826);
   REGISTERS_reg_24_4_inst : DFF_X1 port map( D => n1787, CK => n422, Q => 
                           REGISTERS_24_4_port, QN => n_1827);
   REGISTERS_reg_24_3_inst : DFF_X1 port map( D => n1786, CK => n423, Q => 
                           REGISTERS_24_3_port, QN => n_1828);
   REGISTERS_reg_24_2_inst : DFF_X1 port map( D => n1785, CK => n423, Q => 
                           REGISTERS_24_2_port, QN => n_1829);
   REGISTERS_reg_24_1_inst : DFF_X1 port map( D => n1784, CK => n423, Q => 
                           REGISTERS_24_1_port, QN => n_1830);
   REGISTERS_reg_24_0_inst : DFF_X1 port map( D => n1783, CK => n423, Q => 
                           REGISTERS_24_0_port, QN => n_1831);
   REGISTERS_reg_25_31_inst : DFF_X1 port map( D => n1782, CK => n423, Q => 
                           REGISTERS_25_31_port, QN => n_1832);
   REGISTERS_reg_25_30_inst : DFF_X1 port map( D => n1781, CK => n423, Q => 
                           REGISTERS_25_30_port, QN => n_1833);
   REGISTERS_reg_25_29_inst : DFF_X1 port map( D => n1780, CK => n423, Q => 
                           REGISTERS_25_29_port, QN => n_1834);
   REGISTERS_reg_25_28_inst : DFF_X1 port map( D => n1779, CK => n424, Q => 
                           REGISTERS_25_28_port, QN => n_1835);
   REGISTERS_reg_25_27_inst : DFF_X1 port map( D => n1778, CK => n424, Q => 
                           REGISTERS_25_27_port, QN => n_1836);
   REGISTERS_reg_25_26_inst : DFF_X1 port map( D => n1777, CK => n424, Q => 
                           REGISTERS_25_26_port, QN => n_1837);
   REGISTERS_reg_25_25_inst : DFF_X1 port map( D => n1776, CK => n424, Q => 
                           REGISTERS_25_25_port, QN => n_1838);
   REGISTERS_reg_25_24_inst : DFF_X1 port map( D => n1775, CK => n424, Q => 
                           REGISTERS_25_24_port, QN => n_1839);
   REGISTERS_reg_25_23_inst : DFF_X1 port map( D => n1774, CK => n424, Q => 
                           REGISTERS_25_23_port, QN => n_1840);
   REGISTERS_reg_25_22_inst : DFF_X1 port map( D => n1773, CK => n424, Q => 
                           REGISTERS_25_22_port, QN => n_1841);
   REGISTERS_reg_25_21_inst : DFF_X1 port map( D => n1772, CK => n424, Q => 
                           REGISTERS_25_21_port, QN => n_1842);
   REGISTERS_reg_25_20_inst : DFF_X1 port map( D => n1771, CK => n424, Q => 
                           REGISTERS_25_20_port, QN => n_1843);
   REGISTERS_reg_25_19_inst : DFF_X1 port map( D => n1770, CK => n424, Q => 
                           REGISTERS_25_19_port, QN => n_1844);
   REGISTERS_reg_25_18_inst : DFF_X1 port map( D => n1769, CK => n424, Q => 
                           REGISTERS_25_18_port, QN => n_1845);
   REGISTERS_reg_25_17_inst : DFF_X1 port map( D => n1768, CK => n425, Q => 
                           REGISTERS_25_17_port, QN => n_1846);
   REGISTERS_reg_25_16_inst : DFF_X1 port map( D => n1767, CK => n425, Q => 
                           REGISTERS_25_16_port, QN => n_1847);
   REGISTERS_reg_25_15_inst : DFF_X1 port map( D => n1766, CK => n425, Q => 
                           REGISTERS_25_15_port, QN => n_1848);
   REGISTERS_reg_25_14_inst : DFF_X1 port map( D => n1765, CK => n425, Q => 
                           REGISTERS_25_14_port, QN => n_1849);
   REGISTERS_reg_25_13_inst : DFF_X1 port map( D => n1764, CK => n425, Q => 
                           REGISTERS_25_13_port, QN => n_1850);
   REGISTERS_reg_25_12_inst : DFF_X1 port map( D => n1763, CK => n425, Q => 
                           REGISTERS_25_12_port, QN => n_1851);
   REGISTERS_reg_25_11_inst : DFF_X1 port map( D => n1762, CK => n425, Q => 
                           REGISTERS_25_11_port, QN => n_1852);
   REGISTERS_reg_25_10_inst : DFF_X1 port map( D => n1761, CK => n425, Q => 
                           REGISTERS_25_10_port, QN => n_1853);
   REGISTERS_reg_25_9_inst : DFF_X1 port map( D => n1760, CK => n425, Q => 
                           REGISTERS_25_9_port, QN => n_1854);
   REGISTERS_reg_25_8_inst : DFF_X1 port map( D => n1759, CK => n425, Q => 
                           REGISTERS_25_8_port, QN => n_1855);
   REGISTERS_reg_25_7_inst : DFF_X1 port map( D => n1758, CK => n425, Q => 
                           REGISTERS_25_7_port, QN => n_1856);
   REGISTERS_reg_25_6_inst : DFF_X1 port map( D => n1757, CK => n426, Q => 
                           REGISTERS_25_6_port, QN => n_1857);
   REGISTERS_reg_25_5_inst : DFF_X1 port map( D => n1756, CK => n426, Q => 
                           REGISTERS_25_5_port, QN => n_1858);
   REGISTERS_reg_25_4_inst : DFF_X1 port map( D => n1755, CK => n426, Q => 
                           REGISTERS_25_4_port, QN => n_1859);
   REGISTERS_reg_25_3_inst : DFF_X1 port map( D => n1754, CK => n426, Q => 
                           REGISTERS_25_3_port, QN => n_1860);
   REGISTERS_reg_25_2_inst : DFF_X1 port map( D => n1753, CK => n426, Q => 
                           REGISTERS_25_2_port, QN => n_1861);
   REGISTERS_reg_25_1_inst : DFF_X1 port map( D => n1752, CK => n426, Q => 
                           REGISTERS_25_1_port, QN => n_1862);
   REGISTERS_reg_25_0_inst : DFF_X1 port map( D => n1751, CK => n426, Q => 
                           REGISTERS_25_0_port, QN => n_1863);
   REGISTERS_reg_26_31_inst : DFF_X1 port map( D => n1750, CK => n426, Q => 
                           REGISTERS_26_31_port, QN => n_1864);
   REGISTERS_reg_26_30_inst : DFF_X1 port map( D => n1749, CK => n426, Q => 
                           REGISTERS_26_30_port, QN => n_1865);
   REGISTERS_reg_26_29_inst : DFF_X1 port map( D => n1748, CK => n426, Q => 
                           REGISTERS_26_29_port, QN => n_1866);
   REGISTERS_reg_26_28_inst : DFF_X1 port map( D => n1747, CK => n426, Q => 
                           REGISTERS_26_28_port, QN => n_1867);
   REGISTERS_reg_26_27_inst : DFF_X1 port map( D => n1746, CK => n427, Q => 
                           REGISTERS_26_27_port, QN => n_1868);
   REGISTERS_reg_26_26_inst : DFF_X1 port map( D => n1745, CK => n427, Q => 
                           REGISTERS_26_26_port, QN => n_1869);
   REGISTERS_reg_26_25_inst : DFF_X1 port map( D => n1744, CK => n427, Q => 
                           REGISTERS_26_25_port, QN => n_1870);
   REGISTERS_reg_26_24_inst : DFF_X1 port map( D => n1743, CK => n427, Q => 
                           REGISTERS_26_24_port, QN => n_1871);
   REGISTERS_reg_26_23_inst : DFF_X1 port map( D => n1742, CK => n427, Q => 
                           REGISTERS_26_23_port, QN => n_1872);
   REGISTERS_reg_26_22_inst : DFF_X1 port map( D => n1741, CK => n427, Q => 
                           REGISTERS_26_22_port, QN => n_1873);
   REGISTERS_reg_26_21_inst : DFF_X1 port map( D => n1740, CK => n427, Q => 
                           REGISTERS_26_21_port, QN => n_1874);
   REGISTERS_reg_26_20_inst : DFF_X1 port map( D => n1739, CK => n427, Q => 
                           REGISTERS_26_20_port, QN => n_1875);
   REGISTERS_reg_26_19_inst : DFF_X1 port map( D => n1738, CK => n427, Q => 
                           REGISTERS_26_19_port, QN => n_1876);
   REGISTERS_reg_26_18_inst : DFF_X1 port map( D => n1737, CK => n427, Q => 
                           REGISTERS_26_18_port, QN => n_1877);
   REGISTERS_reg_26_17_inst : DFF_X1 port map( D => n1736, CK => n427, Q => 
                           REGISTERS_26_17_port, QN => n_1878);
   REGISTERS_reg_26_16_inst : DFF_X1 port map( D => n1735, CK => n428, Q => 
                           REGISTERS_26_16_port, QN => n_1879);
   REGISTERS_reg_26_15_inst : DFF_X1 port map( D => n1734, CK => n428, Q => 
                           REGISTERS_26_15_port, QN => n_1880);
   REGISTERS_reg_26_14_inst : DFF_X1 port map( D => n1733, CK => n428, Q => 
                           REGISTERS_26_14_port, QN => n_1881);
   REGISTERS_reg_26_13_inst : DFF_X1 port map( D => n1732, CK => n428, Q => 
                           REGISTERS_26_13_port, QN => n_1882);
   REGISTERS_reg_26_12_inst : DFF_X1 port map( D => n1731, CK => n428, Q => 
                           REGISTERS_26_12_port, QN => n_1883);
   REGISTERS_reg_26_11_inst : DFF_X1 port map( D => n1730, CK => n428, Q => 
                           REGISTERS_26_11_port, QN => n_1884);
   REGISTERS_reg_26_10_inst : DFF_X1 port map( D => n1729, CK => n428, Q => 
                           REGISTERS_26_10_port, QN => n_1885);
   REGISTERS_reg_26_9_inst : DFF_X1 port map( D => n1728, CK => n428, Q => 
                           REGISTERS_26_9_port, QN => n_1886);
   REGISTERS_reg_26_8_inst : DFF_X1 port map( D => n1727, CK => n428, Q => 
                           REGISTERS_26_8_port, QN => n_1887);
   REGISTERS_reg_26_7_inst : DFF_X1 port map( D => n1726, CK => n428, Q => 
                           REGISTERS_26_7_port, QN => n_1888);
   REGISTERS_reg_26_6_inst : DFF_X1 port map( D => n1725, CK => n428, Q => 
                           REGISTERS_26_6_port, QN => n_1889);
   REGISTERS_reg_26_5_inst : DFF_X1 port map( D => n1724, CK => n429, Q => 
                           REGISTERS_26_5_port, QN => n_1890);
   REGISTERS_reg_26_4_inst : DFF_X1 port map( D => n1723, CK => n429, Q => 
                           REGISTERS_26_4_port, QN => n_1891);
   REGISTERS_reg_26_3_inst : DFF_X1 port map( D => n1722, CK => n429, Q => 
                           REGISTERS_26_3_port, QN => n_1892);
   REGISTERS_reg_26_2_inst : DFF_X1 port map( D => n1721, CK => n429, Q => 
                           REGISTERS_26_2_port, QN => n_1893);
   REGISTERS_reg_26_1_inst : DFF_X1 port map( D => n1720, CK => n429, Q => 
                           REGISTERS_26_1_port, QN => n_1894);
   REGISTERS_reg_26_0_inst : DFF_X1 port map( D => n1719, CK => n429, Q => 
                           REGISTERS_26_0_port, QN => n_1895);
   REGISTERS_reg_27_31_inst : DFF_X1 port map( D => n1718, CK => n429, Q => 
                           REGISTERS_27_31_port, QN => n_1896);
   REGISTERS_reg_27_30_inst : DFF_X1 port map( D => n1717, CK => n429, Q => 
                           REGISTERS_27_30_port, QN => n_1897);
   REGISTERS_reg_27_29_inst : DFF_X1 port map( D => n1716, CK => n429, Q => 
                           REGISTERS_27_29_port, QN => n_1898);
   REGISTERS_reg_27_28_inst : DFF_X1 port map( D => n1715, CK => n429, Q => 
                           REGISTERS_27_28_port, QN => n_1899);
   REGISTERS_reg_27_27_inst : DFF_X1 port map( D => n1714, CK => n429, Q => 
                           REGISTERS_27_27_port, QN => n_1900);
   REGISTERS_reg_27_26_inst : DFF_X1 port map( D => n1713, CK => n430, Q => 
                           REGISTERS_27_26_port, QN => n_1901);
   REGISTERS_reg_27_25_inst : DFF_X1 port map( D => n1712, CK => n430, Q => 
                           REGISTERS_27_25_port, QN => n_1902);
   REGISTERS_reg_27_24_inst : DFF_X1 port map( D => n1711, CK => n430, Q => 
                           REGISTERS_27_24_port, QN => n_1903);
   REGISTERS_reg_27_23_inst : DFF_X1 port map( D => n1710, CK => n430, Q => 
                           REGISTERS_27_23_port, QN => n_1904);
   REGISTERS_reg_27_22_inst : DFF_X1 port map( D => n1709, CK => n430, Q => 
                           REGISTERS_27_22_port, QN => n_1905);
   REGISTERS_reg_27_21_inst : DFF_X1 port map( D => n1708, CK => n430, Q => 
                           REGISTERS_27_21_port, QN => n_1906);
   REGISTERS_reg_27_20_inst : DFF_X1 port map( D => n1707, CK => n430, Q => 
                           REGISTERS_27_20_port, QN => n_1907);
   REGISTERS_reg_27_19_inst : DFF_X1 port map( D => n1706, CK => n430, Q => 
                           REGISTERS_27_19_port, QN => n_1908);
   REGISTERS_reg_27_18_inst : DFF_X1 port map( D => n1705, CK => n430, Q => 
                           REGISTERS_27_18_port, QN => n_1909);
   REGISTERS_reg_27_17_inst : DFF_X1 port map( D => n1704, CK => n430, Q => 
                           REGISTERS_27_17_port, QN => n_1910);
   REGISTERS_reg_27_16_inst : DFF_X1 port map( D => n1703, CK => n430, Q => 
                           REGISTERS_27_16_port, QN => n_1911);
   REGISTERS_reg_27_15_inst : DFF_X1 port map( D => n1702, CK => n431, Q => 
                           REGISTERS_27_15_port, QN => n_1912);
   REGISTERS_reg_27_14_inst : DFF_X1 port map( D => n1701, CK => n431, Q => 
                           REGISTERS_27_14_port, QN => n_1913);
   REGISTERS_reg_27_13_inst : DFF_X1 port map( D => n1700, CK => n431, Q => 
                           REGISTERS_27_13_port, QN => n_1914);
   REGISTERS_reg_27_12_inst : DFF_X1 port map( D => n1699, CK => n431, Q => 
                           REGISTERS_27_12_port, QN => n_1915);
   REGISTERS_reg_27_11_inst : DFF_X1 port map( D => n1698, CK => n431, Q => 
                           REGISTERS_27_11_port, QN => n_1916);
   REGISTERS_reg_27_10_inst : DFF_X1 port map( D => n1697, CK => n431, Q => 
                           REGISTERS_27_10_port, QN => n_1917);
   REGISTERS_reg_27_9_inst : DFF_X1 port map( D => n1696, CK => n431, Q => 
                           REGISTERS_27_9_port, QN => n_1918);
   REGISTERS_reg_27_8_inst : DFF_X1 port map( D => n1695, CK => n431, Q => 
                           REGISTERS_27_8_port, QN => n_1919);
   REGISTERS_reg_27_7_inst : DFF_X1 port map( D => n1694, CK => n431, Q => 
                           REGISTERS_27_7_port, QN => n_1920);
   REGISTERS_reg_27_6_inst : DFF_X1 port map( D => n1693, CK => n431, Q => 
                           REGISTERS_27_6_port, QN => n_1921);
   REGISTERS_reg_27_5_inst : DFF_X1 port map( D => n1692, CK => n431, Q => 
                           REGISTERS_27_5_port, QN => n_1922);
   REGISTERS_reg_27_4_inst : DFF_X1 port map( D => n1691, CK => n432, Q => 
                           REGISTERS_27_4_port, QN => n_1923);
   REGISTERS_reg_27_3_inst : DFF_X1 port map( D => n1690, CK => n432, Q => 
                           REGISTERS_27_3_port, QN => n_1924);
   REGISTERS_reg_27_2_inst : DFF_X1 port map( D => n1689, CK => n432, Q => 
                           REGISTERS_27_2_port, QN => n_1925);
   REGISTERS_reg_27_1_inst : DFF_X1 port map( D => n1688, CK => n432, Q => 
                           REGISTERS_27_1_port, QN => n_1926);
   REGISTERS_reg_27_0_inst : DFF_X1 port map( D => n1687, CK => n432, Q => 
                           REGISTERS_27_0_port, QN => n_1927);
   REGISTERS_reg_28_31_inst : DFF_X1 port map( D => n1686, CK => n432, Q => 
                           REGISTERS_28_31_port, QN => n_1928);
   REGISTERS_reg_28_30_inst : DFF_X1 port map( D => n1685, CK => n432, Q => 
                           REGISTERS_28_30_port, QN => n_1929);
   REGISTERS_reg_28_29_inst : DFF_X1 port map( D => n1684, CK => n432, Q => 
                           REGISTERS_28_29_port, QN => n_1930);
   REGISTERS_reg_28_28_inst : DFF_X1 port map( D => n1683, CK => n432, Q => 
                           REGISTERS_28_28_port, QN => n_1931);
   REGISTERS_reg_28_27_inst : DFF_X1 port map( D => n1682, CK => n432, Q => 
                           REGISTERS_28_27_port, QN => n_1932);
   REGISTERS_reg_28_26_inst : DFF_X1 port map( D => n1681, CK => n432, Q => 
                           REGISTERS_28_26_port, QN => n_1933);
   REGISTERS_reg_28_25_inst : DFF_X1 port map( D => n1680, CK => n433, Q => 
                           REGISTERS_28_25_port, QN => n_1934);
   REGISTERS_reg_28_24_inst : DFF_X1 port map( D => n1679, CK => n433, Q => 
                           REGISTERS_28_24_port, QN => n_1935);
   REGISTERS_reg_28_23_inst : DFF_X1 port map( D => n1678, CK => n433, Q => 
                           REGISTERS_28_23_port, QN => n_1936);
   REGISTERS_reg_28_22_inst : DFF_X1 port map( D => n1677, CK => n433, Q => 
                           REGISTERS_28_22_port, QN => n_1937);
   REGISTERS_reg_28_21_inst : DFF_X1 port map( D => n1676, CK => n433, Q => 
                           REGISTERS_28_21_port, QN => n_1938);
   REGISTERS_reg_28_20_inst : DFF_X1 port map( D => n1675, CK => n433, Q => 
                           REGISTERS_28_20_port, QN => n_1939);
   REGISTERS_reg_28_19_inst : DFF_X1 port map( D => n1674, CK => n433, Q => 
                           REGISTERS_28_19_port, QN => n_1940);
   REGISTERS_reg_28_18_inst : DFF_X1 port map( D => n1673, CK => n433, Q => 
                           REGISTERS_28_18_port, QN => n_1941);
   REGISTERS_reg_28_17_inst : DFF_X1 port map( D => n1672, CK => n433, Q => 
                           REGISTERS_28_17_port, QN => n_1942);
   REGISTERS_reg_28_16_inst : DFF_X1 port map( D => n1671, CK => n433, Q => 
                           REGISTERS_28_16_port, QN => n_1943);
   REGISTERS_reg_28_15_inst : DFF_X1 port map( D => n1670, CK => n433, Q => 
                           REGISTERS_28_15_port, QN => n_1944);
   REGISTERS_reg_28_14_inst : DFF_X1 port map( D => n1669, CK => n434, Q => 
                           REGISTERS_28_14_port, QN => n_1945);
   REGISTERS_reg_28_13_inst : DFF_X1 port map( D => n1668, CK => n434, Q => 
                           REGISTERS_28_13_port, QN => n_1946);
   REGISTERS_reg_28_12_inst : DFF_X1 port map( D => n1667, CK => n434, Q => 
                           REGISTERS_28_12_port, QN => n_1947);
   REGISTERS_reg_28_11_inst : DFF_X1 port map( D => n1666, CK => n434, Q => 
                           REGISTERS_28_11_port, QN => n_1948);
   REGISTERS_reg_28_10_inst : DFF_X1 port map( D => n1665, CK => n434, Q => 
                           REGISTERS_28_10_port, QN => n_1949);
   REGISTERS_reg_28_9_inst : DFF_X1 port map( D => n1664, CK => n434, Q => 
                           REGISTERS_28_9_port, QN => n_1950);
   REGISTERS_reg_28_8_inst : DFF_X1 port map( D => n1663, CK => n434, Q => 
                           REGISTERS_28_8_port, QN => n_1951);
   REGISTERS_reg_28_7_inst : DFF_X1 port map( D => n1662, CK => n434, Q => 
                           REGISTERS_28_7_port, QN => n_1952);
   REGISTERS_reg_28_6_inst : DFF_X1 port map( D => n1661, CK => n434, Q => 
                           REGISTERS_28_6_port, QN => n_1953);
   REGISTERS_reg_28_5_inst : DFF_X1 port map( D => n1660, CK => n434, Q => 
                           REGISTERS_28_5_port, QN => n_1954);
   REGISTERS_reg_28_4_inst : DFF_X1 port map( D => n1659, CK => n434, Q => 
                           REGISTERS_28_4_port, QN => n_1955);
   REGISTERS_reg_28_3_inst : DFF_X1 port map( D => n1658, CK => n435, Q => 
                           REGISTERS_28_3_port, QN => n_1956);
   REGISTERS_reg_28_2_inst : DFF_X1 port map( D => n1657, CK => n435, Q => 
                           REGISTERS_28_2_port, QN => n_1957);
   REGISTERS_reg_28_1_inst : DFF_X1 port map( D => n1656, CK => n435, Q => 
                           REGISTERS_28_1_port, QN => n_1958);
   REGISTERS_reg_28_0_inst : DFF_X1 port map( D => n1655, CK => n435, Q => 
                           REGISTERS_28_0_port, QN => n_1959);
   REGISTERS_reg_29_31_inst : DFF_X1 port map( D => n1654, CK => n435, Q => 
                           REGISTERS_29_31_port, QN => n_1960);
   REGISTERS_reg_29_30_inst : DFF_X1 port map( D => n1653, CK => n435, Q => 
                           REGISTERS_29_30_port, QN => n_1961);
   REGISTERS_reg_29_29_inst : DFF_X1 port map( D => n1652, CK => n435, Q => 
                           REGISTERS_29_29_port, QN => n_1962);
   REGISTERS_reg_29_28_inst : DFF_X1 port map( D => n1651, CK => n435, Q => 
                           REGISTERS_29_28_port, QN => n_1963);
   REGISTERS_reg_29_27_inst : DFF_X1 port map( D => n1650, CK => n435, Q => 
                           REGISTERS_29_27_port, QN => n_1964);
   REGISTERS_reg_29_26_inst : DFF_X1 port map( D => n1649, CK => n435, Q => 
                           REGISTERS_29_26_port, QN => n_1965);
   REGISTERS_reg_29_25_inst : DFF_X1 port map( D => n1648, CK => n435, Q => 
                           REGISTERS_29_25_port, QN => n_1966);
   REGISTERS_reg_29_24_inst : DFF_X1 port map( D => n1647, CK => n436, Q => 
                           REGISTERS_29_24_port, QN => n_1967);
   REGISTERS_reg_29_23_inst : DFF_X1 port map( D => n1646, CK => n436, Q => 
                           REGISTERS_29_23_port, QN => n_1968);
   REGISTERS_reg_29_22_inst : DFF_X1 port map( D => n1645, CK => n436, Q => 
                           REGISTERS_29_22_port, QN => n_1969);
   REGISTERS_reg_29_21_inst : DFF_X1 port map( D => n1644, CK => n436, Q => 
                           REGISTERS_29_21_port, QN => n_1970);
   REGISTERS_reg_29_20_inst : DFF_X1 port map( D => n1643, CK => n436, Q => 
                           REGISTERS_29_20_port, QN => n_1971);
   REGISTERS_reg_29_19_inst : DFF_X1 port map( D => n1642, CK => n436, Q => 
                           REGISTERS_29_19_port, QN => n_1972);
   REGISTERS_reg_29_18_inst : DFF_X1 port map( D => n1641, CK => n436, Q => 
                           REGISTERS_29_18_port, QN => n_1973);
   REGISTERS_reg_29_17_inst : DFF_X1 port map( D => n1640, CK => n436, Q => 
                           REGISTERS_29_17_port, QN => n_1974);
   REGISTERS_reg_29_16_inst : DFF_X1 port map( D => n1639, CK => n436, Q => 
                           REGISTERS_29_16_port, QN => n_1975);
   REGISTERS_reg_29_15_inst : DFF_X1 port map( D => n1638, CK => n436, Q => 
                           REGISTERS_29_15_port, QN => n_1976);
   REGISTERS_reg_29_14_inst : DFF_X1 port map( D => n1637, CK => n436, Q => 
                           REGISTERS_29_14_port, QN => n_1977);
   REGISTERS_reg_29_13_inst : DFF_X1 port map( D => n1636, CK => n437, Q => 
                           REGISTERS_29_13_port, QN => n_1978);
   REGISTERS_reg_29_12_inst : DFF_X1 port map( D => n1635, CK => n437, Q => 
                           REGISTERS_29_12_port, QN => n_1979);
   REGISTERS_reg_29_11_inst : DFF_X1 port map( D => n1634, CK => n437, Q => 
                           REGISTERS_29_11_port, QN => n_1980);
   REGISTERS_reg_29_10_inst : DFF_X1 port map( D => n1633, CK => n437, Q => 
                           REGISTERS_29_10_port, QN => n_1981);
   REGISTERS_reg_29_9_inst : DFF_X1 port map( D => n1632, CK => n437, Q => 
                           REGISTERS_29_9_port, QN => n_1982);
   REGISTERS_reg_29_8_inst : DFF_X1 port map( D => n1631, CK => n437, Q => 
                           REGISTERS_29_8_port, QN => n_1983);
   REGISTERS_reg_29_7_inst : DFF_X1 port map( D => n1630, CK => n437, Q => 
                           REGISTERS_29_7_port, QN => n_1984);
   REGISTERS_reg_29_6_inst : DFF_X1 port map( D => n1629, CK => n437, Q => 
                           REGISTERS_29_6_port, QN => n_1985);
   REGISTERS_reg_29_5_inst : DFF_X1 port map( D => n1628, CK => n437, Q => 
                           REGISTERS_29_5_port, QN => n_1986);
   REGISTERS_reg_29_4_inst : DFF_X1 port map( D => n1627, CK => n437, Q => 
                           REGISTERS_29_4_port, QN => n_1987);
   REGISTERS_reg_29_3_inst : DFF_X1 port map( D => n1626, CK => n437, Q => 
                           REGISTERS_29_3_port, QN => n_1988);
   REGISTERS_reg_29_2_inst : DFF_X1 port map( D => n1625, CK => n438, Q => 
                           REGISTERS_29_2_port, QN => n_1989);
   REGISTERS_reg_29_1_inst : DFF_X1 port map( D => n1624, CK => n438, Q => 
                           REGISTERS_29_1_port, QN => n_1990);
   REGISTERS_reg_29_0_inst : DFF_X1 port map( D => n1623, CK => n438, Q => 
                           REGISTERS_29_0_port, QN => n_1991);
   REGISTERS_reg_30_31_inst : DFF_X1 port map( D => n1622, CK => n438, Q => 
                           REGISTERS_30_31_port, QN => n_1992);
   REGISTERS_reg_30_30_inst : DFF_X1 port map( D => n1621, CK => n438, Q => 
                           REGISTERS_30_30_port, QN => n_1993);
   REGISTERS_reg_30_29_inst : DFF_X1 port map( D => n1620, CK => n438, Q => 
                           REGISTERS_30_29_port, QN => n_1994);
   REGISTERS_reg_30_28_inst : DFF_X1 port map( D => n1619, CK => n438, Q => 
                           REGISTERS_30_28_port, QN => n_1995);
   REGISTERS_reg_30_27_inst : DFF_X1 port map( D => n1618, CK => n438, Q => 
                           REGISTERS_30_27_port, QN => n_1996);
   REGISTERS_reg_30_26_inst : DFF_X1 port map( D => n1617, CK => n438, Q => 
                           REGISTERS_30_26_port, QN => n_1997);
   REGISTERS_reg_30_25_inst : DFF_X1 port map( D => n1616, CK => n438, Q => 
                           REGISTERS_30_25_port, QN => n_1998);
   REGISTERS_reg_30_24_inst : DFF_X1 port map( D => n1615, CK => n438, Q => 
                           REGISTERS_30_24_port, QN => n_1999);
   REGISTERS_reg_30_23_inst : DFF_X1 port map( D => n1614, CK => n439, Q => 
                           REGISTERS_30_23_port, QN => n_2000);
   REGISTERS_reg_30_22_inst : DFF_X1 port map( D => n1613, CK => n439, Q => 
                           REGISTERS_30_22_port, QN => n_2001);
   REGISTERS_reg_30_21_inst : DFF_X1 port map( D => n1612, CK => n439, Q => 
                           REGISTERS_30_21_port, QN => n_2002);
   REGISTERS_reg_30_20_inst : DFF_X1 port map( D => n1611, CK => n439, Q => 
                           REGISTERS_30_20_port, QN => n_2003);
   REGISTERS_reg_30_19_inst : DFF_X1 port map( D => n1610, CK => n439, Q => 
                           REGISTERS_30_19_port, QN => n_2004);
   REGISTERS_reg_30_18_inst : DFF_X1 port map( D => n1609, CK => n439, Q => 
                           REGISTERS_30_18_port, QN => n_2005);
   REGISTERS_reg_30_17_inst : DFF_X1 port map( D => n1608, CK => n439, Q => 
                           REGISTERS_30_17_port, QN => n_2006);
   REGISTERS_reg_30_16_inst : DFF_X1 port map( D => n1607, CK => n439, Q => 
                           REGISTERS_30_16_port, QN => n_2007);
   REGISTERS_reg_30_15_inst : DFF_X1 port map( D => n1606, CK => n439, Q => 
                           REGISTERS_30_15_port, QN => n_2008);
   REGISTERS_reg_30_14_inst : DFF_X1 port map( D => n1605, CK => n439, Q => 
                           REGISTERS_30_14_port, QN => n_2009);
   REGISTERS_reg_30_13_inst : DFF_X1 port map( D => n1604, CK => n439, Q => 
                           REGISTERS_30_13_port, QN => n_2010);
   REGISTERS_reg_30_12_inst : DFF_X1 port map( D => n1603, CK => n440, Q => 
                           REGISTERS_30_12_port, QN => n_2011);
   REGISTERS_reg_30_11_inst : DFF_X1 port map( D => n1602, CK => n440, Q => 
                           REGISTERS_30_11_port, QN => n_2012);
   REGISTERS_reg_30_10_inst : DFF_X1 port map( D => n1601, CK => n440, Q => 
                           REGISTERS_30_10_port, QN => n_2013);
   REGISTERS_reg_30_9_inst : DFF_X1 port map( D => n1600, CK => n440, Q => 
                           REGISTERS_30_9_port, QN => n_2014);
   REGISTERS_reg_30_8_inst : DFF_X1 port map( D => n1599, CK => n440, Q => 
                           REGISTERS_30_8_port, QN => n_2015);
   REGISTERS_reg_30_7_inst : DFF_X1 port map( D => n1598, CK => n440, Q => 
                           REGISTERS_30_7_port, QN => n_2016);
   REGISTERS_reg_30_6_inst : DFF_X1 port map( D => n1597, CK => n440, Q => 
                           REGISTERS_30_6_port, QN => n_2017);
   REGISTERS_reg_30_5_inst : DFF_X1 port map( D => n1596, CK => n440, Q => 
                           REGISTERS_30_5_port, QN => n_2018);
   REGISTERS_reg_30_4_inst : DFF_X1 port map( D => n1595, CK => n440, Q => 
                           REGISTERS_30_4_port, QN => n_2019);
   REGISTERS_reg_30_3_inst : DFF_X1 port map( D => n1594, CK => n440, Q => 
                           REGISTERS_30_3_port, QN => n_2020);
   REGISTERS_reg_30_2_inst : DFF_X1 port map( D => n1593, CK => n440, Q => 
                           REGISTERS_30_2_port, QN => n_2021);
   REGISTERS_reg_30_1_inst : DFF_X1 port map( D => n1592, CK => n441, Q => 
                           REGISTERS_30_1_port, QN => n_2022);
   REGISTERS_reg_30_0_inst : DFF_X1 port map( D => n1591, CK => n441, Q => 
                           REGISTERS_30_0_port, QN => n_2023);
   REGISTERS_reg_31_31_inst : DFF_X1 port map( D => n1590, CK => n441, Q => 
                           REGISTERS_31_31_port, QN => n_2024);
   REGISTERS_reg_31_30_inst : DFF_X1 port map( D => n1589, CK => n441, Q => 
                           REGISTERS_31_30_port, QN => n_2025);
   REGISTERS_reg_31_29_inst : DFF_X1 port map( D => n1588, CK => n441, Q => 
                           REGISTERS_31_29_port, QN => n_2026);
   REGISTERS_reg_31_28_inst : DFF_X1 port map( D => n1587, CK => n441, Q => 
                           REGISTERS_31_28_port, QN => n_2027);
   REGISTERS_reg_31_27_inst : DFF_X1 port map( D => n1586, CK => n441, Q => 
                           REGISTERS_31_27_port, QN => n_2028);
   REGISTERS_reg_31_26_inst : DFF_X1 port map( D => n1585, CK => n441, Q => 
                           REGISTERS_31_26_port, QN => n_2029);
   REGISTERS_reg_31_25_inst : DFF_X1 port map( D => n1584, CK => n441, Q => 
                           REGISTERS_31_25_port, QN => n_2030);
   REGISTERS_reg_31_24_inst : DFF_X1 port map( D => n1583, CK => n441, Q => 
                           REGISTERS_31_24_port, QN => n_2031);
   REGISTERS_reg_31_23_inst : DFF_X1 port map( D => n1582, CK => n441, Q => 
                           REGISTERS_31_23_port, QN => n_2032);
   REGISTERS_reg_31_22_inst : DFF_X1 port map( D => n1581, CK => n442, Q => 
                           REGISTERS_31_22_port, QN => n_2033);
   REGISTERS_reg_31_21_inst : DFF_X1 port map( D => n1580, CK => n442, Q => 
                           REGISTERS_31_21_port, QN => n_2034);
   REGISTERS_reg_31_20_inst : DFF_X1 port map( D => n1579, CK => n442, Q => 
                           REGISTERS_31_20_port, QN => n_2035);
   REGISTERS_reg_31_19_inst : DFF_X1 port map( D => n1578, CK => n442, Q => 
                           REGISTERS_31_19_port, QN => n_2036);
   REGISTERS_reg_31_18_inst : DFF_X1 port map( D => n1577, CK => n442, Q => 
                           REGISTERS_31_18_port, QN => n_2037);
   REGISTERS_reg_31_17_inst : DFF_X1 port map( D => n1576, CK => n442, Q => 
                           REGISTERS_31_17_port, QN => n_2038);
   REGISTERS_reg_31_16_inst : DFF_X1 port map( D => n1575, CK => n442, Q => 
                           REGISTERS_31_16_port, QN => n_2039);
   REGISTERS_reg_31_15_inst : DFF_X1 port map( D => n1574, CK => n442, Q => 
                           REGISTERS_31_15_port, QN => n_2040);
   REGISTERS_reg_31_14_inst : DFF_X1 port map( D => n1573, CK => n442, Q => 
                           REGISTERS_31_14_port, QN => n_2041);
   REGISTERS_reg_31_13_inst : DFF_X1 port map( D => n1572, CK => n442, Q => 
                           REGISTERS_31_13_port, QN => n_2042);
   REGISTERS_reg_31_12_inst : DFF_X1 port map( D => n1571, CK => n442, Q => 
                           REGISTERS_31_12_port, QN => n_2043);
   REGISTERS_reg_31_11_inst : DFF_X1 port map( D => n1570, CK => n443, Q => 
                           REGISTERS_31_11_port, QN => n_2044);
   REGISTERS_reg_31_10_inst : DFF_X1 port map( D => n1569, CK => n443, Q => 
                           REGISTERS_31_10_port, QN => n_2045);
   REGISTERS_reg_31_9_inst : DFF_X1 port map( D => n1568, CK => n443, Q => 
                           REGISTERS_31_9_port, QN => n_2046);
   REGISTERS_reg_31_8_inst : DFF_X1 port map( D => n1567, CK => n443, Q => 
                           REGISTERS_31_8_port, QN => n_2047);
   REGISTERS_reg_31_7_inst : DFF_X1 port map( D => n1566, CK => n443, Q => 
                           REGISTERS_31_7_port, QN => n_2048);
   REGISTERS_reg_31_6_inst : DFF_X1 port map( D => n1565, CK => n443, Q => 
                           REGISTERS_31_6_port, QN => n_2049);
   REGISTERS_reg_31_5_inst : DFF_X1 port map( D => n1564, CK => n443, Q => 
                           REGISTERS_31_5_port, QN => n_2050);
   REGISTERS_reg_31_4_inst : DFF_X1 port map( D => n1563, CK => n443, Q => 
                           REGISTERS_31_4_port, QN => n_2051);
   REGISTERS_reg_31_3_inst : DFF_X1 port map( D => n1562, CK => n443, Q => 
                           REGISTERS_31_3_port, QN => n_2052);
   REGISTERS_reg_31_2_inst : DFF_X1 port map( D => n1561, CK => n443, Q => 
                           REGISTERS_31_2_port, QN => n_2053);
   REGISTERS_reg_31_1_inst : DFF_X1 port map( D => n1560, CK => n443, Q => 
                           REGISTERS_31_1_port, QN => n_2054);
   REGISTERS_reg_31_0_inst : DFF_X1 port map( D => n1559, CK => n444, Q => 
                           REGISTERS_31_0_port, QN => n_2055);
   OUT2_reg_31_inst : DFF_X1 port map( D => n1463, CK => n417, Q => n3237, QN 
                           => n_2056);
   OUT2_tri_enable_reg_31_inst : DFF_X1 port map( D => n1558, CK => n516, Q => 
                           n3238, QN => n49);
   OUT2_reg_30_inst : DFF_X1 port map( D => n1464, CK => n418, Q => n3239, QN 
                           => n_2057);
   OUT2_tri_enable_reg_30_inst : DFF_X1 port map( D => n1557, CK => n516, Q => 
                           n3240, QN => n50);
   OUT2_reg_29_inst : DFF_X1 port map( D => n1465, CK => n418, Q => n3241, QN 
                           => n_2058);
   OUT2_tri_enable_reg_29_inst : DFF_X1 port map( D => n1556, CK => n517, Q => 
                           n3242, QN => n51);
   OUT2_reg_28_inst : DFF_X1 port map( D => n1466, CK => n418, Q => n3243, QN 
                           => n_2059);
   OUT2_tri_enable_reg_28_inst : DFF_X1 port map( D => n1555, CK => n517, Q => 
                           n3244, QN => n52);
   OUT2_reg_27_inst : DFF_X1 port map( D => n1467, CK => n418, Q => n3245, QN 
                           => n_2060);
   OUT2_tri_enable_reg_27_inst : DFF_X1 port map( D => n1554, CK => n517, Q => 
                           n3246, QN => n53);
   OUT2_reg_26_inst : DFF_X1 port map( D => n1468, CK => n418, Q => n3247, QN 
                           => n_2061);
   OUT2_tri_enable_reg_26_inst : DFF_X1 port map( D => n1553, CK => n517, Q => 
                           n3248, QN => n54);
   OUT2_reg_25_inst : DFF_X1 port map( D => n1469, CK => n419, Q => n3249, QN 
                           => n_2062);
   OUT2_tri_enable_reg_25_inst : DFF_X1 port map( D => n1552, CK => n517, Q => 
                           n3250, QN => n55);
   OUT2_reg_24_inst : DFF_X1 port map( D => n1470, CK => n419, Q => n3251, QN 
                           => n_2063);
   OUT2_tri_enable_reg_24_inst : DFF_X1 port map( D => n1551, CK => n517, Q => 
                           n3252, QN => n56);
   OUT2_reg_23_inst : DFF_X1 port map( D => n1471, CK => n419, Q => n3253, QN 
                           => n_2064);
   OUT2_tri_enable_reg_23_inst : DFF_X1 port map( D => n1550, CK => n517, Q => 
                           n3254, QN => n57);
   OUT2_reg_22_inst : DFF_X1 port map( D => n1472, CK => n419, Q => n3255, QN 
                           => n_2065);
   OUT2_tri_enable_reg_22_inst : DFF_X1 port map( D => n1549, CK => n517, Q => 
                           n3256, QN => n58);
   OUT2_reg_21_inst : DFF_X1 port map( D => n1473, CK => n419, Q => n3257, QN 
                           => n_2066);
   OUT2_tri_enable_reg_21_inst : DFF_X1 port map( D => n1548, CK => n517, Q => 
                           n3258, QN => n59);
   OUT2_reg_20_inst : DFF_X1 port map( D => n1474, CK => n419, Q => n3259, QN 
                           => n_2067);
   OUT2_tri_enable_reg_20_inst : DFF_X1 port map( D => n1547, CK => n517, Q => 
                           n3260, QN => n60);
   OUT2_reg_19_inst : DFF_X1 port map( D => n1475, CK => n420, Q => n3261, QN 
                           => n_2068);
   OUT2_tri_enable_reg_19_inst : DFF_X1 port map( D => n1546, CK => n517, Q => 
                           n3262, QN => n61);
   OUT2_reg_18_inst : DFF_X1 port map( D => n1476, CK => n420, Q => n3263, QN 
                           => n_2069);
   OUT2_tri_enable_reg_18_inst : DFF_X1 port map( D => n1545, CK => n518, Q => 
                           n3264, QN => n62);
   OUT2_reg_17_inst : DFF_X1 port map( D => n1477, CK => n420, Q => n3265, QN 
                           => n_2070);
   OUT2_tri_enable_reg_17_inst : DFF_X1 port map( D => n1544, CK => n518, Q => 
                           n3266, QN => n63);
   OUT2_reg_16_inst : DFF_X1 port map( D => n1478, CK => n420, Q => n3267, QN 
                           => n_2071);
   OUT2_tri_enable_reg_16_inst : DFF_X1 port map( D => n1543, CK => n518, Q => 
                           n3268, QN => n64);
   OUT2_reg_15_inst : DFF_X1 port map( D => n1479, CK => n420, Q => n3269, QN 
                           => n_2072);
   OUT2_tri_enable_reg_15_inst : DFF_X1 port map( D => n1542, CK => n518, Q => 
                           n3270, QN => n65);
   OUT2_reg_14_inst : DFF_X1 port map( D => n1480, CK => n421, Q => n3271, QN 
                           => n_2073);
   OUT2_tri_enable_reg_14_inst : DFF_X1 port map( D => n1541, CK => n518, Q => 
                           n3272, QN => n66);
   OUT2_reg_13_inst : DFF_X1 port map( D => n1481, CK => n421, Q => n3273, QN 
                           => n_2074);
   OUT2_tri_enable_reg_13_inst : DFF_X1 port map( D => n1540, CK => n518, Q => 
                           n3274, QN => n67);
   OUT2_reg_12_inst : DFF_X1 port map( D => n1482, CK => n421, Q => n3275, QN 
                           => n_2075);
   OUT2_tri_enable_reg_12_inst : DFF_X1 port map( D => n1539, CK => n518, Q => 
                           n3276, QN => n68);
   OUT2_reg_11_inst : DFF_X1 port map( D => n1483, CK => n421, Q => n3277, QN 
                           => n_2076);
   OUT2_tri_enable_reg_11_inst : DFF_X1 port map( D => n1538, CK => n518, Q => 
                           n3278, QN => n69);
   OUT2_reg_10_inst : DFF_X1 port map( D => n1484, CK => n421, Q => n3279, QN 
                           => n_2077);
   OUT2_tri_enable_reg_10_inst : DFF_X1 port map( D => n1537, CK => n518, Q => 
                           n3280, QN => n70);
   OUT2_reg_9_inst : DFF_X1 port map( D => n1485, CK => n421, Q => n3281, QN =>
                           n_2078);
   OUT2_tri_enable_reg_9_inst : DFF_X1 port map( D => n1536, CK => n518, Q => 
                           n3282, QN => n71);
   OUT2_reg_8_inst : DFF_X1 port map( D => n1486, CK => n422, Q => n3283, QN =>
                           n_2079);
   OUT2_tri_enable_reg_8_inst : DFF_X1 port map( D => n1535, CK => n518, Q => 
                           n3284, QN => n72);
   OUT2_reg_7_inst : DFF_X1 port map( D => n1487, CK => n422, Q => n3285, QN =>
                           n_2080);
   OUT2_tri_enable_reg_7_inst : DFF_X1 port map( D => n1534, CK => n519, Q => 
                           n3286, QN => n73);
   OUT2_reg_6_inst : DFF_X1 port map( D => n1488, CK => n422, Q => n3287, QN =>
                           n_2081);
   OUT2_tri_enable_reg_6_inst : DFF_X1 port map( D => n1533, CK => n519, Q => 
                           n3288, QN => n74);
   OUT2_reg_5_inst : DFF_X1 port map( D => n1489, CK => n422, Q => n3289, QN =>
                           n_2082);
   OUT2_tri_enable_reg_5_inst : DFF_X1 port map( D => n1532, CK => n519, Q => 
                           n3290, QN => n75);
   OUT2_reg_4_inst : DFF_X1 port map( D => n1490, CK => n422, Q => n3291, QN =>
                           n_2083);
   OUT2_tri_enable_reg_4_inst : DFF_X1 port map( D => n1531, CK => n519, Q => 
                           n3292, QN => n76);
   OUT2_reg_3_inst : DFF_X1 port map( D => n1491, CK => n423, Q => n3293, QN =>
                           n_2084);
   OUT2_tri_enable_reg_3_inst : DFF_X1 port map( D => n1530, CK => n519, Q => 
                           n3294, QN => n77);
   OUT2_reg_2_inst : DFF_X1 port map( D => n1492, CK => n423, Q => n3295, QN =>
                           n_2085);
   OUT2_tri_enable_reg_2_inst : DFF_X1 port map( D => n1529, CK => n519, Q => 
                           n3296, QN => n78);
   OUT2_reg_1_inst : DFF_X1 port map( D => n1493, CK => n423, Q => n3297, QN =>
                           n_2086);
   OUT2_tri_enable_reg_1_inst : DFF_X1 port map( D => n1528, CK => n519, Q => 
                           n3298, QN => n79);
   OUT2_reg_0_inst : DFF_X1 port map( D => n1494, CK => n423, Q => n3299, QN =>
                           n_2087);
   OUT2_tri_enable_reg_0_inst : DFF_X1 port map( D => n1527, CK => n519, Q => 
                           n3300, QN => n80);
   OUT2_tri_0_inst : TBUF_X1 port map( A => n3299, EN => n3300, Z => OUT2(0));
   OUT2_tri_1_inst : TBUF_X1 port map( A => n3297, EN => n3298, Z => OUT2(1));
   OUT2_tri_2_inst : TBUF_X1 port map( A => n3295, EN => n3296, Z => OUT2(2));
   OUT2_tri_3_inst : TBUF_X1 port map( A => n3293, EN => n3294, Z => OUT2(3));
   OUT2_tri_4_inst : TBUF_X1 port map( A => n3291, EN => n3292, Z => OUT2(4));
   OUT2_tri_5_inst : TBUF_X1 port map( A => n3289, EN => n3290, Z => OUT2(5));
   OUT2_tri_6_inst : TBUF_X1 port map( A => n3287, EN => n3288, Z => OUT2(6));
   OUT2_tri_7_inst : TBUF_X1 port map( A => n3285, EN => n3286, Z => OUT2(7));
   OUT2_tri_8_inst : TBUF_X1 port map( A => n3283, EN => n3284, Z => OUT2(8));
   OUT2_tri_9_inst : TBUF_X1 port map( A => n3281, EN => n3282, Z => OUT2(9));
   OUT2_tri_10_inst : TBUF_X1 port map( A => n3279, EN => n3280, Z => OUT2(10))
                           ;
   OUT2_tri_11_inst : TBUF_X1 port map( A => n3277, EN => n3278, Z => OUT2(11))
                           ;
   OUT2_tri_12_inst : TBUF_X1 port map( A => n3275, EN => n3276, Z => OUT2(12))
                           ;
   OUT2_tri_13_inst : TBUF_X1 port map( A => n3273, EN => n3274, Z => OUT2(13))
                           ;
   OUT2_tri_14_inst : TBUF_X1 port map( A => n3271, EN => n3272, Z => OUT2(14))
                           ;
   OUT2_tri_15_inst : TBUF_X1 port map( A => n3269, EN => n3270, Z => OUT2(15))
                           ;
   OUT2_tri_16_inst : TBUF_X1 port map( A => n3267, EN => n3268, Z => OUT2(16))
                           ;
   OUT2_tri_17_inst : TBUF_X1 port map( A => n3265, EN => n3266, Z => OUT2(17))
                           ;
   OUT2_tri_18_inst : TBUF_X1 port map( A => n3263, EN => n3264, Z => OUT2(18))
                           ;
   OUT2_tri_19_inst : TBUF_X1 port map( A => n3261, EN => n3262, Z => OUT2(19))
                           ;
   OUT2_tri_20_inst : TBUF_X1 port map( A => n3259, EN => n3260, Z => OUT2(20))
                           ;
   OUT2_tri_21_inst : TBUF_X1 port map( A => n3257, EN => n3258, Z => OUT2(21))
                           ;
   OUT2_tri_22_inst : TBUF_X1 port map( A => n3255, EN => n3256, Z => OUT2(22))
                           ;
   OUT2_tri_23_inst : TBUF_X1 port map( A => n3253, EN => n3254, Z => OUT2(23))
                           ;
   OUT2_tri_24_inst : TBUF_X1 port map( A => n3251, EN => n3252, Z => OUT2(24))
                           ;
   OUT2_tri_25_inst : TBUF_X1 port map( A => n3249, EN => n3250, Z => OUT2(25))
                           ;
   OUT2_tri_26_inst : TBUF_X1 port map( A => n3247, EN => n3248, Z => OUT2(26))
                           ;
   OUT2_tri_27_inst : TBUF_X1 port map( A => n3245, EN => n3246, Z => OUT2(27))
                           ;
   OUT2_tri_28_inst : TBUF_X1 port map( A => n3243, EN => n3244, Z => OUT2(28))
                           ;
   OUT2_tri_29_inst : TBUF_X1 port map( A => n3241, EN => n3242, Z => OUT2(29))
                           ;
   OUT2_tri_30_inst : TBUF_X1 port map( A => n3239, EN => n3240, Z => OUT2(30))
                           ;
   OUT2_tri_31_inst : TBUF_X1 port map( A => n3237, EN => n3238, Z => OUT2(31))
                           ;
   OUT1_tri_0_inst : TBUF_X1 port map( A => n3235, EN => n3236, Z => OUT1(0));
   OUT1_tri_1_inst : TBUF_X1 port map( A => n3233, EN => n3234, Z => OUT1(1));
   OUT1_tri_2_inst : TBUF_X1 port map( A => n3231, EN => n3232, Z => OUT1(2));
   OUT1_tri_3_inst : TBUF_X1 port map( A => n3229, EN => n3230, Z => OUT1(3));
   OUT1_tri_4_inst : TBUF_X1 port map( A => n3227, EN => n3228, Z => OUT1(4));
   OUT1_tri_5_inst : TBUF_X1 port map( A => n3225, EN => n3226, Z => OUT1(5));
   OUT1_tri_6_inst : TBUF_X1 port map( A => n3223, EN => n3224, Z => OUT1(6));
   OUT1_tri_7_inst : TBUF_X1 port map( A => n3221, EN => n3222, Z => OUT1(7));
   OUT1_tri_8_inst : TBUF_X1 port map( A => n3219, EN => n3220, Z => OUT1(8));
   OUT1_tri_9_inst : TBUF_X1 port map( A => n3217, EN => n3218, Z => OUT1(9));
   OUT1_tri_10_inst : TBUF_X1 port map( A => n3215, EN => n3216, Z => OUT1(10))
                           ;
   OUT1_tri_11_inst : TBUF_X1 port map( A => n3213, EN => n3214, Z => OUT1(11))
                           ;
   OUT1_tri_12_inst : TBUF_X1 port map( A => n3211, EN => n3212, Z => OUT1(12))
                           ;
   OUT1_tri_13_inst : TBUF_X1 port map( A => n3209, EN => n3210, Z => OUT1(13))
                           ;
   OUT1_tri_14_inst : TBUF_X1 port map( A => n3207, EN => n3208, Z => OUT1(14))
                           ;
   OUT1_tri_15_inst : TBUF_X1 port map( A => n3205, EN => n3206, Z => OUT1(15))
                           ;
   OUT1_tri_16_inst : TBUF_X1 port map( A => n3203, EN => n3204, Z => OUT1(16))
                           ;
   OUT1_tri_17_inst : TBUF_X1 port map( A => n3201, EN => n3202, Z => OUT1(17))
                           ;
   OUT1_tri_18_inst : TBUF_X1 port map( A => n3199, EN => n3200, Z => OUT1(18))
                           ;
   OUT1_tri_19_inst : TBUF_X1 port map( A => n3197, EN => n3198, Z => OUT1(19))
                           ;
   OUT1_tri_20_inst : TBUF_X1 port map( A => n3195, EN => n3196, Z => OUT1(20))
                           ;
   OUT1_tri_21_inst : TBUF_X1 port map( A => n3193, EN => n3194, Z => OUT1(21))
                           ;
   OUT1_tri_22_inst : TBUF_X1 port map( A => n3191, EN => n3192, Z => OUT1(22))
                           ;
   OUT1_tri_23_inst : TBUF_X1 port map( A => n3189, EN => n3190, Z => OUT1(23))
                           ;
   OUT1_tri_24_inst : TBUF_X1 port map( A => n3187, EN => n3188, Z => OUT1(24))
                           ;
   OUT1_tri_25_inst : TBUF_X1 port map( A => n3185, EN => n3186, Z => OUT1(25))
                           ;
   OUT1_tri_26_inst : TBUF_X1 port map( A => n3183, EN => n3184, Z => OUT1(26))
                           ;
   OUT1_tri_27_inst : TBUF_X1 port map( A => n3181, EN => n3182, Z => OUT1(27))
                           ;
   OUT1_tri_28_inst : TBUF_X1 port map( A => n3179, EN => n3180, Z => OUT1(28))
                           ;
   OUT1_tri_29_inst : TBUF_X1 port map( A => n3177, EN => n3178, Z => OUT1(29))
                           ;
   OUT1_tri_30_inst : TBUF_X1 port map( A => n3175, EN => n3176, Z => OUT1(30))
                           ;
   OUT1_tri_31_inst : TBUF_X1 port map( A => n3173, EN => n3174, Z => OUT1(31))
                           ;
   U3 : AND2_X1 port map( A1 => ADD_RD1(0), A2 => n567, ZN => n1);
   U4 : AND2_X1 port map( A1 => ADD_RD2(0), A2 => n1251, ZN => n2);
   U5 : AND2_X1 port map( A1 => n567, A2 => n1246, ZN => n3);
   U6 : AND2_X1 port map( A1 => n1251, A2 => n3082, ZN => n4);
   U7 : AND2_X1 port map( A1 => n566, A2 => ADD_RD1(0), ZN => n5);
   U8 : AND2_X1 port map( A1 => n569, A2 => ADD_RD1(0), ZN => n6);
   U9 : AND2_X1 port map( A1 => n568, A2 => ADD_RD1(0), ZN => n7);
   U10 : AND2_X1 port map( A1 => n566, A2 => n1246, ZN => n8);
   U11 : AND2_X1 port map( A1 => n569, A2 => n1246, ZN => n9);
   U12 : AND2_X1 port map( A1 => n568, A2 => n1246, ZN => n10);
   U13 : AND2_X1 port map( A1 => n1250, A2 => ADD_RD2(0), ZN => n11);
   U14 : AND2_X1 port map( A1 => n1253, A2 => ADD_RD2(0), ZN => n12);
   U15 : AND2_X1 port map( A1 => n1252, A2 => ADD_RD2(0), ZN => n13);
   U16 : AND2_X1 port map( A1 => n1250, A2 => n3082, ZN => n14);
   U17 : AND2_X1 port map( A1 => n1253, A2 => n3082, ZN => n15);
   U18 : AND2_X1 port map( A1 => n1252, A2 => n3082, ZN => n16);
   U19 : OR2_X2 port map( A1 => RD1, A2 => n3088, ZN => n3087);
   U20 : OR2_X2 port map( A1 => RD2, A2 => n3088, ZN => n3172);
   U21 : INV_X1 port map( A => n3159, ZN => n81);
   U22 : INV_X2 port map( A => n81, ZN => n82);
   U23 : INV_X1 port map( A => n3160, ZN => n83);
   U24 : INV_X2 port map( A => n83, ZN => n84);
   U25 : INV_X1 port map( A => n3165, ZN => n85);
   U26 : INV_X2 port map( A => n85, ZN => n86);
   U27 : INV_X1 port map( A => n3166, ZN => n87);
   U28 : INV_X2 port map( A => n87, ZN => n88);
   U29 : INV_X1 port map( A => n3167, ZN => n89);
   U30 : INV_X2 port map( A => n89, ZN => n90);
   U31 : INV_X1 port map( A => n3168, ZN => n91);
   U32 : INV_X2 port map( A => n91, ZN => n92);
   U33 : INV_X1 port map( A => n3169, ZN => n93);
   U34 : INV_X2 port map( A => n93, ZN => n94);
   U35 : INV_X1 port map( A => n3170, ZN => n95);
   U36 : INV_X2 port map( A => n95, ZN => n96);
   U37 : INV_X1 port map( A => n3171, ZN => n97);
   U38 : INV_X2 port map( A => n97, ZN => n98);
   U39 : INV_X1 port map( A => n3157, ZN => n99);
   U40 : INV_X2 port map( A => n99, ZN => n100);
   U41 : INV_X1 port map( A => n3158, ZN => n101);
   U42 : INV_X2 port map( A => n101, ZN => n102);
   U43 : INV_X1 port map( A => n3155, ZN => n103);
   U44 : INV_X2 port map( A => n103, ZN => n104);
   U45 : INV_X1 port map( A => n3156, ZN => n105);
   U46 : INV_X2 port map( A => n105, ZN => n106);
   U47 : INV_X1 port map( A => n3153, ZN => n107);
   U48 : INV_X2 port map( A => n107, ZN => n108);
   U49 : INV_X1 port map( A => n3154, ZN => n109);
   U50 : INV_X2 port map( A => n109, ZN => n110);
   U51 : INV_X1 port map( A => n3150, ZN => n111);
   U52 : INV_X2 port map( A => n111, ZN => n112);
   U53 : INV_X1 port map( A => n3151, ZN => n113);
   U54 : INV_X2 port map( A => n113, ZN => n114);
   U55 : INV_X1 port map( A => n3148, ZN => n115);
   U56 : INV_X2 port map( A => n115, ZN => n116);
   U57 : INV_X1 port map( A => n3149, ZN => n117);
   U58 : INV_X2 port map( A => n117, ZN => n118);
   U59 : INV_X1 port map( A => n3146, ZN => n119);
   U60 : INV_X2 port map( A => n119, ZN => n120);
   U61 : INV_X1 port map( A => n3147, ZN => n121);
   U62 : INV_X2 port map( A => n121, ZN => n122);
   U63 : INV_X1 port map( A => n3144, ZN => n123);
   U64 : INV_X2 port map( A => n123, ZN => n124);
   U65 : INV_X1 port map( A => n3145, ZN => n125);
   U66 : INV_X2 port map( A => n125, ZN => n126);
   U67 : INV_X1 port map( A => n3137, ZN => n127);
   U68 : INV_X2 port map( A => n127, ZN => n128);
   U69 : INV_X1 port map( A => n3142, ZN => n129);
   U70 : INV_X2 port map( A => n129, ZN => n130);
   U71 : INV_X1 port map( A => n3133, ZN => n131);
   U72 : INV_X2 port map( A => n131, ZN => n132);
   U73 : INV_X1 port map( A => n3135, ZN => n133);
   U74 : INV_X2 port map( A => n133, ZN => n134);
   U75 : INV_X1 port map( A => n3129, ZN => n135);
   U76 : INV_X2 port map( A => n135, ZN => n136);
   U77 : INV_X1 port map( A => n3131, ZN => n137);
   U78 : INV_X2 port map( A => n137, ZN => n138);
   U79 : INV_X1 port map( A => n3125, ZN => n139);
   U80 : INV_X2 port map( A => n139, ZN => n140);
   U81 : INV_X1 port map( A => n3127, ZN => n141);
   U82 : INV_X2 port map( A => n141, ZN => n142);
   U83 : OAI21_X4 port map( B1 => n3122, B2 => n3123, A => n3124, ZN => n3090);
   U84 : INV_X4 port map( A => RESET, ZN => n3124);
   U85 : INV_X4 port map( A => n3088, ZN => n3086);
   U86 : NAND2_X4 port map( A1 => ENABLE, A2 => n3124, ZN => n3088);
   U87 : NAND2_X2 port map( A1 => ADD_RD1(4), A2 => ADD_RD1(3), ZN => n1242);
   U88 : NAND2_X2 port map( A1 => ADD_RD2(4), A2 => ADD_RD2(3), ZN => n3078);
   U89 : NAND2_X2 port map( A1 => ADD_RD1(4), A2 => n1249, ZN => n1244);
   U90 : NAND2_X2 port map( A1 => ADD_RD2(4), A2 => n3085, ZN => n3080);
   U91 : NOR2_X4 port map( A1 => n1249, A2 => ADD_RD1(4), ZN => n1238);
   U92 : NOR2_X4 port map( A1 => n3085, A2 => ADD_RD2(4), ZN => n3074);
   U93 : NOR2_X4 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(4), ZN => n1240);
   U94 : NOR2_X4 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(4), ZN => n3076);
   U95 : BUF_X1 port map( A => n413, Z => n411);
   U96 : BUF_X1 port map( A => n396, Z => n394);
   U97 : BUF_X1 port map( A => n379, Z => n377);
   U98 : BUF_X1 port map( A => n362, Z => n360);
   U99 : BUF_X1 port map( A => n413, Z => n410);
   U100 : BUF_X1 port map( A => n396, Z => n393);
   U101 : BUF_X1 port map( A => n379, Z => n376);
   U102 : BUF_X1 port map( A => n362, Z => n359);
   U103 : BUF_X1 port map( A => n277, Z => n275);
   U104 : BUF_X1 port map( A => n260, Z => n258);
   U105 : BUF_X1 port map( A => n243, Z => n241);
   U106 : BUF_X1 port map( A => n226, Z => n224);
   U107 : BUF_X1 port map( A => n277, Z => n274);
   U108 : BUF_X1 port map( A => n260, Z => n257);
   U109 : BUF_X1 port map( A => n243, Z => n240);
   U110 : BUF_X1 port map( A => n226, Z => n223);
   U111 : BUF_X1 port map( A => n563, Z => n557);
   U112 : BUF_X1 port map( A => n563, Z => n556);
   U113 : BUF_X1 port map( A => n562, Z => n560);
   U114 : BUF_X1 port map( A => n562, Z => n559);
   U115 : BUF_X1 port map( A => n563, Z => n558);
   U116 : BUF_X1 port map( A => n562, Z => n561);
   U117 : BUF_X1 port map( A => n16, Z => n413);
   U118 : BUF_X1 port map( A => n15, Z => n396);
   U119 : BUF_X1 port map( A => n14, Z => n379);
   U120 : BUF_X1 port map( A => n4, Z => n362);
   U121 : BUF_X1 port map( A => n10, Z => n277);
   U122 : BUF_X1 port map( A => n9, Z => n260);
   U123 : BUF_X1 port map( A => n8, Z => n243);
   U124 : BUF_X1 port map( A => n3, Z => n226);
   U125 : BUF_X1 port map( A => n345, Z => n343);
   U126 : BUF_X1 port map( A => n328, Z => n326);
   U127 : BUF_X1 port map( A => n311, Z => n309);
   U128 : BUF_X1 port map( A => n294, Z => n292);
   U129 : BUF_X1 port map( A => n345, Z => n342);
   U130 : BUF_X1 port map( A => n328, Z => n325);
   U131 : BUF_X1 port map( A => n311, Z => n308);
   U132 : BUF_X1 port map( A => n294, Z => n291);
   U133 : BUF_X1 port map( A => n209_port, Z => n207_port);
   U134 : BUF_X1 port map( A => n192_port, Z => n190_port);
   U135 : BUF_X1 port map( A => n175_port, Z => n173_port);
   U136 : BUF_X1 port map( A => n158_port, Z => n156_port);
   U137 : BUF_X1 port map( A => n209_port, Z => n206_port);
   U138 : BUF_X1 port map( A => n192_port, Z => n189_port);
   U139 : BUF_X1 port map( A => n175_port, Z => n172_port);
   U140 : BUF_X1 port map( A => n158_port, Z => n155);
   U141 : BUF_X1 port map( A => n414, Z => n409);
   U142 : BUF_X1 port map( A => n397, Z => n392);
   U143 : BUF_X1 port map( A => n380, Z => n375);
   U144 : BUF_X1 port map( A => n363, Z => n358);
   U145 : BUF_X1 port map( A => n278, Z => n273);
   U146 : BUF_X1 port map( A => n261, Z => n256);
   U147 : BUF_X1 port map( A => n244, Z => n239);
   U148 : BUF_X1 port map( A => n227, Z => n222);
   U149 : BUF_X1 port map( A => n564, Z => n555);
   U150 : BUF_X1 port map( A => n565, Z => n563);
   U151 : BUF_X1 port map( A => n565, Z => n562);
   U152 : BUF_X1 port map( A => n13, Z => n345);
   U153 : BUF_X1 port map( A => n12, Z => n328);
   U154 : BUF_X1 port map( A => n11, Z => n311);
   U155 : BUF_X1 port map( A => n2, Z => n294);
   U156 : BUF_X1 port map( A => n7, Z => n209_port);
   U157 : BUF_X1 port map( A => n6, Z => n192_port);
   U158 : BUF_X1 port map( A => n5, Z => n175_port);
   U159 : BUF_X1 port map( A => n1, Z => n158_port);
   U160 : BUF_X1 port map( A => n346, Z => n341);
   U161 : BUF_X1 port map( A => n329, Z => n324);
   U162 : BUF_X1 port map( A => n312, Z => n307);
   U163 : BUF_X1 port map( A => n295, Z => n290);
   U164 : BUF_X1 port map( A => n210_port, Z => n205_port);
   U165 : BUF_X1 port map( A => n193_port, Z => n188);
   U166 : BUF_X1 port map( A => n176_port, Z => n171_port);
   U167 : BUF_X1 port map( A => n159_port, Z => n154);
   U168 : BUF_X1 port map( A => CLK, Z => n565);
   U169 : BUF_X1 port map( A => n411, Z => n400);
   U170 : BUF_X1 port map( A => n377, Z => n366);
   U171 : BUF_X1 port map( A => n411, Z => n401);
   U172 : BUF_X1 port map( A => n377, Z => n367);
   U173 : BUF_X1 port map( A => n411, Z => n402);
   U174 : BUF_X1 port map( A => n377, Z => n368);
   U175 : BUF_X1 port map( A => n410, Z => n403);
   U176 : BUF_X1 port map( A => n376, Z => n369);
   U177 : BUF_X1 port map( A => n410, Z => n404);
   U178 : BUF_X1 port map( A => n376, Z => n370);
   U179 : BUF_X1 port map( A => n410, Z => n405);
   U180 : BUF_X1 port map( A => n376, Z => n371);
   U181 : BUF_X1 port map( A => n275, Z => n264);
   U182 : BUF_X1 port map( A => n241, Z => n230);
   U183 : BUF_X1 port map( A => n275, Z => n265);
   U184 : BUF_X1 port map( A => n241, Z => n231);
   U185 : BUF_X1 port map( A => n275, Z => n266);
   U186 : BUF_X1 port map( A => n241, Z => n232);
   U187 : BUF_X1 port map( A => n274, Z => n267);
   U188 : BUF_X1 port map( A => n240, Z => n233);
   U189 : BUF_X1 port map( A => n274, Z => n268);
   U190 : BUF_X1 port map( A => n240, Z => n234);
   U191 : BUF_X1 port map( A => n274, Z => n269);
   U192 : BUF_X1 port map( A => n240, Z => n235);
   U193 : BUF_X1 port map( A => n520, Z => n518);
   U194 : BUF_X1 port map( A => n520, Z => n517);
   U195 : BUF_X1 port map( A => n545, Z => n443);
   U196 : BUF_X1 port map( A => n545, Z => n442);
   U197 : BUF_X1 port map( A => n546, Z => n441);
   U198 : BUF_X1 port map( A => n546, Z => n440);
   U199 : BUF_X1 port map( A => n546, Z => n439);
   U200 : BUF_X1 port map( A => n547, Z => n438);
   U201 : BUF_X1 port map( A => n547, Z => n437);
   U202 : BUF_X1 port map( A => n547, Z => n436);
   U203 : BUF_X1 port map( A => n548, Z => n435);
   U204 : BUF_X1 port map( A => n548, Z => n434);
   U205 : BUF_X1 port map( A => n548, Z => n433);
   U206 : BUF_X1 port map( A => n549, Z => n432);
   U207 : BUF_X1 port map( A => n549, Z => n431);
   U208 : BUF_X1 port map( A => n549, Z => n430);
   U209 : BUF_X1 port map( A => n537, Z => n466);
   U210 : BUF_X1 port map( A => n538, Z => n465);
   U211 : BUF_X1 port map( A => n538, Z => n464);
   U212 : BUF_X1 port map( A => n538, Z => n463);
   U213 : BUF_X1 port map( A => n539, Z => n462);
   U214 : BUF_X1 port map( A => n539, Z => n461);
   U215 : BUF_X1 port map( A => n539, Z => n460);
   U216 : BUF_X1 port map( A => n540, Z => n459);
   U217 : BUF_X1 port map( A => n540, Z => n458);
   U218 : BUF_X1 port map( A => n540, Z => n457);
   U219 : BUF_X1 port map( A => n541, Z => n456);
   U220 : BUF_X1 port map( A => n541, Z => n455);
   U221 : BUF_X1 port map( A => n541, Z => n454);
   U222 : BUF_X1 port map( A => n542, Z => n453);
   U223 : BUF_X1 port map( A => n542, Z => n452);
   U224 : BUF_X1 port map( A => n542, Z => n451);
   U225 : BUF_X1 port map( A => n543, Z => n450);
   U226 : BUF_X1 port map( A => n543, Z => n449);
   U227 : BUF_X1 port map( A => n543, Z => n448);
   U228 : BUF_X1 port map( A => n544, Z => n447);
   U229 : BUF_X1 port map( A => n544, Z => n446);
   U230 : BUF_X1 port map( A => n544, Z => n445);
   U231 : BUF_X1 port map( A => n545, Z => n444);
   U232 : BUF_X1 port map( A => n522, Z => n512);
   U233 : BUF_X1 port map( A => n522, Z => n511);
   U234 : BUF_X1 port map( A => n523, Z => n510);
   U235 : BUF_X1 port map( A => n523, Z => n509);
   U236 : BUF_X1 port map( A => n523, Z => n508);
   U237 : BUF_X1 port map( A => n524, Z => n507);
   U238 : BUF_X1 port map( A => n524, Z => n506);
   U239 : BUF_X1 port map( A => n524, Z => n505);
   U240 : BUF_X1 port map( A => n525, Z => n504);
   U241 : BUF_X1 port map( A => n525, Z => n503);
   U242 : BUF_X1 port map( A => n525, Z => n502);
   U243 : BUF_X1 port map( A => n526, Z => n501);
   U244 : BUF_X1 port map( A => n526, Z => n500);
   U245 : BUF_X1 port map( A => n526, Z => n499);
   U246 : BUF_X1 port map( A => n527, Z => n498);
   U247 : BUF_X1 port map( A => n527, Z => n497);
   U248 : BUF_X1 port map( A => n527, Z => n496);
   U249 : BUF_X1 port map( A => n528, Z => n495);
   U250 : BUF_X1 port map( A => n528, Z => n494);
   U251 : BUF_X1 port map( A => n528, Z => n493);
   U252 : BUF_X1 port map( A => n529, Z => n492);
   U253 : BUF_X1 port map( A => n529, Z => n491);
   U254 : BUF_X1 port map( A => n529, Z => n490);
   U255 : BUF_X1 port map( A => n530, Z => n489);
   U256 : BUF_X1 port map( A => n530, Z => n488);
   U257 : BUF_X1 port map( A => n530, Z => n487);
   U258 : BUF_X1 port map( A => n531, Z => n486);
   U259 : BUF_X1 port map( A => n531, Z => n485);
   U260 : BUF_X1 port map( A => n531, Z => n484);
   U261 : BUF_X1 port map( A => n532, Z => n483);
   U262 : BUF_X1 port map( A => n532, Z => n482);
   U263 : BUF_X1 port map( A => n532, Z => n481);
   U264 : BUF_X1 port map( A => n533, Z => n480);
   U265 : BUF_X1 port map( A => n533, Z => n479);
   U266 : BUF_X1 port map( A => n533, Z => n478);
   U267 : BUF_X1 port map( A => n534, Z => n477);
   U268 : BUF_X1 port map( A => n534, Z => n476);
   U269 : BUF_X1 port map( A => n534, Z => n475);
   U270 : BUF_X1 port map( A => n535, Z => n474);
   U271 : BUF_X1 port map( A => n535, Z => n473);
   U272 : BUF_X1 port map( A => n535, Z => n472);
   U273 : BUF_X1 port map( A => n536, Z => n471);
   U274 : BUF_X1 port map( A => n536, Z => n470);
   U275 : BUF_X1 port map( A => n536, Z => n469);
   U276 : BUF_X1 port map( A => n537, Z => n468);
   U277 : BUF_X1 port map( A => n537, Z => n467);
   U278 : BUF_X1 port map( A => n521, Z => n516);
   U279 : BUF_X1 port map( A => n521, Z => n515);
   U280 : BUF_X1 port map( A => n521, Z => n514);
   U281 : BUF_X1 port map( A => n522, Z => n513);
   U282 : BUF_X1 port map( A => n412, Z => n398);
   U283 : BUF_X1 port map( A => n378, Z => n364);
   U284 : BUF_X1 port map( A => n412, Z => n399);
   U285 : BUF_X1 port map( A => n378, Z => n365);
   U286 : BUF_X1 port map( A => n276, Z => n262);
   U287 : BUF_X1 port map( A => n242, Z => n228);
   U288 : BUF_X1 port map( A => n276, Z => n263);
   U289 : BUF_X1 port map( A => n242, Z => n229);
   U290 : BUF_X1 port map( A => n394, Z => n383);
   U291 : BUF_X1 port map( A => n360, Z => n349);
   U292 : BUF_X1 port map( A => n394, Z => n384);
   U293 : BUF_X1 port map( A => n360, Z => n350);
   U294 : BUF_X1 port map( A => n394, Z => n385);
   U295 : BUF_X1 port map( A => n360, Z => n351);
   U296 : BUF_X1 port map( A => n393, Z => n386);
   U297 : BUF_X1 port map( A => n359, Z => n352);
   U298 : BUF_X1 port map( A => n393, Z => n387);
   U299 : BUF_X1 port map( A => n359, Z => n353);
   U300 : BUF_X1 port map( A => n393, Z => n388);
   U301 : BUF_X1 port map( A => n359, Z => n354);
   U302 : BUF_X1 port map( A => n258, Z => n247);
   U303 : BUF_X1 port map( A => n224, Z => n213_port);
   U304 : BUF_X1 port map( A => n258, Z => n248);
   U305 : BUF_X1 port map( A => n224, Z => n214_port);
   U306 : BUF_X1 port map( A => n258, Z => n249);
   U307 : BUF_X1 port map( A => n224, Z => n215_port);
   U308 : BUF_X1 port map( A => n257, Z => n250);
   U309 : BUF_X1 port map( A => n223, Z => n216_port);
   U310 : BUF_X1 port map( A => n257, Z => n251);
   U311 : BUF_X1 port map( A => n223, Z => n217_port);
   U312 : BUF_X1 port map( A => n257, Z => n252);
   U313 : BUF_X1 port map( A => n223, Z => n218_port);
   U314 : BUF_X1 port map( A => n395, Z => n381);
   U315 : BUF_X1 port map( A => n361, Z => n347);
   U316 : BUF_X1 port map( A => n395, Z => n382);
   U317 : BUF_X1 port map( A => n361, Z => n348);
   U318 : BUF_X1 port map( A => n259, Z => n245);
   U319 : BUF_X1 port map( A => n225, Z => n211_port);
   U320 : BUF_X1 port map( A => n259, Z => n246);
   U321 : BUF_X1 port map( A => n225, Z => n212_port);
   U322 : BUF_X1 port map( A => n520, Z => n519);
   U323 : BUF_X1 port map( A => n561, Z => n520);
   U324 : BUF_X1 port map( A => n556, Z => n546);
   U325 : BUF_X1 port map( A => n556, Z => n547);
   U326 : BUF_X1 port map( A => n556, Z => n548);
   U327 : BUF_X1 port map( A => n556, Z => n549);
   U328 : BUF_X1 port map( A => n558, Z => n538);
   U329 : BUF_X1 port map( A => n558, Z => n539);
   U330 : BUF_X1 port map( A => n557, Z => n540);
   U331 : BUF_X1 port map( A => n557, Z => n541);
   U332 : BUF_X1 port map( A => n557, Z => n542);
   U333 : BUF_X1 port map( A => n557, Z => n543);
   U334 : BUF_X1 port map( A => n557, Z => n544);
   U335 : BUF_X1 port map( A => n556, Z => n545);
   U336 : BUF_X1 port map( A => n561, Z => n523);
   U337 : BUF_X1 port map( A => n561, Z => n524);
   U338 : BUF_X1 port map( A => n560, Z => n525);
   U339 : BUF_X1 port map( A => n560, Z => n526);
   U340 : BUF_X1 port map( A => n560, Z => n527);
   U341 : BUF_X1 port map( A => n560, Z => n528);
   U342 : BUF_X1 port map( A => n560, Z => n529);
   U343 : BUF_X1 port map( A => n559, Z => n530);
   U344 : BUF_X1 port map( A => n559, Z => n531);
   U345 : BUF_X1 port map( A => n559, Z => n532);
   U346 : BUF_X1 port map( A => n559, Z => n533);
   U347 : BUF_X1 port map( A => n559, Z => n534);
   U348 : BUF_X1 port map( A => n558, Z => n535);
   U349 : BUF_X1 port map( A => n558, Z => n536);
   U350 : BUF_X1 port map( A => n558, Z => n537);
   U351 : BUF_X1 port map( A => n561, Z => n521);
   U352 : BUF_X1 port map( A => n561, Z => n522);
   U353 : BUF_X1 port map( A => n413, Z => n412);
   U354 : BUF_X1 port map( A => n396, Z => n395);
   U355 : BUF_X1 port map( A => n379, Z => n378);
   U356 : BUF_X1 port map( A => n362, Z => n361);
   U357 : BUF_X1 port map( A => n277, Z => n276);
   U358 : BUF_X1 port map( A => n260, Z => n259);
   U359 : BUF_X1 port map( A => n243, Z => n242);
   U360 : BUF_X1 port map( A => n226, Z => n225);
   U361 : BUF_X1 port map( A => n343, Z => n332);
   U362 : BUF_X1 port map( A => n309, Z => n298);
   U363 : BUF_X1 port map( A => n343, Z => n333);
   U364 : BUF_X1 port map( A => n309, Z => n299);
   U365 : BUF_X1 port map( A => n343, Z => n334);
   U366 : BUF_X1 port map( A => n309, Z => n300);
   U367 : BUF_X1 port map( A => n342, Z => n335);
   U368 : BUF_X1 port map( A => n308, Z => n301);
   U369 : BUF_X1 port map( A => n342, Z => n336);
   U370 : BUF_X1 port map( A => n308, Z => n302);
   U371 : BUF_X1 port map( A => n342, Z => n337);
   U372 : BUF_X1 port map( A => n308, Z => n303);
   U373 : BUF_X1 port map( A => n207_port, Z => n196_port);
   U374 : BUF_X1 port map( A => n173_port, Z => n162_port);
   U375 : BUF_X1 port map( A => n207_port, Z => n197_port);
   U376 : BUF_X1 port map( A => n173_port, Z => n163_port);
   U377 : BUF_X1 port map( A => n207_port, Z => n198_port);
   U378 : BUF_X1 port map( A => n173_port, Z => n164_port);
   U379 : BUF_X1 port map( A => n206_port, Z => n199_port);
   U380 : BUF_X1 port map( A => n172_port, Z => n165_port);
   U381 : BUF_X1 port map( A => n206_port, Z => n200_port);
   U382 : BUF_X1 port map( A => n172_port, Z => n166_port);
   U383 : BUF_X1 port map( A => n206_port, Z => n201_port);
   U384 : BUF_X1 port map( A => n172_port, Z => n167_port);
   U385 : BUF_X1 port map( A => n409, Z => n406);
   U386 : BUF_X1 port map( A => n375, Z => n372);
   U387 : BUF_X1 port map( A => n409, Z => n407);
   U388 : BUF_X1 port map( A => n375, Z => n373);
   U389 : BUF_X1 port map( A => n273, Z => n270);
   U390 : BUF_X1 port map( A => n239, Z => n236);
   U391 : BUF_X1 port map( A => n273, Z => n271);
   U392 : BUF_X1 port map( A => n239, Z => n237);
   U393 : BUF_X1 port map( A => n550, Z => n429);
   U394 : BUF_X1 port map( A => n550, Z => n428);
   U395 : BUF_X1 port map( A => n550, Z => n427);
   U396 : BUF_X1 port map( A => n551, Z => n426);
   U397 : BUF_X1 port map( A => n551, Z => n425);
   U398 : BUF_X1 port map( A => n551, Z => n424);
   U399 : BUF_X1 port map( A => n552, Z => n423);
   U400 : BUF_X1 port map( A => n552, Z => n422);
   U401 : BUF_X1 port map( A => n552, Z => n421);
   U402 : BUF_X1 port map( A => n553, Z => n420);
   U403 : BUF_X1 port map( A => n553, Z => n419);
   U404 : BUF_X1 port map( A => n553, Z => n418);
   U405 : BUF_X1 port map( A => n554, Z => n417);
   U406 : BUF_X1 port map( A => n554, Z => n416);
   U407 : BUF_X1 port map( A => n554, Z => n415);
   U408 : BUF_X1 port map( A => n344, Z => n330);
   U409 : BUF_X1 port map( A => n310, Z => n296);
   U410 : BUF_X1 port map( A => n344, Z => n331);
   U411 : BUF_X1 port map( A => n310, Z => n297);
   U412 : BUF_X1 port map( A => n208_port, Z => n194_port);
   U413 : BUF_X1 port map( A => n174_port, Z => n160_port);
   U414 : BUF_X1 port map( A => n208_port, Z => n195_port);
   U415 : BUF_X1 port map( A => n174_port, Z => n161_port);
   U416 : BUF_X1 port map( A => n326, Z => n315);
   U417 : BUF_X1 port map( A => n292, Z => n281);
   U418 : BUF_X1 port map( A => n326, Z => n316);
   U419 : BUF_X1 port map( A => n292, Z => n282);
   U420 : BUF_X1 port map( A => n326, Z => n317);
   U421 : BUF_X1 port map( A => n292, Z => n283);
   U422 : BUF_X1 port map( A => n325, Z => n318);
   U423 : BUF_X1 port map( A => n291, Z => n284);
   U424 : BUF_X1 port map( A => n325, Z => n319);
   U425 : BUF_X1 port map( A => n291, Z => n285);
   U426 : BUF_X1 port map( A => n325, Z => n320);
   U427 : BUF_X1 port map( A => n291, Z => n286);
   U428 : BUF_X1 port map( A => n392, Z => n389);
   U429 : BUF_X1 port map( A => n358, Z => n355);
   U430 : BUF_X1 port map( A => n392, Z => n390);
   U431 : BUF_X1 port map( A => n358, Z => n356);
   U432 : BUF_X1 port map( A => n190_port, Z => n179_port);
   U433 : BUF_X1 port map( A => n156_port, Z => n145);
   U434 : BUF_X1 port map( A => n190_port, Z => n180_port);
   U435 : BUF_X1 port map( A => n156_port, Z => n146);
   U436 : BUF_X1 port map( A => n190_port, Z => n181_port);
   U437 : BUF_X1 port map( A => n156_port, Z => n147);
   U438 : BUF_X1 port map( A => n189_port, Z => n182_port);
   U439 : BUF_X1 port map( A => n155, Z => n148);
   U440 : BUF_X1 port map( A => n189_port, Z => n183_port);
   U441 : BUF_X1 port map( A => n155, Z => n149);
   U442 : BUF_X1 port map( A => n189_port, Z => n184_port);
   U443 : BUF_X1 port map( A => n155, Z => n150);
   U444 : BUF_X1 port map( A => n256, Z => n253);
   U445 : BUF_X1 port map( A => n222, Z => n219_port);
   U446 : BUF_X1 port map( A => n256, Z => n254);
   U447 : BUF_X1 port map( A => n222, Z => n220_port);
   U448 : BUF_X1 port map( A => n327, Z => n313);
   U449 : BUF_X1 port map( A => n293, Z => n279);
   U450 : BUF_X1 port map( A => n327, Z => n314);
   U451 : BUF_X1 port map( A => n293, Z => n280);
   U452 : BUF_X1 port map( A => n191_port, Z => n177_port);
   U453 : BUF_X1 port map( A => n157_port, Z => n143);
   U454 : BUF_X1 port map( A => n191_port, Z => n178_port);
   U455 : BUF_X1 port map( A => n157_port, Z => n144);
   U456 : BUF_X1 port map( A => n409, Z => n408);
   U457 : BUF_X1 port map( A => n375, Z => n374);
   U458 : BUF_X1 port map( A => n273, Z => n272);
   U459 : BUF_X1 port map( A => n239, Z => n238);
   U460 : BUF_X1 port map( A => n392, Z => n391);
   U461 : BUF_X1 port map( A => n358, Z => n357);
   U462 : BUF_X1 port map( A => n256, Z => n255);
   U463 : BUF_X1 port map( A => n222, Z => n221);
   U464 : BUF_X1 port map( A => n16, Z => n414);
   U465 : BUF_X1 port map( A => n15, Z => n397);
   U466 : BUF_X1 port map( A => n14, Z => n380);
   U467 : BUF_X1 port map( A => n4, Z => n363);
   U468 : BUF_X1 port map( A => n10, Z => n278);
   U469 : BUF_X1 port map( A => n9, Z => n261);
   U470 : BUF_X1 port map( A => n8, Z => n244);
   U471 : BUF_X1 port map( A => n3, Z => n227);
   U472 : BUF_X1 port map( A => n555, Z => n550);
   U473 : BUF_X1 port map( A => n555, Z => n551);
   U474 : BUF_X1 port map( A => n555, Z => n552);
   U475 : BUF_X1 port map( A => n555, Z => n553);
   U476 : BUF_X1 port map( A => n555, Z => n554);
   U477 : BUF_X1 port map( A => n345, Z => n344);
   U478 : BUF_X1 port map( A => n328, Z => n327);
   U479 : BUF_X1 port map( A => n311, Z => n310);
   U480 : BUF_X1 port map( A => n294, Z => n293);
   U481 : BUF_X1 port map( A => n209_port, Z => n208_port);
   U482 : BUF_X1 port map( A => n192_port, Z => n191_port);
   U483 : BUF_X1 port map( A => n175_port, Z => n174_port);
   U484 : BUF_X1 port map( A => n158_port, Z => n157_port);
   U485 : BUF_X1 port map( A => n341, Z => n338);
   U486 : BUF_X1 port map( A => n307, Z => n304);
   U487 : BUF_X1 port map( A => n341, Z => n339);
   U488 : BUF_X1 port map( A => n307, Z => n305);
   U489 : BUF_X1 port map( A => n205_port, Z => n202_port);
   U490 : BUF_X1 port map( A => n171_port, Z => n168_port);
   U491 : BUF_X1 port map( A => n205_port, Z => n203_port);
   U492 : BUF_X1 port map( A => n171_port, Z => n169_port);
   U493 : BUF_X1 port map( A => n324, Z => n321);
   U494 : BUF_X1 port map( A => n290, Z => n287);
   U495 : BUF_X1 port map( A => n324, Z => n322);
   U496 : BUF_X1 port map( A => n290, Z => n288);
   U497 : BUF_X1 port map( A => n188, Z => n185_port);
   U498 : BUF_X1 port map( A => n154, Z => n151);
   U499 : BUF_X1 port map( A => n188, Z => n186_port);
   U500 : BUF_X1 port map( A => n154, Z => n152);
   U501 : BUF_X1 port map( A => n341, Z => n340);
   U502 : BUF_X1 port map( A => n307, Z => n306);
   U503 : BUF_X1 port map( A => n205_port, Z => n204_port);
   U504 : BUF_X1 port map( A => n171_port, Z => n170_port);
   U505 : BUF_X1 port map( A => n324, Z => n323);
   U506 : BUF_X1 port map( A => n290, Z => n289);
   U507 : BUF_X1 port map( A => n188, Z => n187_port);
   U508 : BUF_X1 port map( A => n154, Z => n153);
   U509 : BUF_X1 port map( A => n13, Z => n346);
   U510 : BUF_X1 port map( A => n12, Z => n329);
   U511 : BUF_X1 port map( A => n11, Z => n312);
   U512 : BUF_X1 port map( A => n2, Z => n295);
   U513 : BUF_X1 port map( A => n7, Z => n210_port);
   U514 : BUF_X1 port map( A => n6, Z => n193_port);
   U515 : BUF_X1 port map( A => n5, Z => n176_port);
   U516 : BUF_X1 port map( A => n1, Z => n159_port);
   U517 : BUF_X1 port map( A => n565, Z => n564);
   U518 : INV_X1 port map( A => ADD_RD2(0), ZN => n3082);
   U519 : INV_X1 port map( A => ADD_RD1(0), ZN => n1246);
   U520 : INV_X1 port map( A => ADD_RD2(2), ZN => n3084);
   U521 : INV_X1 port map( A => ADD_RD1(2), ZN => n1248);
   U522 : INV_X1 port map( A => ADD_RD2(1), ZN => n3083);
   U523 : INV_X1 port map( A => ADD_RD1(1), ZN => n1247);
   U524 : INV_X1 port map( A => ADD_RD2(3), ZN => n3085);
   U525 : INV_X1 port map( A => ADD_RD1(3), ZN => n1249);
   U526 : NOR2_X1 port map( A1 => n1248, A2 => ADD_RD1(1), ZN => n566);
   U527 : NOR2_X1 port map( A1 => n1248, A2 => n1247, ZN => n567);
   U528 : AOI22_X1 port map( A1 => REGISTERS_21_0_port, A2 => n160_port, B1 => 
                           REGISTERS_23_0_port, B2 => n143, ZN => n573);
   U529 : NOR2_X1 port map( A1 => ADD_RD1(1), A2 => ADD_RD1(2), ZN => n568);
   U530 : NOR2_X1 port map( A1 => n1247, A2 => ADD_RD1(2), ZN => n569);
   U531 : AOI22_X1 port map( A1 => REGISTERS_17_0_port, A2 => n194_port, B1 => 
                           REGISTERS_19_0_port, B2 => n177_port, ZN => n572);
   U532 : AOI22_X1 port map( A1 => REGISTERS_20_0_port, A2 => n228, B1 => 
                           REGISTERS_22_0_port, B2 => n211_port, ZN => n571);
   U533 : AOI22_X1 port map( A1 => REGISTERS_16_0_port, A2 => n262, B1 => 
                           REGISTERS_18_0_port, B2 => n245, ZN => n570);
   U534 : AND4_X1 port map( A1 => n573, A2 => n572, A3 => n571, A4 => n570, ZN 
                           => n590);
   U535 : AOI22_X1 port map( A1 => REGISTERS_29_0_port, A2 => n160_port, B1 => 
                           REGISTERS_31_0_port, B2 => n143, ZN => n577);
   U536 : AOI22_X1 port map( A1 => REGISTERS_25_0_port, A2 => n194_port, B1 => 
                           REGISTERS_27_0_port, B2 => n177_port, ZN => n576);
   U537 : AOI22_X1 port map( A1 => REGISTERS_28_0_port, A2 => n228, B1 => 
                           REGISTERS_30_0_port, B2 => n211_port, ZN => n575);
   U538 : AOI22_X1 port map( A1 => REGISTERS_24_0_port, A2 => n262, B1 => 
                           REGISTERS_26_0_port, B2 => n245, ZN => n574);
   U539 : AND4_X1 port map( A1 => n577, A2 => n576, A3 => n575, A4 => n574, ZN 
                           => n589);
   U540 : AOI22_X1 port map( A1 => REGISTERS_5_0_port, A2 => n160_port, B1 => 
                           REGISTERS_7_0_port, B2 => n143, ZN => n581);
   U541 : AOI22_X1 port map( A1 => REGISTERS_1_0_port, A2 => n194_port, B1 => 
                           REGISTERS_3_0_port, B2 => n177_port, ZN => n580);
   U542 : AOI22_X1 port map( A1 => REGISTERS_4_0_port, A2 => n228, B1 => 
                           REGISTERS_6_0_port, B2 => n211_port, ZN => n579);
   U543 : AOI22_X1 port map( A1 => REGISTERS_0_0_port, A2 => n262, B1 => 
                           REGISTERS_2_0_port, B2 => n245, ZN => n578);
   U544 : NAND4_X1 port map( A1 => n581, A2 => n580, A3 => n579, A4 => n578, ZN
                           => n587);
   U545 : AOI22_X1 port map( A1 => REGISTERS_13_0_port, A2 => n160_port, B1 => 
                           REGISTERS_15_0_port, B2 => n143, ZN => n585);
   U546 : AOI22_X1 port map( A1 => REGISTERS_9_0_port, A2 => n194_port, B1 => 
                           REGISTERS_11_0_port, B2 => n177_port, ZN => n584);
   U547 : AOI22_X1 port map( A1 => REGISTERS_12_0_port, A2 => n228, B1 => 
                           REGISTERS_14_0_port, B2 => n211_port, ZN => n583);
   U548 : AOI22_X1 port map( A1 => REGISTERS_8_0_port, A2 => n262, B1 => 
                           REGISTERS_10_0_port, B2 => n245, ZN => n582);
   U549 : NAND4_X1 port map( A1 => n585, A2 => n584, A3 => n583, A4 => n582, ZN
                           => n586);
   U550 : AOI22_X1 port map( A1 => n587, A2 => n1240, B1 => n586, B2 => n1238, 
                           ZN => n588);
   U551 : OAI221_X1 port map( B1 => n1244, B2 => n590, C1 => n1242, C2 => n589,
                           A => n588, ZN => N187);
   U552 : AOI22_X1 port map( A1 => REGISTERS_21_1_port, A2 => n160_port, B1 => 
                           REGISTERS_23_1_port, B2 => n143, ZN => n594);
   U553 : AOI22_X1 port map( A1 => REGISTERS_17_1_port, A2 => n194_port, B1 => 
                           REGISTERS_19_1_port, B2 => n177_port, ZN => n593);
   U554 : AOI22_X1 port map( A1 => REGISTERS_20_1_port, A2 => n228, B1 => 
                           REGISTERS_22_1_port, B2 => n211_port, ZN => n592);
   U555 : AOI22_X1 port map( A1 => REGISTERS_16_1_port, A2 => n262, B1 => 
                           REGISTERS_18_1_port, B2 => n245, ZN => n591);
   U556 : AND4_X1 port map( A1 => n594, A2 => n593, A3 => n592, A4 => n591, ZN 
                           => n611);
   U557 : AOI22_X1 port map( A1 => REGISTERS_29_1_port, A2 => n160_port, B1 => 
                           REGISTERS_31_1_port, B2 => n143, ZN => n598);
   U558 : AOI22_X1 port map( A1 => REGISTERS_25_1_port, A2 => n194_port, B1 => 
                           REGISTERS_27_1_port, B2 => n177_port, ZN => n597);
   U559 : AOI22_X1 port map( A1 => REGISTERS_28_1_port, A2 => n228, B1 => 
                           REGISTERS_30_1_port, B2 => n211_port, ZN => n596);
   U560 : AOI22_X1 port map( A1 => REGISTERS_24_1_port, A2 => n262, B1 => 
                           REGISTERS_26_1_port, B2 => n245, ZN => n595);
   U561 : AND4_X1 port map( A1 => n598, A2 => n597, A3 => n596, A4 => n595, ZN 
                           => n610);
   U562 : AOI22_X1 port map( A1 => REGISTERS_5_1_port, A2 => n160_port, B1 => 
                           REGISTERS_7_1_port, B2 => n143, ZN => n602);
   U563 : AOI22_X1 port map( A1 => REGISTERS_1_1_port, A2 => n194_port, B1 => 
                           REGISTERS_3_1_port, B2 => n177_port, ZN => n601);
   U564 : AOI22_X1 port map( A1 => REGISTERS_4_1_port, A2 => n228, B1 => 
                           REGISTERS_6_1_port, B2 => n211_port, ZN => n600);
   U565 : AOI22_X1 port map( A1 => REGISTERS_0_1_port, A2 => n262, B1 => 
                           REGISTERS_2_1_port, B2 => n245, ZN => n599);
   U566 : NAND4_X1 port map( A1 => n602, A2 => n601, A3 => n600, A4 => n599, ZN
                           => n608);
   U567 : AOI22_X1 port map( A1 => REGISTERS_13_1_port, A2 => n160_port, B1 => 
                           REGISTERS_15_1_port, B2 => n143, ZN => n606);
   U568 : AOI22_X1 port map( A1 => REGISTERS_9_1_port, A2 => n194_port, B1 => 
                           REGISTERS_11_1_port, B2 => n177_port, ZN => n605);
   U569 : AOI22_X1 port map( A1 => REGISTERS_12_1_port, A2 => n228, B1 => 
                           REGISTERS_14_1_port, B2 => n211_port, ZN => n604);
   U570 : AOI22_X1 port map( A1 => REGISTERS_8_1_port, A2 => n262, B1 => 
                           REGISTERS_10_1_port, B2 => n245, ZN => n603);
   U571 : NAND4_X1 port map( A1 => n606, A2 => n605, A3 => n604, A4 => n603, ZN
                           => n607);
   U572 : AOI22_X1 port map( A1 => n608, A2 => n1240, B1 => n607, B2 => n1238, 
                           ZN => n609);
   U573 : OAI221_X1 port map( B1 => n1244, B2 => n611, C1 => n1242, C2 => n610,
                           A => n609, ZN => N186);
   U574 : AOI22_X1 port map( A1 => REGISTERS_21_2_port, A2 => n160_port, B1 => 
                           REGISTERS_23_2_port, B2 => n143, ZN => n615);
   U575 : AOI22_X1 port map( A1 => REGISTERS_17_2_port, A2 => n194_port, B1 => 
                           REGISTERS_19_2_port, B2 => n177_port, ZN => n614);
   U576 : AOI22_X1 port map( A1 => REGISTERS_20_2_port, A2 => n228, B1 => 
                           REGISTERS_22_2_port, B2 => n211_port, ZN => n613);
   U577 : AOI22_X1 port map( A1 => REGISTERS_16_2_port, A2 => n262, B1 => 
                           REGISTERS_18_2_port, B2 => n245, ZN => n612);
   U578 : AND4_X1 port map( A1 => n615, A2 => n614, A3 => n613, A4 => n612, ZN 
                           => n632);
   U579 : AOI22_X1 port map( A1 => REGISTERS_29_2_port, A2 => n160_port, B1 => 
                           REGISTERS_31_2_port, B2 => n143, ZN => n619);
   U580 : AOI22_X1 port map( A1 => REGISTERS_25_2_port, A2 => n194_port, B1 => 
                           REGISTERS_27_2_port, B2 => n177_port, ZN => n618);
   U581 : AOI22_X1 port map( A1 => REGISTERS_28_2_port, A2 => n228, B1 => 
                           REGISTERS_30_2_port, B2 => n211_port, ZN => n617);
   U582 : AOI22_X1 port map( A1 => REGISTERS_24_2_port, A2 => n262, B1 => 
                           REGISTERS_26_2_port, B2 => n245, ZN => n616);
   U583 : AND4_X1 port map( A1 => n619, A2 => n618, A3 => n617, A4 => n616, ZN 
                           => n631);
   U584 : AOI22_X1 port map( A1 => REGISTERS_5_2_port, A2 => n160_port, B1 => 
                           REGISTERS_7_2_port, B2 => n143, ZN => n623);
   U585 : AOI22_X1 port map( A1 => REGISTERS_1_2_port, A2 => n194_port, B1 => 
                           REGISTERS_3_2_port, B2 => n177_port, ZN => n622);
   U586 : AOI22_X1 port map( A1 => REGISTERS_4_2_port, A2 => n228, B1 => 
                           REGISTERS_6_2_port, B2 => n211_port, ZN => n621);
   U587 : AOI22_X1 port map( A1 => REGISTERS_0_2_port, A2 => n262, B1 => 
                           REGISTERS_2_2_port, B2 => n245, ZN => n620);
   U588 : NAND4_X1 port map( A1 => n623, A2 => n622, A3 => n621, A4 => n620, ZN
                           => n629);
   U589 : AOI22_X1 port map( A1 => REGISTERS_13_2_port, A2 => n160_port, B1 => 
                           REGISTERS_15_2_port, B2 => n143, ZN => n627);
   U590 : AOI22_X1 port map( A1 => REGISTERS_9_2_port, A2 => n194_port, B1 => 
                           REGISTERS_11_2_port, B2 => n177_port, ZN => n626);
   U591 : AOI22_X1 port map( A1 => REGISTERS_12_2_port, A2 => n228, B1 => 
                           REGISTERS_14_2_port, B2 => n211_port, ZN => n625);
   U592 : AOI22_X1 port map( A1 => REGISTERS_8_2_port, A2 => n262, B1 => 
                           REGISTERS_10_2_port, B2 => n245, ZN => n624);
   U593 : NAND4_X1 port map( A1 => n627, A2 => n626, A3 => n625, A4 => n624, ZN
                           => n628);
   U594 : AOI22_X1 port map( A1 => n629, A2 => n1240, B1 => n628, B2 => n1238, 
                           ZN => n630);
   U595 : OAI221_X1 port map( B1 => n1244, B2 => n632, C1 => n1242, C2 => n631,
                           A => n630, ZN => N185);
   U596 : AOI22_X1 port map( A1 => REGISTERS_21_3_port, A2 => n161_port, B1 => 
                           REGISTERS_23_3_port, B2 => n144, ZN => n636);
   U597 : AOI22_X1 port map( A1 => REGISTERS_17_3_port, A2 => n195_port, B1 => 
                           REGISTERS_19_3_port, B2 => n178_port, ZN => n635);
   U598 : AOI22_X1 port map( A1 => REGISTERS_20_3_port, A2 => n229, B1 => 
                           REGISTERS_22_3_port, B2 => n212_port, ZN => n634);
   U599 : AOI22_X1 port map( A1 => REGISTERS_16_3_port, A2 => n263, B1 => 
                           REGISTERS_18_3_port, B2 => n246, ZN => n633);
   U600 : AND4_X1 port map( A1 => n636, A2 => n635, A3 => n634, A4 => n633, ZN 
                           => n653);
   U601 : AOI22_X1 port map( A1 => REGISTERS_29_3_port, A2 => n161_port, B1 => 
                           REGISTERS_31_3_port, B2 => n144, ZN => n640);
   U602 : AOI22_X1 port map( A1 => REGISTERS_25_3_port, A2 => n195_port, B1 => 
                           REGISTERS_27_3_port, B2 => n178_port, ZN => n639);
   U603 : AOI22_X1 port map( A1 => REGISTERS_28_3_port, A2 => n229, B1 => 
                           REGISTERS_30_3_port, B2 => n212_port, ZN => n638);
   U604 : AOI22_X1 port map( A1 => REGISTERS_24_3_port, A2 => n263, B1 => 
                           REGISTERS_26_3_port, B2 => n246, ZN => n637);
   U605 : AND4_X1 port map( A1 => n640, A2 => n639, A3 => n638, A4 => n637, ZN 
                           => n652);
   U606 : AOI22_X1 port map( A1 => REGISTERS_5_3_port, A2 => n161_port, B1 => 
                           REGISTERS_7_3_port, B2 => n144, ZN => n644);
   U607 : AOI22_X1 port map( A1 => REGISTERS_1_3_port, A2 => n195_port, B1 => 
                           REGISTERS_3_3_port, B2 => n178_port, ZN => n643);
   U608 : AOI22_X1 port map( A1 => REGISTERS_4_3_port, A2 => n229, B1 => 
                           REGISTERS_6_3_port, B2 => n212_port, ZN => n642);
   U609 : AOI22_X1 port map( A1 => REGISTERS_0_3_port, A2 => n263, B1 => 
                           REGISTERS_2_3_port, B2 => n246, ZN => n641);
   U610 : NAND4_X1 port map( A1 => n644, A2 => n643, A3 => n642, A4 => n641, ZN
                           => n650);
   U611 : AOI22_X1 port map( A1 => REGISTERS_13_3_port, A2 => n161_port, B1 => 
                           REGISTERS_15_3_port, B2 => n144, ZN => n648);
   U612 : AOI22_X1 port map( A1 => REGISTERS_9_3_port, A2 => n195_port, B1 => 
                           REGISTERS_11_3_port, B2 => n178_port, ZN => n647);
   U613 : AOI22_X1 port map( A1 => REGISTERS_12_3_port, A2 => n229, B1 => 
                           REGISTERS_14_3_port, B2 => n212_port, ZN => n646);
   U614 : AOI22_X1 port map( A1 => REGISTERS_8_3_port, A2 => n263, B1 => 
                           REGISTERS_10_3_port, B2 => n246, ZN => n645);
   U615 : NAND4_X1 port map( A1 => n648, A2 => n647, A3 => n646, A4 => n645, ZN
                           => n649);
   U616 : AOI22_X1 port map( A1 => n650, A2 => n1240, B1 => n649, B2 => n1238, 
                           ZN => n651);
   U617 : OAI221_X1 port map( B1 => n1244, B2 => n653, C1 => n1242, C2 => n652,
                           A => n651, ZN => N184);
   U618 : AOI22_X1 port map( A1 => REGISTERS_21_4_port, A2 => n161_port, B1 => 
                           REGISTERS_23_4_port, B2 => n144, ZN => n657);
   U619 : AOI22_X1 port map( A1 => REGISTERS_17_4_port, A2 => n195_port, B1 => 
                           REGISTERS_19_4_port, B2 => n178_port, ZN => n656);
   U620 : AOI22_X1 port map( A1 => REGISTERS_20_4_port, A2 => n229, B1 => 
                           REGISTERS_22_4_port, B2 => n212_port, ZN => n655);
   U621 : AOI22_X1 port map( A1 => REGISTERS_16_4_port, A2 => n263, B1 => 
                           REGISTERS_18_4_port, B2 => n246, ZN => n654);
   U622 : AND4_X1 port map( A1 => n657, A2 => n656, A3 => n655, A4 => n654, ZN 
                           => n674);
   U623 : AOI22_X1 port map( A1 => REGISTERS_29_4_port, A2 => n161_port, B1 => 
                           REGISTERS_31_4_port, B2 => n144, ZN => n661);
   U624 : AOI22_X1 port map( A1 => REGISTERS_25_4_port, A2 => n195_port, B1 => 
                           REGISTERS_27_4_port, B2 => n178_port, ZN => n660);
   U625 : AOI22_X1 port map( A1 => REGISTERS_28_4_port, A2 => n229, B1 => 
                           REGISTERS_30_4_port, B2 => n212_port, ZN => n659);
   U626 : AOI22_X1 port map( A1 => REGISTERS_24_4_port, A2 => n263, B1 => 
                           REGISTERS_26_4_port, B2 => n246, ZN => n658);
   U627 : AND4_X1 port map( A1 => n661, A2 => n660, A3 => n659, A4 => n658, ZN 
                           => n673);
   U628 : AOI22_X1 port map( A1 => REGISTERS_5_4_port, A2 => n161_port, B1 => 
                           REGISTERS_7_4_port, B2 => n144, ZN => n665);
   U629 : AOI22_X1 port map( A1 => REGISTERS_1_4_port, A2 => n195_port, B1 => 
                           REGISTERS_3_4_port, B2 => n178_port, ZN => n664);
   U630 : AOI22_X1 port map( A1 => REGISTERS_4_4_port, A2 => n229, B1 => 
                           REGISTERS_6_4_port, B2 => n212_port, ZN => n663);
   U631 : AOI22_X1 port map( A1 => REGISTERS_0_4_port, A2 => n263, B1 => 
                           REGISTERS_2_4_port, B2 => n246, ZN => n662);
   U632 : NAND4_X1 port map( A1 => n665, A2 => n664, A3 => n663, A4 => n662, ZN
                           => n671);
   U633 : AOI22_X1 port map( A1 => REGISTERS_13_4_port, A2 => n161_port, B1 => 
                           REGISTERS_15_4_port, B2 => n144, ZN => n669);
   U634 : AOI22_X1 port map( A1 => REGISTERS_9_4_port, A2 => n195_port, B1 => 
                           REGISTERS_11_4_port, B2 => n178_port, ZN => n668);
   U635 : AOI22_X1 port map( A1 => REGISTERS_12_4_port, A2 => n229, B1 => 
                           REGISTERS_14_4_port, B2 => n212_port, ZN => n667);
   U636 : AOI22_X1 port map( A1 => REGISTERS_8_4_port, A2 => n263, B1 => 
                           REGISTERS_10_4_port, B2 => n246, ZN => n666);
   U637 : NAND4_X1 port map( A1 => n669, A2 => n668, A3 => n667, A4 => n666, ZN
                           => n670);
   U638 : AOI22_X1 port map( A1 => n671, A2 => n1240, B1 => n670, B2 => n1238, 
                           ZN => n672);
   U639 : OAI221_X1 port map( B1 => n1244, B2 => n674, C1 => n1242, C2 => n673,
                           A => n672, ZN => N183);
   U640 : AOI22_X1 port map( A1 => REGISTERS_21_5_port, A2 => n161_port, B1 => 
                           REGISTERS_23_5_port, B2 => n144, ZN => n678);
   U641 : AOI22_X1 port map( A1 => REGISTERS_17_5_port, A2 => n195_port, B1 => 
                           REGISTERS_19_5_port, B2 => n178_port, ZN => n677);
   U642 : AOI22_X1 port map( A1 => REGISTERS_20_5_port, A2 => n229, B1 => 
                           REGISTERS_22_5_port, B2 => n212_port, ZN => n676);
   U643 : AOI22_X1 port map( A1 => REGISTERS_16_5_port, A2 => n263, B1 => 
                           REGISTERS_18_5_port, B2 => n246, ZN => n675);
   U644 : AND4_X1 port map( A1 => n678, A2 => n677, A3 => n676, A4 => n675, ZN 
                           => n695);
   U645 : AOI22_X1 port map( A1 => REGISTERS_29_5_port, A2 => n161_port, B1 => 
                           REGISTERS_31_5_port, B2 => n144, ZN => n682);
   U646 : AOI22_X1 port map( A1 => REGISTERS_25_5_port, A2 => n195_port, B1 => 
                           REGISTERS_27_5_port, B2 => n178_port, ZN => n681);
   U647 : AOI22_X1 port map( A1 => REGISTERS_28_5_port, A2 => n229, B1 => 
                           REGISTERS_30_5_port, B2 => n212_port, ZN => n680);
   U648 : AOI22_X1 port map( A1 => REGISTERS_24_5_port, A2 => n263, B1 => 
                           REGISTERS_26_5_port, B2 => n246, ZN => n679);
   U649 : AND4_X1 port map( A1 => n682, A2 => n681, A3 => n680, A4 => n679, ZN 
                           => n694);
   U650 : AOI22_X1 port map( A1 => REGISTERS_5_5_port, A2 => n161_port, B1 => 
                           REGISTERS_7_5_port, B2 => n144, ZN => n686);
   U651 : AOI22_X1 port map( A1 => REGISTERS_1_5_port, A2 => n195_port, B1 => 
                           REGISTERS_3_5_port, B2 => n178_port, ZN => n685);
   U652 : AOI22_X1 port map( A1 => REGISTERS_4_5_port, A2 => n229, B1 => 
                           REGISTERS_6_5_port, B2 => n212_port, ZN => n684);
   U653 : AOI22_X1 port map( A1 => REGISTERS_0_5_port, A2 => n263, B1 => 
                           REGISTERS_2_5_port, B2 => n246, ZN => n683);
   U654 : NAND4_X1 port map( A1 => n686, A2 => n685, A3 => n684, A4 => n683, ZN
                           => n692);
   U655 : AOI22_X1 port map( A1 => REGISTERS_13_5_port, A2 => n161_port, B1 => 
                           REGISTERS_15_5_port, B2 => n144, ZN => n690);
   U656 : AOI22_X1 port map( A1 => REGISTERS_9_5_port, A2 => n195_port, B1 => 
                           REGISTERS_11_5_port, B2 => n178_port, ZN => n689);
   U657 : AOI22_X1 port map( A1 => REGISTERS_12_5_port, A2 => n229, B1 => 
                           REGISTERS_14_5_port, B2 => n212_port, ZN => n688);
   U658 : AOI22_X1 port map( A1 => REGISTERS_8_5_port, A2 => n263, B1 => 
                           REGISTERS_10_5_port, B2 => n246, ZN => n687);
   U659 : NAND4_X1 port map( A1 => n690, A2 => n689, A3 => n688, A4 => n687, ZN
                           => n691);
   U660 : AOI22_X1 port map( A1 => n692, A2 => n1240, B1 => n691, B2 => n1238, 
                           ZN => n693);
   U661 : OAI221_X1 port map( B1 => n1244, B2 => n695, C1 => n1242, C2 => n694,
                           A => n693, ZN => N182);
   U662 : AOI22_X1 port map( A1 => REGISTERS_21_6_port, A2 => n162_port, B1 => 
                           REGISTERS_23_6_port, B2 => n145, ZN => n699);
   U663 : AOI22_X1 port map( A1 => REGISTERS_17_6_port, A2 => n196_port, B1 => 
                           REGISTERS_19_6_port, B2 => n179_port, ZN => n698);
   U664 : AOI22_X1 port map( A1 => REGISTERS_20_6_port, A2 => n230, B1 => 
                           REGISTERS_22_6_port, B2 => n213_port, ZN => n697);
   U665 : AOI22_X1 port map( A1 => REGISTERS_16_6_port, A2 => n264, B1 => 
                           REGISTERS_18_6_port, B2 => n247, ZN => n696);
   U666 : AND4_X1 port map( A1 => n699, A2 => n698, A3 => n697, A4 => n696, ZN 
                           => n716);
   U667 : AOI22_X1 port map( A1 => REGISTERS_29_6_port, A2 => n162_port, B1 => 
                           REGISTERS_31_6_port, B2 => n145, ZN => n703);
   U668 : AOI22_X1 port map( A1 => REGISTERS_25_6_port, A2 => n196_port, B1 => 
                           REGISTERS_27_6_port, B2 => n179_port, ZN => n702);
   U669 : AOI22_X1 port map( A1 => REGISTERS_28_6_port, A2 => n230, B1 => 
                           REGISTERS_30_6_port, B2 => n213_port, ZN => n701);
   U670 : AOI22_X1 port map( A1 => REGISTERS_24_6_port, A2 => n264, B1 => 
                           REGISTERS_26_6_port, B2 => n247, ZN => n700);
   U671 : AND4_X1 port map( A1 => n703, A2 => n702, A3 => n701, A4 => n700, ZN 
                           => n715);
   U672 : AOI22_X1 port map( A1 => REGISTERS_5_6_port, A2 => n162_port, B1 => 
                           REGISTERS_7_6_port, B2 => n145, ZN => n707);
   U673 : AOI22_X1 port map( A1 => REGISTERS_1_6_port, A2 => n196_port, B1 => 
                           REGISTERS_3_6_port, B2 => n179_port, ZN => n706);
   U674 : AOI22_X1 port map( A1 => REGISTERS_4_6_port, A2 => n230, B1 => 
                           REGISTERS_6_6_port, B2 => n213_port, ZN => n705);
   U675 : AOI22_X1 port map( A1 => REGISTERS_0_6_port, A2 => n264, B1 => 
                           REGISTERS_2_6_port, B2 => n247, ZN => n704);
   U676 : NAND4_X1 port map( A1 => n707, A2 => n706, A3 => n705, A4 => n704, ZN
                           => n713);
   U677 : AOI22_X1 port map( A1 => REGISTERS_13_6_port, A2 => n162_port, B1 => 
                           REGISTERS_15_6_port, B2 => n145, ZN => n711);
   U678 : AOI22_X1 port map( A1 => REGISTERS_9_6_port, A2 => n196_port, B1 => 
                           REGISTERS_11_6_port, B2 => n179_port, ZN => n710);
   U679 : AOI22_X1 port map( A1 => REGISTERS_12_6_port, A2 => n230, B1 => 
                           REGISTERS_14_6_port, B2 => n213_port, ZN => n709);
   U680 : AOI22_X1 port map( A1 => REGISTERS_8_6_port, A2 => n264, B1 => 
                           REGISTERS_10_6_port, B2 => n247, ZN => n708);
   U681 : NAND4_X1 port map( A1 => n711, A2 => n710, A3 => n709, A4 => n708, ZN
                           => n712);
   U682 : AOI22_X1 port map( A1 => n713, A2 => n1240, B1 => n712, B2 => n1238, 
                           ZN => n714);
   U683 : OAI221_X1 port map( B1 => n1244, B2 => n716, C1 => n1242, C2 => n715,
                           A => n714, ZN => N181);
   U684 : AOI22_X1 port map( A1 => REGISTERS_21_7_port, A2 => n162_port, B1 => 
                           REGISTERS_23_7_port, B2 => n145, ZN => n720);
   U685 : AOI22_X1 port map( A1 => REGISTERS_17_7_port, A2 => n196_port, B1 => 
                           REGISTERS_19_7_port, B2 => n179_port, ZN => n719);
   U686 : AOI22_X1 port map( A1 => REGISTERS_20_7_port, A2 => n230, B1 => 
                           REGISTERS_22_7_port, B2 => n213_port, ZN => n718);
   U687 : AOI22_X1 port map( A1 => REGISTERS_16_7_port, A2 => n264, B1 => 
                           REGISTERS_18_7_port, B2 => n247, ZN => n717);
   U688 : AND4_X1 port map( A1 => n720, A2 => n719, A3 => n718, A4 => n717, ZN 
                           => n737);
   U689 : AOI22_X1 port map( A1 => REGISTERS_29_7_port, A2 => n162_port, B1 => 
                           REGISTERS_31_7_port, B2 => n145, ZN => n724);
   U690 : AOI22_X1 port map( A1 => REGISTERS_25_7_port, A2 => n196_port, B1 => 
                           REGISTERS_27_7_port, B2 => n179_port, ZN => n723);
   U691 : AOI22_X1 port map( A1 => REGISTERS_28_7_port, A2 => n230, B1 => 
                           REGISTERS_30_7_port, B2 => n213_port, ZN => n722);
   U692 : AOI22_X1 port map( A1 => REGISTERS_24_7_port, A2 => n264, B1 => 
                           REGISTERS_26_7_port, B2 => n247, ZN => n721);
   U693 : AND4_X1 port map( A1 => n724, A2 => n723, A3 => n722, A4 => n721, ZN 
                           => n736);
   U694 : AOI22_X1 port map( A1 => REGISTERS_5_7_port, A2 => n162_port, B1 => 
                           REGISTERS_7_7_port, B2 => n145, ZN => n728);
   U695 : AOI22_X1 port map( A1 => REGISTERS_1_7_port, A2 => n196_port, B1 => 
                           REGISTERS_3_7_port, B2 => n179_port, ZN => n727);
   U696 : AOI22_X1 port map( A1 => REGISTERS_4_7_port, A2 => n230, B1 => 
                           REGISTERS_6_7_port, B2 => n213_port, ZN => n726);
   U697 : AOI22_X1 port map( A1 => REGISTERS_0_7_port, A2 => n264, B1 => 
                           REGISTERS_2_7_port, B2 => n247, ZN => n725);
   U698 : NAND4_X1 port map( A1 => n728, A2 => n727, A3 => n726, A4 => n725, ZN
                           => n734);
   U699 : AOI22_X1 port map( A1 => REGISTERS_13_7_port, A2 => n162_port, B1 => 
                           REGISTERS_15_7_port, B2 => n145, ZN => n732);
   U700 : AOI22_X1 port map( A1 => REGISTERS_9_7_port, A2 => n196_port, B1 => 
                           REGISTERS_11_7_port, B2 => n179_port, ZN => n731);
   U701 : AOI22_X1 port map( A1 => REGISTERS_12_7_port, A2 => n230, B1 => 
                           REGISTERS_14_7_port, B2 => n213_port, ZN => n730);
   U702 : AOI22_X1 port map( A1 => REGISTERS_8_7_port, A2 => n264, B1 => 
                           REGISTERS_10_7_port, B2 => n247, ZN => n729);
   U703 : NAND4_X1 port map( A1 => n732, A2 => n731, A3 => n730, A4 => n729, ZN
                           => n733);
   U704 : AOI22_X1 port map( A1 => n734, A2 => n1240, B1 => n733, B2 => n1238, 
                           ZN => n735);
   U705 : OAI221_X1 port map( B1 => n1244, B2 => n737, C1 => n1242, C2 => n736,
                           A => n735, ZN => N180);
   U706 : AOI22_X1 port map( A1 => REGISTERS_21_8_port, A2 => n162_port, B1 => 
                           REGISTERS_23_8_port, B2 => n145, ZN => n741);
   U707 : AOI22_X1 port map( A1 => REGISTERS_17_8_port, A2 => n196_port, B1 => 
                           REGISTERS_19_8_port, B2 => n179_port, ZN => n740);
   U708 : AOI22_X1 port map( A1 => REGISTERS_20_8_port, A2 => n230, B1 => 
                           REGISTERS_22_8_port, B2 => n213_port, ZN => n739);
   U709 : AOI22_X1 port map( A1 => REGISTERS_16_8_port, A2 => n264, B1 => 
                           REGISTERS_18_8_port, B2 => n247, ZN => n738);
   U710 : AND4_X1 port map( A1 => n741, A2 => n740, A3 => n739, A4 => n738, ZN 
                           => n758);
   U711 : AOI22_X1 port map( A1 => REGISTERS_29_8_port, A2 => n162_port, B1 => 
                           REGISTERS_31_8_port, B2 => n145, ZN => n745);
   U712 : AOI22_X1 port map( A1 => REGISTERS_25_8_port, A2 => n196_port, B1 => 
                           REGISTERS_27_8_port, B2 => n179_port, ZN => n744);
   U713 : AOI22_X1 port map( A1 => REGISTERS_28_8_port, A2 => n230, B1 => 
                           REGISTERS_30_8_port, B2 => n213_port, ZN => n743);
   U714 : AOI22_X1 port map( A1 => REGISTERS_24_8_port, A2 => n264, B1 => 
                           REGISTERS_26_8_port, B2 => n247, ZN => n742);
   U715 : AND4_X1 port map( A1 => n745, A2 => n744, A3 => n743, A4 => n742, ZN 
                           => n757);
   U716 : AOI22_X1 port map( A1 => REGISTERS_5_8_port, A2 => n162_port, B1 => 
                           REGISTERS_7_8_port, B2 => n145, ZN => n749);
   U717 : AOI22_X1 port map( A1 => REGISTERS_1_8_port, A2 => n196_port, B1 => 
                           REGISTERS_3_8_port, B2 => n179_port, ZN => n748);
   U718 : AOI22_X1 port map( A1 => REGISTERS_4_8_port, A2 => n230, B1 => 
                           REGISTERS_6_8_port, B2 => n213_port, ZN => n747);
   U719 : AOI22_X1 port map( A1 => REGISTERS_0_8_port, A2 => n264, B1 => 
                           REGISTERS_2_8_port, B2 => n247, ZN => n746);
   U720 : NAND4_X1 port map( A1 => n749, A2 => n748, A3 => n747, A4 => n746, ZN
                           => n755);
   U721 : AOI22_X1 port map( A1 => REGISTERS_13_8_port, A2 => n162_port, B1 => 
                           REGISTERS_15_8_port, B2 => n145, ZN => n753);
   U722 : AOI22_X1 port map( A1 => REGISTERS_9_8_port, A2 => n196_port, B1 => 
                           REGISTERS_11_8_port, B2 => n179_port, ZN => n752);
   U723 : AOI22_X1 port map( A1 => REGISTERS_12_8_port, A2 => n230, B1 => 
                           REGISTERS_14_8_port, B2 => n213_port, ZN => n751);
   U724 : AOI22_X1 port map( A1 => REGISTERS_8_8_port, A2 => n264, B1 => 
                           REGISTERS_10_8_port, B2 => n247, ZN => n750);
   U725 : NAND4_X1 port map( A1 => n753, A2 => n752, A3 => n751, A4 => n750, ZN
                           => n754);
   U726 : AOI22_X1 port map( A1 => n755, A2 => n1240, B1 => n754, B2 => n1238, 
                           ZN => n756);
   U727 : OAI221_X1 port map( B1 => n1244, B2 => n758, C1 => n1242, C2 => n757,
                           A => n756, ZN => N179);
   U728 : AOI22_X1 port map( A1 => REGISTERS_21_9_port, A2 => n163_port, B1 => 
                           REGISTERS_23_9_port, B2 => n146, ZN => n762);
   U729 : AOI22_X1 port map( A1 => REGISTERS_17_9_port, A2 => n197_port, B1 => 
                           REGISTERS_19_9_port, B2 => n180_port, ZN => n761);
   U730 : AOI22_X1 port map( A1 => REGISTERS_20_9_port, A2 => n231, B1 => 
                           REGISTERS_22_9_port, B2 => n214_port, ZN => n760);
   U731 : AOI22_X1 port map( A1 => REGISTERS_16_9_port, A2 => n265, B1 => 
                           REGISTERS_18_9_port, B2 => n248, ZN => n759);
   U732 : AND4_X1 port map( A1 => n762, A2 => n761, A3 => n760, A4 => n759, ZN 
                           => n779);
   U733 : AOI22_X1 port map( A1 => REGISTERS_29_9_port, A2 => n163_port, B1 => 
                           REGISTERS_31_9_port, B2 => n146, ZN => n766);
   U734 : AOI22_X1 port map( A1 => REGISTERS_25_9_port, A2 => n197_port, B1 => 
                           REGISTERS_27_9_port, B2 => n180_port, ZN => n765);
   U735 : AOI22_X1 port map( A1 => REGISTERS_28_9_port, A2 => n231, B1 => 
                           REGISTERS_30_9_port, B2 => n214_port, ZN => n764);
   U736 : AOI22_X1 port map( A1 => REGISTERS_24_9_port, A2 => n265, B1 => 
                           REGISTERS_26_9_port, B2 => n248, ZN => n763);
   U737 : AND4_X1 port map( A1 => n766, A2 => n765, A3 => n764, A4 => n763, ZN 
                           => n778);
   U738 : AOI22_X1 port map( A1 => REGISTERS_5_9_port, A2 => n163_port, B1 => 
                           REGISTERS_7_9_port, B2 => n146, ZN => n770);
   U739 : AOI22_X1 port map( A1 => REGISTERS_1_9_port, A2 => n197_port, B1 => 
                           REGISTERS_3_9_port, B2 => n180_port, ZN => n769);
   U740 : AOI22_X1 port map( A1 => REGISTERS_4_9_port, A2 => n231, B1 => 
                           REGISTERS_6_9_port, B2 => n214_port, ZN => n768);
   U741 : AOI22_X1 port map( A1 => REGISTERS_0_9_port, A2 => n265, B1 => 
                           REGISTERS_2_9_port, B2 => n248, ZN => n767);
   U742 : NAND4_X1 port map( A1 => n770, A2 => n769, A3 => n768, A4 => n767, ZN
                           => n776);
   U743 : AOI22_X1 port map( A1 => REGISTERS_13_9_port, A2 => n163_port, B1 => 
                           REGISTERS_15_9_port, B2 => n146, ZN => n774);
   U744 : AOI22_X1 port map( A1 => REGISTERS_9_9_port, A2 => n197_port, B1 => 
                           REGISTERS_11_9_port, B2 => n180_port, ZN => n773);
   U745 : AOI22_X1 port map( A1 => REGISTERS_12_9_port, A2 => n231, B1 => 
                           REGISTERS_14_9_port, B2 => n214_port, ZN => n772);
   U746 : AOI22_X1 port map( A1 => REGISTERS_8_9_port, A2 => n265, B1 => 
                           REGISTERS_10_9_port, B2 => n248, ZN => n771);
   U747 : NAND4_X1 port map( A1 => n774, A2 => n773, A3 => n772, A4 => n771, ZN
                           => n775);
   U748 : AOI22_X1 port map( A1 => n776, A2 => n1240, B1 => n775, B2 => n1238, 
                           ZN => n777);
   U749 : OAI221_X1 port map( B1 => n1244, B2 => n779, C1 => n1242, C2 => n778,
                           A => n777, ZN => N178);
   U750 : AOI22_X1 port map( A1 => REGISTERS_21_10_port, A2 => n163_port, B1 =>
                           REGISTERS_23_10_port, B2 => n146, ZN => n783);
   U751 : AOI22_X1 port map( A1 => REGISTERS_17_10_port, A2 => n197_port, B1 =>
                           REGISTERS_19_10_port, B2 => n180_port, ZN => n782);
   U752 : AOI22_X1 port map( A1 => REGISTERS_20_10_port, A2 => n231, B1 => 
                           REGISTERS_22_10_port, B2 => n214_port, ZN => n781);
   U753 : AOI22_X1 port map( A1 => REGISTERS_16_10_port, A2 => n265, B1 => 
                           REGISTERS_18_10_port, B2 => n248, ZN => n780);
   U754 : AND4_X1 port map( A1 => n783, A2 => n782, A3 => n781, A4 => n780, ZN 
                           => n800);
   U755 : AOI22_X1 port map( A1 => REGISTERS_29_10_port, A2 => n163_port, B1 =>
                           REGISTERS_31_10_port, B2 => n146, ZN => n787);
   U756 : AOI22_X1 port map( A1 => REGISTERS_25_10_port, A2 => n197_port, B1 =>
                           REGISTERS_27_10_port, B2 => n180_port, ZN => n786);
   U757 : AOI22_X1 port map( A1 => REGISTERS_28_10_port, A2 => n231, B1 => 
                           REGISTERS_30_10_port, B2 => n214_port, ZN => n785);
   U758 : AOI22_X1 port map( A1 => REGISTERS_24_10_port, A2 => n265, B1 => 
                           REGISTERS_26_10_port, B2 => n248, ZN => n784);
   U759 : AND4_X1 port map( A1 => n787, A2 => n786, A3 => n785, A4 => n784, ZN 
                           => n799);
   U760 : AOI22_X1 port map( A1 => REGISTERS_5_10_port, A2 => n163_port, B1 => 
                           REGISTERS_7_10_port, B2 => n146, ZN => n791);
   U761 : AOI22_X1 port map( A1 => REGISTERS_1_10_port, A2 => n197_port, B1 => 
                           REGISTERS_3_10_port, B2 => n180_port, ZN => n790);
   U762 : AOI22_X1 port map( A1 => REGISTERS_4_10_port, A2 => n231, B1 => 
                           REGISTERS_6_10_port, B2 => n214_port, ZN => n789);
   U763 : AOI22_X1 port map( A1 => REGISTERS_0_10_port, A2 => n265, B1 => 
                           REGISTERS_2_10_port, B2 => n248, ZN => n788);
   U764 : NAND4_X1 port map( A1 => n791, A2 => n790, A3 => n789, A4 => n788, ZN
                           => n797);
   U765 : AOI22_X1 port map( A1 => REGISTERS_13_10_port, A2 => n163_port, B1 =>
                           REGISTERS_15_10_port, B2 => n146, ZN => n795);
   U766 : AOI22_X1 port map( A1 => REGISTERS_9_10_port, A2 => n197_port, B1 => 
                           REGISTERS_11_10_port, B2 => n180_port, ZN => n794);
   U767 : AOI22_X1 port map( A1 => REGISTERS_12_10_port, A2 => n231, B1 => 
                           REGISTERS_14_10_port, B2 => n214_port, ZN => n793);
   U768 : AOI22_X1 port map( A1 => REGISTERS_8_10_port, A2 => n265, B1 => 
                           REGISTERS_10_10_port, B2 => n248, ZN => n792);
   U769 : NAND4_X1 port map( A1 => n795, A2 => n794, A3 => n793, A4 => n792, ZN
                           => n796);
   U770 : AOI22_X1 port map( A1 => n797, A2 => n1240, B1 => n796, B2 => n1238, 
                           ZN => n798);
   U771 : OAI221_X1 port map( B1 => n1244, B2 => n800, C1 => n1242, C2 => n799,
                           A => n798, ZN => N177);
   U772 : AOI22_X1 port map( A1 => REGISTERS_21_11_port, A2 => n163_port, B1 =>
                           REGISTERS_23_11_port, B2 => n146, ZN => n804);
   U773 : AOI22_X1 port map( A1 => REGISTERS_17_11_port, A2 => n197_port, B1 =>
                           REGISTERS_19_11_port, B2 => n180_port, ZN => n803);
   U774 : AOI22_X1 port map( A1 => REGISTERS_20_11_port, A2 => n231, B1 => 
                           REGISTERS_22_11_port, B2 => n214_port, ZN => n802);
   U775 : AOI22_X1 port map( A1 => REGISTERS_16_11_port, A2 => n265, B1 => 
                           REGISTERS_18_11_port, B2 => n248, ZN => n801);
   U776 : AND4_X1 port map( A1 => n804, A2 => n803, A3 => n802, A4 => n801, ZN 
                           => n821);
   U777 : AOI22_X1 port map( A1 => REGISTERS_29_11_port, A2 => n163_port, B1 =>
                           REGISTERS_31_11_port, B2 => n146, ZN => n808);
   U778 : AOI22_X1 port map( A1 => REGISTERS_25_11_port, A2 => n197_port, B1 =>
                           REGISTERS_27_11_port, B2 => n180_port, ZN => n807);
   U779 : AOI22_X1 port map( A1 => REGISTERS_28_11_port, A2 => n231, B1 => 
                           REGISTERS_30_11_port, B2 => n214_port, ZN => n806);
   U780 : AOI22_X1 port map( A1 => REGISTERS_24_11_port, A2 => n265, B1 => 
                           REGISTERS_26_11_port, B2 => n248, ZN => n805);
   U781 : AND4_X1 port map( A1 => n808, A2 => n807, A3 => n806, A4 => n805, ZN 
                           => n820);
   U782 : AOI22_X1 port map( A1 => REGISTERS_5_11_port, A2 => n163_port, B1 => 
                           REGISTERS_7_11_port, B2 => n146, ZN => n812);
   U783 : AOI22_X1 port map( A1 => REGISTERS_1_11_port, A2 => n197_port, B1 => 
                           REGISTERS_3_11_port, B2 => n180_port, ZN => n811);
   U784 : AOI22_X1 port map( A1 => REGISTERS_4_11_port, A2 => n231, B1 => 
                           REGISTERS_6_11_port, B2 => n214_port, ZN => n810);
   U785 : AOI22_X1 port map( A1 => REGISTERS_0_11_port, A2 => n265, B1 => 
                           REGISTERS_2_11_port, B2 => n248, ZN => n809);
   U786 : NAND4_X1 port map( A1 => n812, A2 => n811, A3 => n810, A4 => n809, ZN
                           => n818);
   U787 : AOI22_X1 port map( A1 => REGISTERS_13_11_port, A2 => n163_port, B1 =>
                           REGISTERS_15_11_port, B2 => n146, ZN => n816);
   U788 : AOI22_X1 port map( A1 => REGISTERS_9_11_port, A2 => n197_port, B1 => 
                           REGISTERS_11_11_port, B2 => n180_port, ZN => n815);
   U789 : AOI22_X1 port map( A1 => REGISTERS_12_11_port, A2 => n231, B1 => 
                           REGISTERS_14_11_port, B2 => n214_port, ZN => n814);
   U790 : AOI22_X1 port map( A1 => REGISTERS_8_11_port, A2 => n265, B1 => 
                           REGISTERS_10_11_port, B2 => n248, ZN => n813);
   U791 : NAND4_X1 port map( A1 => n816, A2 => n815, A3 => n814, A4 => n813, ZN
                           => n817);
   U792 : AOI22_X1 port map( A1 => n818, A2 => n1240, B1 => n817, B2 => n1238, 
                           ZN => n819);
   U793 : OAI221_X1 port map( B1 => n1244, B2 => n821, C1 => n1242, C2 => n820,
                           A => n819, ZN => N176);
   U794 : AOI22_X1 port map( A1 => REGISTERS_21_12_port, A2 => n164_port, B1 =>
                           REGISTERS_23_12_port, B2 => n147, ZN => n825);
   U795 : AOI22_X1 port map( A1 => REGISTERS_17_12_port, A2 => n198_port, B1 =>
                           REGISTERS_19_12_port, B2 => n181_port, ZN => n824);
   U796 : AOI22_X1 port map( A1 => REGISTERS_20_12_port, A2 => n232, B1 => 
                           REGISTERS_22_12_port, B2 => n215_port, ZN => n823);
   U797 : AOI22_X1 port map( A1 => REGISTERS_16_12_port, A2 => n266, B1 => 
                           REGISTERS_18_12_port, B2 => n249, ZN => n822);
   U798 : AND4_X1 port map( A1 => n825, A2 => n824, A3 => n823, A4 => n822, ZN 
                           => n842);
   U799 : AOI22_X1 port map( A1 => REGISTERS_29_12_port, A2 => n164_port, B1 =>
                           REGISTERS_31_12_port, B2 => n147, ZN => n829);
   U800 : AOI22_X1 port map( A1 => REGISTERS_25_12_port, A2 => n198_port, B1 =>
                           REGISTERS_27_12_port, B2 => n181_port, ZN => n828);
   U801 : AOI22_X1 port map( A1 => REGISTERS_28_12_port, A2 => n232, B1 => 
                           REGISTERS_30_12_port, B2 => n215_port, ZN => n827);
   U802 : AOI22_X1 port map( A1 => REGISTERS_24_12_port, A2 => n266, B1 => 
                           REGISTERS_26_12_port, B2 => n249, ZN => n826);
   U803 : AND4_X1 port map( A1 => n829, A2 => n828, A3 => n827, A4 => n826, ZN 
                           => n841);
   U804 : AOI22_X1 port map( A1 => REGISTERS_5_12_port, A2 => n164_port, B1 => 
                           REGISTERS_7_12_port, B2 => n147, ZN => n833);
   U805 : AOI22_X1 port map( A1 => REGISTERS_1_12_port, A2 => n198_port, B1 => 
                           REGISTERS_3_12_port, B2 => n181_port, ZN => n832);
   U806 : AOI22_X1 port map( A1 => REGISTERS_4_12_port, A2 => n232, B1 => 
                           REGISTERS_6_12_port, B2 => n215_port, ZN => n831);
   U807 : AOI22_X1 port map( A1 => REGISTERS_0_12_port, A2 => n266, B1 => 
                           REGISTERS_2_12_port, B2 => n249, ZN => n830);
   U808 : NAND4_X1 port map( A1 => n833, A2 => n832, A3 => n831, A4 => n830, ZN
                           => n839);
   U809 : AOI22_X1 port map( A1 => REGISTERS_13_12_port, A2 => n164_port, B1 =>
                           REGISTERS_15_12_port, B2 => n147, ZN => n837);
   U810 : AOI22_X1 port map( A1 => REGISTERS_9_12_port, A2 => n198_port, B1 => 
                           REGISTERS_11_12_port, B2 => n181_port, ZN => n836);
   U811 : AOI22_X1 port map( A1 => REGISTERS_12_12_port, A2 => n232, B1 => 
                           REGISTERS_14_12_port, B2 => n215_port, ZN => n835);
   U812 : AOI22_X1 port map( A1 => REGISTERS_8_12_port, A2 => n266, B1 => 
                           REGISTERS_10_12_port, B2 => n249, ZN => n834);
   U813 : NAND4_X1 port map( A1 => n837, A2 => n836, A3 => n835, A4 => n834, ZN
                           => n838);
   U814 : AOI22_X1 port map( A1 => n839, A2 => n1240, B1 => n838, B2 => n1238, 
                           ZN => n840);
   U815 : OAI221_X1 port map( B1 => n1244, B2 => n842, C1 => n1242, C2 => n841,
                           A => n840, ZN => N175);
   U816 : AOI22_X1 port map( A1 => REGISTERS_21_13_port, A2 => n164_port, B1 =>
                           REGISTERS_23_13_port, B2 => n147, ZN => n846);
   U817 : AOI22_X1 port map( A1 => REGISTERS_17_13_port, A2 => n198_port, B1 =>
                           REGISTERS_19_13_port, B2 => n181_port, ZN => n845);
   U818 : AOI22_X1 port map( A1 => REGISTERS_20_13_port, A2 => n232, B1 => 
                           REGISTERS_22_13_port, B2 => n215_port, ZN => n844);
   U819 : AOI22_X1 port map( A1 => REGISTERS_16_13_port, A2 => n266, B1 => 
                           REGISTERS_18_13_port, B2 => n249, ZN => n843);
   U820 : AND4_X1 port map( A1 => n846, A2 => n845, A3 => n844, A4 => n843, ZN 
                           => n863);
   U821 : AOI22_X1 port map( A1 => REGISTERS_29_13_port, A2 => n164_port, B1 =>
                           REGISTERS_31_13_port, B2 => n147, ZN => n850);
   U822 : AOI22_X1 port map( A1 => REGISTERS_25_13_port, A2 => n198_port, B1 =>
                           REGISTERS_27_13_port, B2 => n181_port, ZN => n849);
   U823 : AOI22_X1 port map( A1 => REGISTERS_28_13_port, A2 => n232, B1 => 
                           REGISTERS_30_13_port, B2 => n215_port, ZN => n848);
   U824 : AOI22_X1 port map( A1 => REGISTERS_24_13_port, A2 => n266, B1 => 
                           REGISTERS_26_13_port, B2 => n249, ZN => n847);
   U825 : AND4_X1 port map( A1 => n850, A2 => n849, A3 => n848, A4 => n847, ZN 
                           => n862);
   U826 : AOI22_X1 port map( A1 => REGISTERS_5_13_port, A2 => n164_port, B1 => 
                           REGISTERS_7_13_port, B2 => n147, ZN => n854);
   U827 : AOI22_X1 port map( A1 => REGISTERS_1_13_port, A2 => n198_port, B1 => 
                           REGISTERS_3_13_port, B2 => n181_port, ZN => n853);
   U828 : AOI22_X1 port map( A1 => REGISTERS_4_13_port, A2 => n232, B1 => 
                           REGISTERS_6_13_port, B2 => n215_port, ZN => n852);
   U829 : AOI22_X1 port map( A1 => REGISTERS_0_13_port, A2 => n266, B1 => 
                           REGISTERS_2_13_port, B2 => n249, ZN => n851);
   U830 : NAND4_X1 port map( A1 => n854, A2 => n853, A3 => n852, A4 => n851, ZN
                           => n860);
   U831 : AOI22_X1 port map( A1 => REGISTERS_13_13_port, A2 => n164_port, B1 =>
                           REGISTERS_15_13_port, B2 => n147, ZN => n858);
   U832 : AOI22_X1 port map( A1 => REGISTERS_9_13_port, A2 => n198_port, B1 => 
                           REGISTERS_11_13_port, B2 => n181_port, ZN => n857);
   U833 : AOI22_X1 port map( A1 => REGISTERS_12_13_port, A2 => n232, B1 => 
                           REGISTERS_14_13_port, B2 => n215_port, ZN => n856);
   U834 : AOI22_X1 port map( A1 => REGISTERS_8_13_port, A2 => n266, B1 => 
                           REGISTERS_10_13_port, B2 => n249, ZN => n855);
   U835 : NAND4_X1 port map( A1 => n858, A2 => n857, A3 => n856, A4 => n855, ZN
                           => n859);
   U836 : AOI22_X1 port map( A1 => n860, A2 => n1240, B1 => n859, B2 => n1238, 
                           ZN => n861);
   U837 : OAI221_X1 port map( B1 => n1244, B2 => n863, C1 => n1242, C2 => n862,
                           A => n861, ZN => N174);
   U838 : AOI22_X1 port map( A1 => REGISTERS_21_14_port, A2 => n164_port, B1 =>
                           REGISTERS_23_14_port, B2 => n147, ZN => n867);
   U839 : AOI22_X1 port map( A1 => REGISTERS_17_14_port, A2 => n198_port, B1 =>
                           REGISTERS_19_14_port, B2 => n181_port, ZN => n866);
   U840 : AOI22_X1 port map( A1 => REGISTERS_20_14_port, A2 => n232, B1 => 
                           REGISTERS_22_14_port, B2 => n215_port, ZN => n865);
   U841 : AOI22_X1 port map( A1 => REGISTERS_16_14_port, A2 => n266, B1 => 
                           REGISTERS_18_14_port, B2 => n249, ZN => n864);
   U842 : AND4_X1 port map( A1 => n867, A2 => n866, A3 => n865, A4 => n864, ZN 
                           => n884);
   U843 : AOI22_X1 port map( A1 => REGISTERS_29_14_port, A2 => n164_port, B1 =>
                           REGISTERS_31_14_port, B2 => n147, ZN => n871);
   U844 : AOI22_X1 port map( A1 => REGISTERS_25_14_port, A2 => n198_port, B1 =>
                           REGISTERS_27_14_port, B2 => n181_port, ZN => n870);
   U845 : AOI22_X1 port map( A1 => REGISTERS_28_14_port, A2 => n232, B1 => 
                           REGISTERS_30_14_port, B2 => n215_port, ZN => n869);
   U846 : AOI22_X1 port map( A1 => REGISTERS_24_14_port, A2 => n266, B1 => 
                           REGISTERS_26_14_port, B2 => n249, ZN => n868);
   U847 : AND4_X1 port map( A1 => n871, A2 => n870, A3 => n869, A4 => n868, ZN 
                           => n883);
   U848 : AOI22_X1 port map( A1 => REGISTERS_5_14_port, A2 => n164_port, B1 => 
                           REGISTERS_7_14_port, B2 => n147, ZN => n875);
   U849 : AOI22_X1 port map( A1 => REGISTERS_1_14_port, A2 => n198_port, B1 => 
                           REGISTERS_3_14_port, B2 => n181_port, ZN => n874);
   U850 : AOI22_X1 port map( A1 => REGISTERS_4_14_port, A2 => n232, B1 => 
                           REGISTERS_6_14_port, B2 => n215_port, ZN => n873);
   U851 : AOI22_X1 port map( A1 => REGISTERS_0_14_port, A2 => n266, B1 => 
                           REGISTERS_2_14_port, B2 => n249, ZN => n872);
   U852 : NAND4_X1 port map( A1 => n875, A2 => n874, A3 => n873, A4 => n872, ZN
                           => n881);
   U853 : AOI22_X1 port map( A1 => REGISTERS_13_14_port, A2 => n164_port, B1 =>
                           REGISTERS_15_14_port, B2 => n147, ZN => n879);
   U854 : AOI22_X1 port map( A1 => REGISTERS_9_14_port, A2 => n198_port, B1 => 
                           REGISTERS_11_14_port, B2 => n181_port, ZN => n878);
   U855 : AOI22_X1 port map( A1 => REGISTERS_12_14_port, A2 => n232, B1 => 
                           REGISTERS_14_14_port, B2 => n215_port, ZN => n877);
   U856 : AOI22_X1 port map( A1 => REGISTERS_8_14_port, A2 => n266, B1 => 
                           REGISTERS_10_14_port, B2 => n249, ZN => n876);
   U857 : NAND4_X1 port map( A1 => n879, A2 => n878, A3 => n877, A4 => n876, ZN
                           => n880);
   U858 : AOI22_X1 port map( A1 => n881, A2 => n1240, B1 => n880, B2 => n1238, 
                           ZN => n882);
   U859 : OAI221_X1 port map( B1 => n1244, B2 => n884, C1 => n1242, C2 => n883,
                           A => n882, ZN => N173);
   U860 : AOI22_X1 port map( A1 => REGISTERS_21_15_port, A2 => n165_port, B1 =>
                           REGISTERS_23_15_port, B2 => n148, ZN => n888);
   U861 : AOI22_X1 port map( A1 => REGISTERS_17_15_port, A2 => n199_port, B1 =>
                           REGISTERS_19_15_port, B2 => n182_port, ZN => n887);
   U862 : AOI22_X1 port map( A1 => REGISTERS_20_15_port, A2 => n233, B1 => 
                           REGISTERS_22_15_port, B2 => n216_port, ZN => n886);
   U863 : AOI22_X1 port map( A1 => REGISTERS_16_15_port, A2 => n267, B1 => 
                           REGISTERS_18_15_port, B2 => n250, ZN => n885);
   U864 : AND4_X1 port map( A1 => n888, A2 => n887, A3 => n886, A4 => n885, ZN 
                           => n905);
   U865 : AOI22_X1 port map( A1 => REGISTERS_29_15_port, A2 => n165_port, B1 =>
                           REGISTERS_31_15_port, B2 => n148, ZN => n892);
   U866 : AOI22_X1 port map( A1 => REGISTERS_25_15_port, A2 => n199_port, B1 =>
                           REGISTERS_27_15_port, B2 => n182_port, ZN => n891);
   U867 : AOI22_X1 port map( A1 => REGISTERS_28_15_port, A2 => n233, B1 => 
                           REGISTERS_30_15_port, B2 => n216_port, ZN => n890);
   U868 : AOI22_X1 port map( A1 => REGISTERS_24_15_port, A2 => n267, B1 => 
                           REGISTERS_26_15_port, B2 => n250, ZN => n889);
   U869 : AND4_X1 port map( A1 => n892, A2 => n891, A3 => n890, A4 => n889, ZN 
                           => n904);
   U870 : AOI22_X1 port map( A1 => REGISTERS_5_15_port, A2 => n165_port, B1 => 
                           REGISTERS_7_15_port, B2 => n148, ZN => n896);
   U871 : AOI22_X1 port map( A1 => REGISTERS_1_15_port, A2 => n199_port, B1 => 
                           REGISTERS_3_15_port, B2 => n182_port, ZN => n895);
   U872 : AOI22_X1 port map( A1 => REGISTERS_4_15_port, A2 => n233, B1 => 
                           REGISTERS_6_15_port, B2 => n216_port, ZN => n894);
   U873 : AOI22_X1 port map( A1 => REGISTERS_0_15_port, A2 => n267, B1 => 
                           REGISTERS_2_15_port, B2 => n250, ZN => n893);
   U874 : NAND4_X1 port map( A1 => n896, A2 => n895, A3 => n894, A4 => n893, ZN
                           => n902);
   U875 : AOI22_X1 port map( A1 => REGISTERS_13_15_port, A2 => n165_port, B1 =>
                           REGISTERS_15_15_port, B2 => n148, ZN => n900);
   U876 : AOI22_X1 port map( A1 => REGISTERS_9_15_port, A2 => n199_port, B1 => 
                           REGISTERS_11_15_port, B2 => n182_port, ZN => n899);
   U877 : AOI22_X1 port map( A1 => REGISTERS_12_15_port, A2 => n233, B1 => 
                           REGISTERS_14_15_port, B2 => n216_port, ZN => n898);
   U878 : AOI22_X1 port map( A1 => REGISTERS_8_15_port, A2 => n267, B1 => 
                           REGISTERS_10_15_port, B2 => n250, ZN => n897);
   U879 : NAND4_X1 port map( A1 => n900, A2 => n899, A3 => n898, A4 => n897, ZN
                           => n901);
   U880 : AOI22_X1 port map( A1 => n902, A2 => n1240, B1 => n901, B2 => n1238, 
                           ZN => n903);
   U881 : OAI221_X1 port map( B1 => n1244, B2 => n905, C1 => n1242, C2 => n904,
                           A => n903, ZN => N172);
   U882 : AOI22_X1 port map( A1 => REGISTERS_21_16_port, A2 => n165_port, B1 =>
                           REGISTERS_23_16_port, B2 => n148, ZN => n909);
   U883 : AOI22_X1 port map( A1 => REGISTERS_17_16_port, A2 => n199_port, B1 =>
                           REGISTERS_19_16_port, B2 => n182_port, ZN => n908);
   U884 : AOI22_X1 port map( A1 => REGISTERS_20_16_port, A2 => n233, B1 => 
                           REGISTERS_22_16_port, B2 => n216_port, ZN => n907);
   U885 : AOI22_X1 port map( A1 => REGISTERS_16_16_port, A2 => n267, B1 => 
                           REGISTERS_18_16_port, B2 => n250, ZN => n906);
   U886 : AND4_X1 port map( A1 => n909, A2 => n908, A3 => n907, A4 => n906, ZN 
                           => n926);
   U887 : AOI22_X1 port map( A1 => REGISTERS_29_16_port, A2 => n165_port, B1 =>
                           REGISTERS_31_16_port, B2 => n148, ZN => n913);
   U888 : AOI22_X1 port map( A1 => REGISTERS_25_16_port, A2 => n199_port, B1 =>
                           REGISTERS_27_16_port, B2 => n182_port, ZN => n912);
   U889 : AOI22_X1 port map( A1 => REGISTERS_28_16_port, A2 => n233, B1 => 
                           REGISTERS_30_16_port, B2 => n216_port, ZN => n911);
   U890 : AOI22_X1 port map( A1 => REGISTERS_24_16_port, A2 => n267, B1 => 
                           REGISTERS_26_16_port, B2 => n250, ZN => n910);
   U891 : AND4_X1 port map( A1 => n913, A2 => n912, A3 => n911, A4 => n910, ZN 
                           => n925);
   U892 : AOI22_X1 port map( A1 => REGISTERS_5_16_port, A2 => n165_port, B1 => 
                           REGISTERS_7_16_port, B2 => n148, ZN => n917);
   U893 : AOI22_X1 port map( A1 => REGISTERS_1_16_port, A2 => n199_port, B1 => 
                           REGISTERS_3_16_port, B2 => n182_port, ZN => n916);
   U894 : AOI22_X1 port map( A1 => REGISTERS_4_16_port, A2 => n233, B1 => 
                           REGISTERS_6_16_port, B2 => n216_port, ZN => n915);
   U895 : AOI22_X1 port map( A1 => REGISTERS_0_16_port, A2 => n267, B1 => 
                           REGISTERS_2_16_port, B2 => n250, ZN => n914);
   U896 : NAND4_X1 port map( A1 => n917, A2 => n916, A3 => n915, A4 => n914, ZN
                           => n923);
   U897 : AOI22_X1 port map( A1 => REGISTERS_13_16_port, A2 => n165_port, B1 =>
                           REGISTERS_15_16_port, B2 => n148, ZN => n921);
   U898 : AOI22_X1 port map( A1 => REGISTERS_9_16_port, A2 => n199_port, B1 => 
                           REGISTERS_11_16_port, B2 => n182_port, ZN => n920);
   U899 : AOI22_X1 port map( A1 => REGISTERS_12_16_port, A2 => n233, B1 => 
                           REGISTERS_14_16_port, B2 => n216_port, ZN => n919);
   U900 : AOI22_X1 port map( A1 => REGISTERS_8_16_port, A2 => n267, B1 => 
                           REGISTERS_10_16_port, B2 => n250, ZN => n918);
   U901 : NAND4_X1 port map( A1 => n921, A2 => n920, A3 => n919, A4 => n918, ZN
                           => n922);
   U902 : AOI22_X1 port map( A1 => n923, A2 => n1240, B1 => n922, B2 => n1238, 
                           ZN => n924);
   U903 : OAI221_X1 port map( B1 => n1244, B2 => n926, C1 => n1242, C2 => n925,
                           A => n924, ZN => N171);
   U904 : AOI22_X1 port map( A1 => REGISTERS_21_17_port, A2 => n165_port, B1 =>
                           REGISTERS_23_17_port, B2 => n148, ZN => n930);
   U905 : AOI22_X1 port map( A1 => REGISTERS_17_17_port, A2 => n199_port, B1 =>
                           REGISTERS_19_17_port, B2 => n182_port, ZN => n929);
   U906 : AOI22_X1 port map( A1 => REGISTERS_20_17_port, A2 => n233, B1 => 
                           REGISTERS_22_17_port, B2 => n216_port, ZN => n928);
   U907 : AOI22_X1 port map( A1 => REGISTERS_16_17_port, A2 => n267, B1 => 
                           REGISTERS_18_17_port, B2 => n250, ZN => n927);
   U908 : AND4_X1 port map( A1 => n930, A2 => n929, A3 => n928, A4 => n927, ZN 
                           => n947);
   U909 : AOI22_X1 port map( A1 => REGISTERS_29_17_port, A2 => n165_port, B1 =>
                           REGISTERS_31_17_port, B2 => n148, ZN => n934);
   U910 : AOI22_X1 port map( A1 => REGISTERS_25_17_port, A2 => n199_port, B1 =>
                           REGISTERS_27_17_port, B2 => n182_port, ZN => n933);
   U911 : AOI22_X1 port map( A1 => REGISTERS_28_17_port, A2 => n233, B1 => 
                           REGISTERS_30_17_port, B2 => n216_port, ZN => n932);
   U912 : AOI22_X1 port map( A1 => REGISTERS_24_17_port, A2 => n267, B1 => 
                           REGISTERS_26_17_port, B2 => n250, ZN => n931);
   U913 : AND4_X1 port map( A1 => n934, A2 => n933, A3 => n932, A4 => n931, ZN 
                           => n946);
   U914 : AOI22_X1 port map( A1 => REGISTERS_5_17_port, A2 => n165_port, B1 => 
                           REGISTERS_7_17_port, B2 => n148, ZN => n938);
   U915 : AOI22_X1 port map( A1 => REGISTERS_1_17_port, A2 => n199_port, B1 => 
                           REGISTERS_3_17_port, B2 => n182_port, ZN => n937);
   U916 : AOI22_X1 port map( A1 => REGISTERS_4_17_port, A2 => n233, B1 => 
                           REGISTERS_6_17_port, B2 => n216_port, ZN => n936);
   U917 : AOI22_X1 port map( A1 => REGISTERS_0_17_port, A2 => n267, B1 => 
                           REGISTERS_2_17_port, B2 => n250, ZN => n935);
   U918 : NAND4_X1 port map( A1 => n938, A2 => n937, A3 => n936, A4 => n935, ZN
                           => n944);
   U919 : AOI22_X1 port map( A1 => REGISTERS_13_17_port, A2 => n165_port, B1 =>
                           REGISTERS_15_17_port, B2 => n148, ZN => n942);
   U920 : AOI22_X1 port map( A1 => REGISTERS_9_17_port, A2 => n199_port, B1 => 
                           REGISTERS_11_17_port, B2 => n182_port, ZN => n941);
   U921 : AOI22_X1 port map( A1 => REGISTERS_12_17_port, A2 => n233, B1 => 
                           REGISTERS_14_17_port, B2 => n216_port, ZN => n940);
   U922 : AOI22_X1 port map( A1 => REGISTERS_8_17_port, A2 => n267, B1 => 
                           REGISTERS_10_17_port, B2 => n250, ZN => n939);
   U923 : NAND4_X1 port map( A1 => n942, A2 => n941, A3 => n940, A4 => n939, ZN
                           => n943);
   U924 : AOI22_X1 port map( A1 => n944, A2 => n1240, B1 => n943, B2 => n1238, 
                           ZN => n945);
   U925 : OAI221_X1 port map( B1 => n1244, B2 => n947, C1 => n1242, C2 => n946,
                           A => n945, ZN => N170);
   U926 : AOI22_X1 port map( A1 => REGISTERS_21_18_port, A2 => n166_port, B1 =>
                           REGISTERS_23_18_port, B2 => n149, ZN => n951);
   U927 : AOI22_X1 port map( A1 => REGISTERS_17_18_port, A2 => n200_port, B1 =>
                           REGISTERS_19_18_port, B2 => n183_port, ZN => n950);
   U928 : AOI22_X1 port map( A1 => REGISTERS_20_18_port, A2 => n234, B1 => 
                           REGISTERS_22_18_port, B2 => n217_port, ZN => n949);
   U929 : AOI22_X1 port map( A1 => REGISTERS_16_18_port, A2 => n268, B1 => 
                           REGISTERS_18_18_port, B2 => n251, ZN => n948);
   U930 : AND4_X1 port map( A1 => n951, A2 => n950, A3 => n949, A4 => n948, ZN 
                           => n968);
   U931 : AOI22_X1 port map( A1 => REGISTERS_29_18_port, A2 => n166_port, B1 =>
                           REGISTERS_31_18_port, B2 => n149, ZN => n955);
   U932 : AOI22_X1 port map( A1 => REGISTERS_25_18_port, A2 => n200_port, B1 =>
                           REGISTERS_27_18_port, B2 => n183_port, ZN => n954);
   U933 : AOI22_X1 port map( A1 => REGISTERS_28_18_port, A2 => n234, B1 => 
                           REGISTERS_30_18_port, B2 => n217_port, ZN => n953);
   U934 : AOI22_X1 port map( A1 => REGISTERS_24_18_port, A2 => n268, B1 => 
                           REGISTERS_26_18_port, B2 => n251, ZN => n952);
   U935 : AND4_X1 port map( A1 => n955, A2 => n954, A3 => n953, A4 => n952, ZN 
                           => n967);
   U936 : AOI22_X1 port map( A1 => REGISTERS_5_18_port, A2 => n166_port, B1 => 
                           REGISTERS_7_18_port, B2 => n149, ZN => n959);
   U937 : AOI22_X1 port map( A1 => REGISTERS_1_18_port, A2 => n200_port, B1 => 
                           REGISTERS_3_18_port, B2 => n183_port, ZN => n958);
   U938 : AOI22_X1 port map( A1 => REGISTERS_4_18_port, A2 => n234, B1 => 
                           REGISTERS_6_18_port, B2 => n217_port, ZN => n957);
   U939 : AOI22_X1 port map( A1 => REGISTERS_0_18_port, A2 => n268, B1 => 
                           REGISTERS_2_18_port, B2 => n251, ZN => n956);
   U940 : NAND4_X1 port map( A1 => n959, A2 => n958, A3 => n957, A4 => n956, ZN
                           => n965);
   U941 : AOI22_X1 port map( A1 => REGISTERS_13_18_port, A2 => n166_port, B1 =>
                           REGISTERS_15_18_port, B2 => n149, ZN => n963);
   U942 : AOI22_X1 port map( A1 => REGISTERS_9_18_port, A2 => n200_port, B1 => 
                           REGISTERS_11_18_port, B2 => n183_port, ZN => n962);
   U943 : AOI22_X1 port map( A1 => REGISTERS_12_18_port, A2 => n234, B1 => 
                           REGISTERS_14_18_port, B2 => n217_port, ZN => n961);
   U944 : AOI22_X1 port map( A1 => REGISTERS_8_18_port, A2 => n268, B1 => 
                           REGISTERS_10_18_port, B2 => n251, ZN => n960);
   U945 : NAND4_X1 port map( A1 => n963, A2 => n962, A3 => n961, A4 => n960, ZN
                           => n964);
   U946 : AOI22_X1 port map( A1 => n965, A2 => n1240, B1 => n964, B2 => n1238, 
                           ZN => n966);
   U947 : OAI221_X1 port map( B1 => n1244, B2 => n968, C1 => n1242, C2 => n967,
                           A => n966, ZN => N169);
   U948 : AOI22_X1 port map( A1 => REGISTERS_21_19_port, A2 => n166_port, B1 =>
                           REGISTERS_23_19_port, B2 => n149, ZN => n972);
   U949 : AOI22_X1 port map( A1 => REGISTERS_17_19_port, A2 => n200_port, B1 =>
                           REGISTERS_19_19_port, B2 => n183_port, ZN => n971);
   U950 : AOI22_X1 port map( A1 => REGISTERS_20_19_port, A2 => n234, B1 => 
                           REGISTERS_22_19_port, B2 => n217_port, ZN => n970);
   U951 : AOI22_X1 port map( A1 => REGISTERS_16_19_port, A2 => n268, B1 => 
                           REGISTERS_18_19_port, B2 => n251, ZN => n969);
   U952 : AND4_X1 port map( A1 => n972, A2 => n971, A3 => n970, A4 => n969, ZN 
                           => n989);
   U953 : AOI22_X1 port map( A1 => REGISTERS_29_19_port, A2 => n166_port, B1 =>
                           REGISTERS_31_19_port, B2 => n149, ZN => n976);
   U954 : AOI22_X1 port map( A1 => REGISTERS_25_19_port, A2 => n200_port, B1 =>
                           REGISTERS_27_19_port, B2 => n183_port, ZN => n975);
   U955 : AOI22_X1 port map( A1 => REGISTERS_28_19_port, A2 => n234, B1 => 
                           REGISTERS_30_19_port, B2 => n217_port, ZN => n974);
   U956 : AOI22_X1 port map( A1 => REGISTERS_24_19_port, A2 => n268, B1 => 
                           REGISTERS_26_19_port, B2 => n251, ZN => n973);
   U957 : AND4_X1 port map( A1 => n976, A2 => n975, A3 => n974, A4 => n973, ZN 
                           => n988);
   U958 : AOI22_X1 port map( A1 => REGISTERS_5_19_port, A2 => n166_port, B1 => 
                           REGISTERS_7_19_port, B2 => n149, ZN => n980);
   U959 : AOI22_X1 port map( A1 => REGISTERS_1_19_port, A2 => n200_port, B1 => 
                           REGISTERS_3_19_port, B2 => n183_port, ZN => n979);
   U960 : AOI22_X1 port map( A1 => REGISTERS_4_19_port, A2 => n234, B1 => 
                           REGISTERS_6_19_port, B2 => n217_port, ZN => n978);
   U961 : AOI22_X1 port map( A1 => REGISTERS_0_19_port, A2 => n268, B1 => 
                           REGISTERS_2_19_port, B2 => n251, ZN => n977);
   U962 : NAND4_X1 port map( A1 => n980, A2 => n979, A3 => n978, A4 => n977, ZN
                           => n986);
   U963 : AOI22_X1 port map( A1 => REGISTERS_13_19_port, A2 => n166_port, B1 =>
                           REGISTERS_15_19_port, B2 => n149, ZN => n984);
   U964 : AOI22_X1 port map( A1 => REGISTERS_9_19_port, A2 => n200_port, B1 => 
                           REGISTERS_11_19_port, B2 => n183_port, ZN => n983);
   U965 : AOI22_X1 port map( A1 => REGISTERS_12_19_port, A2 => n234, B1 => 
                           REGISTERS_14_19_port, B2 => n217_port, ZN => n982);
   U966 : AOI22_X1 port map( A1 => REGISTERS_8_19_port, A2 => n268, B1 => 
                           REGISTERS_10_19_port, B2 => n251, ZN => n981);
   U967 : NAND4_X1 port map( A1 => n984, A2 => n983, A3 => n982, A4 => n981, ZN
                           => n985);
   U968 : AOI22_X1 port map( A1 => n986, A2 => n1240, B1 => n985, B2 => n1238, 
                           ZN => n987);
   U969 : OAI221_X1 port map( B1 => n1244, B2 => n989, C1 => n1242, C2 => n988,
                           A => n987, ZN => N168);
   U970 : AOI22_X1 port map( A1 => REGISTERS_21_20_port, A2 => n166_port, B1 =>
                           REGISTERS_23_20_port, B2 => n149, ZN => n993);
   U971 : AOI22_X1 port map( A1 => REGISTERS_17_20_port, A2 => n200_port, B1 =>
                           REGISTERS_19_20_port, B2 => n183_port, ZN => n992);
   U972 : AOI22_X1 port map( A1 => REGISTERS_20_20_port, A2 => n234, B1 => 
                           REGISTERS_22_20_port, B2 => n217_port, ZN => n991);
   U973 : AOI22_X1 port map( A1 => REGISTERS_16_20_port, A2 => n268, B1 => 
                           REGISTERS_18_20_port, B2 => n251, ZN => n990);
   U974 : AND4_X1 port map( A1 => n993, A2 => n992, A3 => n991, A4 => n990, ZN 
                           => n1010);
   U975 : AOI22_X1 port map( A1 => REGISTERS_29_20_port, A2 => n166_port, B1 =>
                           REGISTERS_31_20_port, B2 => n149, ZN => n997);
   U976 : AOI22_X1 port map( A1 => REGISTERS_25_20_port, A2 => n200_port, B1 =>
                           REGISTERS_27_20_port, B2 => n183_port, ZN => n996);
   U977 : AOI22_X1 port map( A1 => REGISTERS_28_20_port, A2 => n234, B1 => 
                           REGISTERS_30_20_port, B2 => n217_port, ZN => n995);
   U978 : AOI22_X1 port map( A1 => REGISTERS_24_20_port, A2 => n268, B1 => 
                           REGISTERS_26_20_port, B2 => n251, ZN => n994);
   U979 : AND4_X1 port map( A1 => n997, A2 => n996, A3 => n995, A4 => n994, ZN 
                           => n1009);
   U980 : AOI22_X1 port map( A1 => REGISTERS_5_20_port, A2 => n166_port, B1 => 
                           REGISTERS_7_20_port, B2 => n149, ZN => n1001);
   U981 : AOI22_X1 port map( A1 => REGISTERS_1_20_port, A2 => n200_port, B1 => 
                           REGISTERS_3_20_port, B2 => n183_port, ZN => n1000);
   U982 : AOI22_X1 port map( A1 => REGISTERS_4_20_port, A2 => n234, B1 => 
                           REGISTERS_6_20_port, B2 => n217_port, ZN => n999);
   U983 : AOI22_X1 port map( A1 => REGISTERS_0_20_port, A2 => n268, B1 => 
                           REGISTERS_2_20_port, B2 => n251, ZN => n998);
   U984 : NAND4_X1 port map( A1 => n1001, A2 => n1000, A3 => n999, A4 => n998, 
                           ZN => n1007);
   U985 : AOI22_X1 port map( A1 => REGISTERS_13_20_port, A2 => n166_port, B1 =>
                           REGISTERS_15_20_port, B2 => n149, ZN => n1005);
   U986 : AOI22_X1 port map( A1 => REGISTERS_9_20_port, A2 => n200_port, B1 => 
                           REGISTERS_11_20_port, B2 => n183_port, ZN => n1004);
   U987 : AOI22_X1 port map( A1 => REGISTERS_12_20_port, A2 => n234, B1 => 
                           REGISTERS_14_20_port, B2 => n217_port, ZN => n1003);
   U988 : AOI22_X1 port map( A1 => REGISTERS_8_20_port, A2 => n268, B1 => 
                           REGISTERS_10_20_port, B2 => n251, ZN => n1002);
   U989 : NAND4_X1 port map( A1 => n1005, A2 => n1004, A3 => n1003, A4 => n1002
                           , ZN => n1006);
   U990 : AOI22_X1 port map( A1 => n1007, A2 => n1240, B1 => n1006, B2 => n1238
                           , ZN => n1008);
   U991 : OAI221_X1 port map( B1 => n1244, B2 => n1010, C1 => n1242, C2 => 
                           n1009, A => n1008, ZN => N167);
   U992 : AOI22_X1 port map( A1 => REGISTERS_21_21_port, A2 => n167_port, B1 =>
                           REGISTERS_23_21_port, B2 => n150, ZN => n1014);
   U993 : AOI22_X1 port map( A1 => REGISTERS_17_21_port, A2 => n201_port, B1 =>
                           REGISTERS_19_21_port, B2 => n184_port, ZN => n1013);
   U994 : AOI22_X1 port map( A1 => REGISTERS_20_21_port, A2 => n235, B1 => 
                           REGISTERS_22_21_port, B2 => n218_port, ZN => n1012);
   U995 : AOI22_X1 port map( A1 => REGISTERS_16_21_port, A2 => n269, B1 => 
                           REGISTERS_18_21_port, B2 => n252, ZN => n1011);
   U996 : AND4_X1 port map( A1 => n1014, A2 => n1013, A3 => n1012, A4 => n1011,
                           ZN => n1031);
   U997 : AOI22_X1 port map( A1 => REGISTERS_29_21_port, A2 => n167_port, B1 =>
                           REGISTERS_31_21_port, B2 => n150, ZN => n1018);
   U998 : AOI22_X1 port map( A1 => REGISTERS_25_21_port, A2 => n201_port, B1 =>
                           REGISTERS_27_21_port, B2 => n184_port, ZN => n1017);
   U999 : AOI22_X1 port map( A1 => REGISTERS_28_21_port, A2 => n235, B1 => 
                           REGISTERS_30_21_port, B2 => n218_port, ZN => n1016);
   U1000 : AOI22_X1 port map( A1 => REGISTERS_24_21_port, A2 => n269, B1 => 
                           REGISTERS_26_21_port, B2 => n252, ZN => n1015);
   U1001 : AND4_X1 port map( A1 => n1018, A2 => n1017, A3 => n1016, A4 => n1015
                           , ZN => n1030);
   U1002 : AOI22_X1 port map( A1 => REGISTERS_5_21_port, A2 => n167_port, B1 =>
                           REGISTERS_7_21_port, B2 => n150, ZN => n1022);
   U1003 : AOI22_X1 port map( A1 => REGISTERS_1_21_port, A2 => n201_port, B1 =>
                           REGISTERS_3_21_port, B2 => n184_port, ZN => n1021);
   U1004 : AOI22_X1 port map( A1 => REGISTERS_4_21_port, A2 => n235, B1 => 
                           REGISTERS_6_21_port, B2 => n218_port, ZN => n1020);
   U1005 : AOI22_X1 port map( A1 => REGISTERS_0_21_port, A2 => n269, B1 => 
                           REGISTERS_2_21_port, B2 => n252, ZN => n1019);
   U1006 : NAND4_X1 port map( A1 => n1022, A2 => n1021, A3 => n1020, A4 => 
                           n1019, ZN => n1028);
   U1007 : AOI22_X1 port map( A1 => REGISTERS_13_21_port, A2 => n167_port, B1 
                           => REGISTERS_15_21_port, B2 => n150, ZN => n1026);
   U1008 : AOI22_X1 port map( A1 => REGISTERS_9_21_port, A2 => n201_port, B1 =>
                           REGISTERS_11_21_port, B2 => n184_port, ZN => n1025);
   U1009 : AOI22_X1 port map( A1 => REGISTERS_12_21_port, A2 => n235, B1 => 
                           REGISTERS_14_21_port, B2 => n218_port, ZN => n1024);
   U1010 : AOI22_X1 port map( A1 => REGISTERS_8_21_port, A2 => n269, B1 => 
                           REGISTERS_10_21_port, B2 => n252, ZN => n1023);
   U1011 : NAND4_X1 port map( A1 => n1026, A2 => n1025, A3 => n1024, A4 => 
                           n1023, ZN => n1027);
   U1012 : AOI22_X1 port map( A1 => n1028, A2 => n1240, B1 => n1027, B2 => 
                           n1238, ZN => n1029);
   U1013 : OAI221_X1 port map( B1 => n1244, B2 => n1031, C1 => n1242, C2 => 
                           n1030, A => n1029, ZN => N166);
   U1014 : AOI22_X1 port map( A1 => REGISTERS_21_22_port, A2 => n167_port, B1 
                           => REGISTERS_23_22_port, B2 => n150, ZN => n1035);
   U1015 : AOI22_X1 port map( A1 => REGISTERS_17_22_port, A2 => n201_port, B1 
                           => REGISTERS_19_22_port, B2 => n184_port, ZN => 
                           n1034);
   U1016 : AOI22_X1 port map( A1 => REGISTERS_20_22_port, A2 => n235, B1 => 
                           REGISTERS_22_22_port, B2 => n218_port, ZN => n1033);
   U1017 : AOI22_X1 port map( A1 => REGISTERS_16_22_port, A2 => n269, B1 => 
                           REGISTERS_18_22_port, B2 => n252, ZN => n1032);
   U1018 : AND4_X1 port map( A1 => n1035, A2 => n1034, A3 => n1033, A4 => n1032
                           , ZN => n1052);
   U1019 : AOI22_X1 port map( A1 => REGISTERS_29_22_port, A2 => n167_port, B1 
                           => REGISTERS_31_22_port, B2 => n150, ZN => n1039);
   U1020 : AOI22_X1 port map( A1 => REGISTERS_25_22_port, A2 => n201_port, B1 
                           => REGISTERS_27_22_port, B2 => n184_port, ZN => 
                           n1038);
   U1021 : AOI22_X1 port map( A1 => REGISTERS_28_22_port, A2 => n235, B1 => 
                           REGISTERS_30_22_port, B2 => n218_port, ZN => n1037);
   U1022 : AOI22_X1 port map( A1 => REGISTERS_24_22_port, A2 => n269, B1 => 
                           REGISTERS_26_22_port, B2 => n252, ZN => n1036);
   U1023 : AND4_X1 port map( A1 => n1039, A2 => n1038, A3 => n1037, A4 => n1036
                           , ZN => n1051);
   U1024 : AOI22_X1 port map( A1 => REGISTERS_5_22_port, A2 => n167_port, B1 =>
                           REGISTERS_7_22_port, B2 => n150, ZN => n1043);
   U1025 : AOI22_X1 port map( A1 => REGISTERS_1_22_port, A2 => n201_port, B1 =>
                           REGISTERS_3_22_port, B2 => n184_port, ZN => n1042);
   U1026 : AOI22_X1 port map( A1 => REGISTERS_4_22_port, A2 => n235, B1 => 
                           REGISTERS_6_22_port, B2 => n218_port, ZN => n1041);
   U1027 : AOI22_X1 port map( A1 => REGISTERS_0_22_port, A2 => n269, B1 => 
                           REGISTERS_2_22_port, B2 => n252, ZN => n1040);
   U1028 : NAND4_X1 port map( A1 => n1043, A2 => n1042, A3 => n1041, A4 => 
                           n1040, ZN => n1049);
   U1029 : AOI22_X1 port map( A1 => REGISTERS_13_22_port, A2 => n167_port, B1 
                           => REGISTERS_15_22_port, B2 => n150, ZN => n1047);
   U1030 : AOI22_X1 port map( A1 => REGISTERS_9_22_port, A2 => n201_port, B1 =>
                           REGISTERS_11_22_port, B2 => n184_port, ZN => n1046);
   U1031 : AOI22_X1 port map( A1 => REGISTERS_12_22_port, A2 => n235, B1 => 
                           REGISTERS_14_22_port, B2 => n218_port, ZN => n1045);
   U1032 : AOI22_X1 port map( A1 => REGISTERS_8_22_port, A2 => n269, B1 => 
                           REGISTERS_10_22_port, B2 => n252, ZN => n1044);
   U1033 : NAND4_X1 port map( A1 => n1047, A2 => n1046, A3 => n1045, A4 => 
                           n1044, ZN => n1048);
   U1034 : AOI22_X1 port map( A1 => n1049, A2 => n1240, B1 => n1048, B2 => 
                           n1238, ZN => n1050);
   U1035 : OAI221_X1 port map( B1 => n1244, B2 => n1052, C1 => n1242, C2 => 
                           n1051, A => n1050, ZN => N165);
   U1036 : AOI22_X1 port map( A1 => REGISTERS_21_23_port, A2 => n167_port, B1 
                           => REGISTERS_23_23_port, B2 => n150, ZN => n1056);
   U1037 : AOI22_X1 port map( A1 => REGISTERS_17_23_port, A2 => n201_port, B1 
                           => REGISTERS_19_23_port, B2 => n184_port, ZN => 
                           n1055);
   U1038 : AOI22_X1 port map( A1 => REGISTERS_20_23_port, A2 => n235, B1 => 
                           REGISTERS_22_23_port, B2 => n218_port, ZN => n1054);
   U1039 : AOI22_X1 port map( A1 => REGISTERS_16_23_port, A2 => n269, B1 => 
                           REGISTERS_18_23_port, B2 => n252, ZN => n1053);
   U1040 : AND4_X1 port map( A1 => n1056, A2 => n1055, A3 => n1054, A4 => n1053
                           , ZN => n1073);
   U1041 : AOI22_X1 port map( A1 => REGISTERS_29_23_port, A2 => n167_port, B1 
                           => REGISTERS_31_23_port, B2 => n150, ZN => n1060);
   U1042 : AOI22_X1 port map( A1 => REGISTERS_25_23_port, A2 => n201_port, B1 
                           => REGISTERS_27_23_port, B2 => n184_port, ZN => 
                           n1059);
   U1043 : AOI22_X1 port map( A1 => REGISTERS_28_23_port, A2 => n235, B1 => 
                           REGISTERS_30_23_port, B2 => n218_port, ZN => n1058);
   U1044 : AOI22_X1 port map( A1 => REGISTERS_24_23_port, A2 => n269, B1 => 
                           REGISTERS_26_23_port, B2 => n252, ZN => n1057);
   U1045 : AND4_X1 port map( A1 => n1060, A2 => n1059, A3 => n1058, A4 => n1057
                           , ZN => n1072);
   U1046 : AOI22_X1 port map( A1 => REGISTERS_5_23_port, A2 => n167_port, B1 =>
                           REGISTERS_7_23_port, B2 => n150, ZN => n1064);
   U1047 : AOI22_X1 port map( A1 => REGISTERS_1_23_port, A2 => n201_port, B1 =>
                           REGISTERS_3_23_port, B2 => n184_port, ZN => n1063);
   U1048 : AOI22_X1 port map( A1 => REGISTERS_4_23_port, A2 => n235, B1 => 
                           REGISTERS_6_23_port, B2 => n218_port, ZN => n1062);
   U1049 : AOI22_X1 port map( A1 => REGISTERS_0_23_port, A2 => n269, B1 => 
                           REGISTERS_2_23_port, B2 => n252, ZN => n1061);
   U1050 : NAND4_X1 port map( A1 => n1064, A2 => n1063, A3 => n1062, A4 => 
                           n1061, ZN => n1070);
   U1051 : AOI22_X1 port map( A1 => REGISTERS_13_23_port, A2 => n167_port, B1 
                           => REGISTERS_15_23_port, B2 => n150, ZN => n1068);
   U1052 : AOI22_X1 port map( A1 => REGISTERS_9_23_port, A2 => n201_port, B1 =>
                           REGISTERS_11_23_port, B2 => n184_port, ZN => n1067);
   U1053 : AOI22_X1 port map( A1 => REGISTERS_12_23_port, A2 => n235, B1 => 
                           REGISTERS_14_23_port, B2 => n218_port, ZN => n1066);
   U1054 : AOI22_X1 port map( A1 => REGISTERS_8_23_port, A2 => n269, B1 => 
                           REGISTERS_10_23_port, B2 => n252, ZN => n1065);
   U1055 : NAND4_X1 port map( A1 => n1068, A2 => n1067, A3 => n1066, A4 => 
                           n1065, ZN => n1069);
   U1056 : AOI22_X1 port map( A1 => n1070, A2 => n1240, B1 => n1069, B2 => 
                           n1238, ZN => n1071);
   U1057 : OAI221_X1 port map( B1 => n1244, B2 => n1073, C1 => n1242, C2 => 
                           n1072, A => n1071, ZN => N164);
   U1058 : AOI22_X1 port map( A1 => REGISTERS_21_24_port, A2 => n168_port, B1 
                           => REGISTERS_23_24_port, B2 => n151, ZN => n1077);
   U1059 : AOI22_X1 port map( A1 => REGISTERS_17_24_port, A2 => n202_port, B1 
                           => REGISTERS_19_24_port, B2 => n185_port, ZN => 
                           n1076);
   U1060 : AOI22_X1 port map( A1 => REGISTERS_20_24_port, A2 => n236, B1 => 
                           REGISTERS_22_24_port, B2 => n219_port, ZN => n1075);
   U1061 : AOI22_X1 port map( A1 => REGISTERS_16_24_port, A2 => n270, B1 => 
                           REGISTERS_18_24_port, B2 => n253, ZN => n1074);
   U1062 : AND4_X1 port map( A1 => n1077, A2 => n1076, A3 => n1075, A4 => n1074
                           , ZN => n1094);
   U1063 : AOI22_X1 port map( A1 => REGISTERS_29_24_port, A2 => n168_port, B1 
                           => REGISTERS_31_24_port, B2 => n151, ZN => n1081);
   U1064 : AOI22_X1 port map( A1 => REGISTERS_25_24_port, A2 => n202_port, B1 
                           => REGISTERS_27_24_port, B2 => n185_port, ZN => 
                           n1080);
   U1065 : AOI22_X1 port map( A1 => REGISTERS_28_24_port, A2 => n236, B1 => 
                           REGISTERS_30_24_port, B2 => n219_port, ZN => n1079);
   U1066 : AOI22_X1 port map( A1 => REGISTERS_24_24_port, A2 => n270, B1 => 
                           REGISTERS_26_24_port, B2 => n253, ZN => n1078);
   U1067 : AND4_X1 port map( A1 => n1081, A2 => n1080, A3 => n1079, A4 => n1078
                           , ZN => n1093);
   U1068 : AOI22_X1 port map( A1 => REGISTERS_5_24_port, A2 => n168_port, B1 =>
                           REGISTERS_7_24_port, B2 => n151, ZN => n1085);
   U1069 : AOI22_X1 port map( A1 => REGISTERS_1_24_port, A2 => n202_port, B1 =>
                           REGISTERS_3_24_port, B2 => n185_port, ZN => n1084);
   U1070 : AOI22_X1 port map( A1 => REGISTERS_4_24_port, A2 => n236, B1 => 
                           REGISTERS_6_24_port, B2 => n219_port, ZN => n1083);
   U1071 : AOI22_X1 port map( A1 => REGISTERS_0_24_port, A2 => n270, B1 => 
                           REGISTERS_2_24_port, B2 => n253, ZN => n1082);
   U1072 : NAND4_X1 port map( A1 => n1085, A2 => n1084, A3 => n1083, A4 => 
                           n1082, ZN => n1091);
   U1073 : AOI22_X1 port map( A1 => REGISTERS_13_24_port, A2 => n168_port, B1 
                           => REGISTERS_15_24_port, B2 => n151, ZN => n1089);
   U1074 : AOI22_X1 port map( A1 => REGISTERS_9_24_port, A2 => n202_port, B1 =>
                           REGISTERS_11_24_port, B2 => n185_port, ZN => n1088);
   U1075 : AOI22_X1 port map( A1 => REGISTERS_12_24_port, A2 => n236, B1 => 
                           REGISTERS_14_24_port, B2 => n219_port, ZN => n1087);
   U1076 : AOI22_X1 port map( A1 => REGISTERS_8_24_port, A2 => n270, B1 => 
                           REGISTERS_10_24_port, B2 => n253, ZN => n1086);
   U1077 : NAND4_X1 port map( A1 => n1089, A2 => n1088, A3 => n1087, A4 => 
                           n1086, ZN => n1090);
   U1078 : AOI22_X1 port map( A1 => n1091, A2 => n1240, B1 => n1090, B2 => 
                           n1238, ZN => n1092);
   U1079 : OAI221_X1 port map( B1 => n1244, B2 => n1094, C1 => n1242, C2 => 
                           n1093, A => n1092, ZN => N163);
   U1080 : AOI22_X1 port map( A1 => REGISTERS_21_25_port, A2 => n168_port, B1 
                           => REGISTERS_23_25_port, B2 => n151, ZN => n1098);
   U1081 : AOI22_X1 port map( A1 => REGISTERS_17_25_port, A2 => n202_port, B1 
                           => REGISTERS_19_25_port, B2 => n185_port, ZN => 
                           n1097);
   U1082 : AOI22_X1 port map( A1 => REGISTERS_20_25_port, A2 => n236, B1 => 
                           REGISTERS_22_25_port, B2 => n219_port, ZN => n1096);
   U1083 : AOI22_X1 port map( A1 => REGISTERS_16_25_port, A2 => n270, B1 => 
                           REGISTERS_18_25_port, B2 => n253, ZN => n1095);
   U1084 : AND4_X1 port map( A1 => n1098, A2 => n1097, A3 => n1096, A4 => n1095
                           , ZN => n1115);
   U1085 : AOI22_X1 port map( A1 => REGISTERS_29_25_port, A2 => n168_port, B1 
                           => REGISTERS_31_25_port, B2 => n151, ZN => n1102);
   U1086 : AOI22_X1 port map( A1 => REGISTERS_25_25_port, A2 => n202_port, B1 
                           => REGISTERS_27_25_port, B2 => n185_port, ZN => 
                           n1101);
   U1087 : AOI22_X1 port map( A1 => REGISTERS_28_25_port, A2 => n236, B1 => 
                           REGISTERS_30_25_port, B2 => n219_port, ZN => n1100);
   U1088 : AOI22_X1 port map( A1 => REGISTERS_24_25_port, A2 => n270, B1 => 
                           REGISTERS_26_25_port, B2 => n253, ZN => n1099);
   U1089 : AND4_X1 port map( A1 => n1102, A2 => n1101, A3 => n1100, A4 => n1099
                           , ZN => n1114);
   U1090 : AOI22_X1 port map( A1 => REGISTERS_5_25_port, A2 => n168_port, B1 =>
                           REGISTERS_7_25_port, B2 => n151, ZN => n1106);
   U1091 : AOI22_X1 port map( A1 => REGISTERS_1_25_port, A2 => n202_port, B1 =>
                           REGISTERS_3_25_port, B2 => n185_port, ZN => n1105);
   U1092 : AOI22_X1 port map( A1 => REGISTERS_4_25_port, A2 => n236, B1 => 
                           REGISTERS_6_25_port, B2 => n219_port, ZN => n1104);
   U1093 : AOI22_X1 port map( A1 => REGISTERS_0_25_port, A2 => n270, B1 => 
                           REGISTERS_2_25_port, B2 => n253, ZN => n1103);
   U1094 : NAND4_X1 port map( A1 => n1106, A2 => n1105, A3 => n1104, A4 => 
                           n1103, ZN => n1112);
   U1095 : AOI22_X1 port map( A1 => REGISTERS_13_25_port, A2 => n168_port, B1 
                           => REGISTERS_15_25_port, B2 => n151, ZN => n1110);
   U1096 : AOI22_X1 port map( A1 => REGISTERS_9_25_port, A2 => n202_port, B1 =>
                           REGISTERS_11_25_port, B2 => n185_port, ZN => n1109);
   U1097 : AOI22_X1 port map( A1 => REGISTERS_12_25_port, A2 => n236, B1 => 
                           REGISTERS_14_25_port, B2 => n219_port, ZN => n1108);
   U1098 : AOI22_X1 port map( A1 => REGISTERS_8_25_port, A2 => n270, B1 => 
                           REGISTERS_10_25_port, B2 => n253, ZN => n1107);
   U1099 : NAND4_X1 port map( A1 => n1110, A2 => n1109, A3 => n1108, A4 => 
                           n1107, ZN => n1111);
   U1100 : AOI22_X1 port map( A1 => n1112, A2 => n1240, B1 => n1111, B2 => 
                           n1238, ZN => n1113);
   U1101 : OAI221_X1 port map( B1 => n1244, B2 => n1115, C1 => n1242, C2 => 
                           n1114, A => n1113, ZN => N162);
   U1102 : AOI22_X1 port map( A1 => REGISTERS_21_26_port, A2 => n168_port, B1 
                           => REGISTERS_23_26_port, B2 => n151, ZN => n1119);
   U1103 : AOI22_X1 port map( A1 => REGISTERS_17_26_port, A2 => n202_port, B1 
                           => REGISTERS_19_26_port, B2 => n185_port, ZN => 
                           n1118);
   U1104 : AOI22_X1 port map( A1 => REGISTERS_20_26_port, A2 => n236, B1 => 
                           REGISTERS_22_26_port, B2 => n219_port, ZN => n1117);
   U1105 : AOI22_X1 port map( A1 => REGISTERS_16_26_port, A2 => n270, B1 => 
                           REGISTERS_18_26_port, B2 => n253, ZN => n1116);
   U1106 : AND4_X1 port map( A1 => n1119, A2 => n1118, A3 => n1117, A4 => n1116
                           , ZN => n1136);
   U1107 : AOI22_X1 port map( A1 => REGISTERS_29_26_port, A2 => n168_port, B1 
                           => REGISTERS_31_26_port, B2 => n151, ZN => n1123);
   U1108 : AOI22_X1 port map( A1 => REGISTERS_25_26_port, A2 => n202_port, B1 
                           => REGISTERS_27_26_port, B2 => n185_port, ZN => 
                           n1122);
   U1109 : AOI22_X1 port map( A1 => REGISTERS_28_26_port, A2 => n236, B1 => 
                           REGISTERS_30_26_port, B2 => n219_port, ZN => n1121);
   U1110 : AOI22_X1 port map( A1 => REGISTERS_24_26_port, A2 => n270, B1 => 
                           REGISTERS_26_26_port, B2 => n253, ZN => n1120);
   U1111 : AND4_X1 port map( A1 => n1123, A2 => n1122, A3 => n1121, A4 => n1120
                           , ZN => n1135);
   U1112 : AOI22_X1 port map( A1 => REGISTERS_5_26_port, A2 => n168_port, B1 =>
                           REGISTERS_7_26_port, B2 => n151, ZN => n1127);
   U1113 : AOI22_X1 port map( A1 => REGISTERS_1_26_port, A2 => n202_port, B1 =>
                           REGISTERS_3_26_port, B2 => n185_port, ZN => n1126);
   U1114 : AOI22_X1 port map( A1 => REGISTERS_4_26_port, A2 => n236, B1 => 
                           REGISTERS_6_26_port, B2 => n219_port, ZN => n1125);
   U1115 : AOI22_X1 port map( A1 => REGISTERS_0_26_port, A2 => n270, B1 => 
                           REGISTERS_2_26_port, B2 => n253, ZN => n1124);
   U1116 : NAND4_X1 port map( A1 => n1127, A2 => n1126, A3 => n1125, A4 => 
                           n1124, ZN => n1133);
   U1117 : AOI22_X1 port map( A1 => REGISTERS_13_26_port, A2 => n168_port, B1 
                           => REGISTERS_15_26_port, B2 => n151, ZN => n1131);
   U1118 : AOI22_X1 port map( A1 => REGISTERS_9_26_port, A2 => n202_port, B1 =>
                           REGISTERS_11_26_port, B2 => n185_port, ZN => n1130);
   U1119 : AOI22_X1 port map( A1 => REGISTERS_12_26_port, A2 => n236, B1 => 
                           REGISTERS_14_26_port, B2 => n219_port, ZN => n1129);
   U1120 : AOI22_X1 port map( A1 => REGISTERS_8_26_port, A2 => n270, B1 => 
                           REGISTERS_10_26_port, B2 => n253, ZN => n1128);
   U1121 : NAND4_X1 port map( A1 => n1131, A2 => n1130, A3 => n1129, A4 => 
                           n1128, ZN => n1132);
   U1122 : AOI22_X1 port map( A1 => n1133, A2 => n1240, B1 => n1132, B2 => 
                           n1238, ZN => n1134);
   U1123 : OAI221_X1 port map( B1 => n1244, B2 => n1136, C1 => n1242, C2 => 
                           n1135, A => n1134, ZN => N161);
   U1124 : AOI22_X1 port map( A1 => REGISTERS_21_27_port, A2 => n169_port, B1 
                           => REGISTERS_23_27_port, B2 => n152, ZN => n1140);
   U1125 : AOI22_X1 port map( A1 => REGISTERS_17_27_port, A2 => n203_port, B1 
                           => REGISTERS_19_27_port, B2 => n186_port, ZN => 
                           n1139);
   U1126 : AOI22_X1 port map( A1 => REGISTERS_20_27_port, A2 => n237, B1 => 
                           REGISTERS_22_27_port, B2 => n220_port, ZN => n1138);
   U1127 : AOI22_X1 port map( A1 => REGISTERS_16_27_port, A2 => n271, B1 => 
                           REGISTERS_18_27_port, B2 => n254, ZN => n1137);
   U1128 : AND4_X1 port map( A1 => n1140, A2 => n1139, A3 => n1138, A4 => n1137
                           , ZN => n1157);
   U1129 : AOI22_X1 port map( A1 => REGISTERS_29_27_port, A2 => n169_port, B1 
                           => REGISTERS_31_27_port, B2 => n152, ZN => n1144);
   U1130 : AOI22_X1 port map( A1 => REGISTERS_25_27_port, A2 => n203_port, B1 
                           => REGISTERS_27_27_port, B2 => n186_port, ZN => 
                           n1143);
   U1131 : AOI22_X1 port map( A1 => REGISTERS_28_27_port, A2 => n237, B1 => 
                           REGISTERS_30_27_port, B2 => n220_port, ZN => n1142);
   U1132 : AOI22_X1 port map( A1 => REGISTERS_24_27_port, A2 => n271, B1 => 
                           REGISTERS_26_27_port, B2 => n254, ZN => n1141);
   U1133 : AND4_X1 port map( A1 => n1144, A2 => n1143, A3 => n1142, A4 => n1141
                           , ZN => n1156);
   U1134 : AOI22_X1 port map( A1 => REGISTERS_5_27_port, A2 => n169_port, B1 =>
                           REGISTERS_7_27_port, B2 => n152, ZN => n1148);
   U1135 : AOI22_X1 port map( A1 => REGISTERS_1_27_port, A2 => n203_port, B1 =>
                           REGISTERS_3_27_port, B2 => n186_port, ZN => n1147);
   U1136 : AOI22_X1 port map( A1 => REGISTERS_4_27_port, A2 => n237, B1 => 
                           REGISTERS_6_27_port, B2 => n220_port, ZN => n1146);
   U1137 : AOI22_X1 port map( A1 => REGISTERS_0_27_port, A2 => n271, B1 => 
                           REGISTERS_2_27_port, B2 => n254, ZN => n1145);
   U1138 : NAND4_X1 port map( A1 => n1148, A2 => n1147, A3 => n1146, A4 => 
                           n1145, ZN => n1154);
   U1139 : AOI22_X1 port map( A1 => REGISTERS_13_27_port, A2 => n169_port, B1 
                           => REGISTERS_15_27_port, B2 => n152, ZN => n1152);
   U1140 : AOI22_X1 port map( A1 => REGISTERS_9_27_port, A2 => n203_port, B1 =>
                           REGISTERS_11_27_port, B2 => n186_port, ZN => n1151);
   U1141 : AOI22_X1 port map( A1 => REGISTERS_12_27_port, A2 => n237, B1 => 
                           REGISTERS_14_27_port, B2 => n220_port, ZN => n1150);
   U1142 : AOI22_X1 port map( A1 => REGISTERS_8_27_port, A2 => n271, B1 => 
                           REGISTERS_10_27_port, B2 => n254, ZN => n1149);
   U1143 : NAND4_X1 port map( A1 => n1152, A2 => n1151, A3 => n1150, A4 => 
                           n1149, ZN => n1153);
   U1144 : AOI22_X1 port map( A1 => n1154, A2 => n1240, B1 => n1153, B2 => 
                           n1238, ZN => n1155);
   U1145 : OAI221_X1 port map( B1 => n1244, B2 => n1157, C1 => n1242, C2 => 
                           n1156, A => n1155, ZN => N160);
   U1146 : AOI22_X1 port map( A1 => REGISTERS_21_28_port, A2 => n169_port, B1 
                           => REGISTERS_23_28_port, B2 => n152, ZN => n1161);
   U1147 : AOI22_X1 port map( A1 => REGISTERS_17_28_port, A2 => n203_port, B1 
                           => REGISTERS_19_28_port, B2 => n186_port, ZN => 
                           n1160);
   U1148 : AOI22_X1 port map( A1 => REGISTERS_20_28_port, A2 => n237, B1 => 
                           REGISTERS_22_28_port, B2 => n220_port, ZN => n1159);
   U1149 : AOI22_X1 port map( A1 => REGISTERS_16_28_port, A2 => n271, B1 => 
                           REGISTERS_18_28_port, B2 => n254, ZN => n1158);
   U1150 : AND4_X1 port map( A1 => n1161, A2 => n1160, A3 => n1159, A4 => n1158
                           , ZN => n1178);
   U1151 : AOI22_X1 port map( A1 => REGISTERS_29_28_port, A2 => n169_port, B1 
                           => REGISTERS_31_28_port, B2 => n152, ZN => n1165);
   U1152 : AOI22_X1 port map( A1 => REGISTERS_25_28_port, A2 => n203_port, B1 
                           => REGISTERS_27_28_port, B2 => n186_port, ZN => 
                           n1164);
   U1153 : AOI22_X1 port map( A1 => REGISTERS_28_28_port, A2 => n237, B1 => 
                           REGISTERS_30_28_port, B2 => n220_port, ZN => n1163);
   U1154 : AOI22_X1 port map( A1 => REGISTERS_24_28_port, A2 => n271, B1 => 
                           REGISTERS_26_28_port, B2 => n254, ZN => n1162);
   U1155 : AND4_X1 port map( A1 => n1165, A2 => n1164, A3 => n1163, A4 => n1162
                           , ZN => n1177);
   U1156 : AOI22_X1 port map( A1 => REGISTERS_5_28_port, A2 => n169_port, B1 =>
                           REGISTERS_7_28_port, B2 => n152, ZN => n1169);
   U1157 : AOI22_X1 port map( A1 => REGISTERS_1_28_port, A2 => n203_port, B1 =>
                           REGISTERS_3_28_port, B2 => n186_port, ZN => n1168);
   U1158 : AOI22_X1 port map( A1 => REGISTERS_4_28_port, A2 => n237, B1 => 
                           REGISTERS_6_28_port, B2 => n220_port, ZN => n1167);
   U1159 : AOI22_X1 port map( A1 => REGISTERS_0_28_port, A2 => n271, B1 => 
                           REGISTERS_2_28_port, B2 => n254, ZN => n1166);
   U1160 : NAND4_X1 port map( A1 => n1169, A2 => n1168, A3 => n1167, A4 => 
                           n1166, ZN => n1175);
   U1161 : AOI22_X1 port map( A1 => REGISTERS_13_28_port, A2 => n169_port, B1 
                           => REGISTERS_15_28_port, B2 => n152, ZN => n1173);
   U1162 : AOI22_X1 port map( A1 => REGISTERS_9_28_port, A2 => n203_port, B1 =>
                           REGISTERS_11_28_port, B2 => n186_port, ZN => n1172);
   U1163 : AOI22_X1 port map( A1 => REGISTERS_12_28_port, A2 => n237, B1 => 
                           REGISTERS_14_28_port, B2 => n220_port, ZN => n1171);
   U1164 : AOI22_X1 port map( A1 => REGISTERS_8_28_port, A2 => n271, B1 => 
                           REGISTERS_10_28_port, B2 => n254, ZN => n1170);
   U1165 : NAND4_X1 port map( A1 => n1173, A2 => n1172, A3 => n1171, A4 => 
                           n1170, ZN => n1174);
   U1166 : AOI22_X1 port map( A1 => n1175, A2 => n1240, B1 => n1174, B2 => 
                           n1238, ZN => n1176);
   U1167 : OAI221_X1 port map( B1 => n1244, B2 => n1178, C1 => n1242, C2 => 
                           n1177, A => n1176, ZN => N159);
   U1168 : AOI22_X1 port map( A1 => REGISTERS_21_29_port, A2 => n169_port, B1 
                           => REGISTERS_23_29_port, B2 => n152, ZN => n1182);
   U1169 : AOI22_X1 port map( A1 => REGISTERS_17_29_port, A2 => n203_port, B1 
                           => REGISTERS_19_29_port, B2 => n186_port, ZN => 
                           n1181);
   U1170 : AOI22_X1 port map( A1 => REGISTERS_20_29_port, A2 => n237, B1 => 
                           REGISTERS_22_29_port, B2 => n220_port, ZN => n1180);
   U1171 : AOI22_X1 port map( A1 => REGISTERS_16_29_port, A2 => n271, B1 => 
                           REGISTERS_18_29_port, B2 => n254, ZN => n1179);
   U1172 : AND4_X1 port map( A1 => n1182, A2 => n1181, A3 => n1180, A4 => n1179
                           , ZN => n1199);
   U1173 : AOI22_X1 port map( A1 => REGISTERS_29_29_port, A2 => n169_port, B1 
                           => REGISTERS_31_29_port, B2 => n152, ZN => n1186);
   U1174 : AOI22_X1 port map( A1 => REGISTERS_25_29_port, A2 => n203_port, B1 
                           => REGISTERS_27_29_port, B2 => n186_port, ZN => 
                           n1185);
   U1175 : AOI22_X1 port map( A1 => REGISTERS_28_29_port, A2 => n237, B1 => 
                           REGISTERS_30_29_port, B2 => n220_port, ZN => n1184);
   U1176 : AOI22_X1 port map( A1 => REGISTERS_24_29_port, A2 => n271, B1 => 
                           REGISTERS_26_29_port, B2 => n254, ZN => n1183);
   U1177 : AND4_X1 port map( A1 => n1186, A2 => n1185, A3 => n1184, A4 => n1183
                           , ZN => n1198);
   U1178 : AOI22_X1 port map( A1 => REGISTERS_5_29_port, A2 => n169_port, B1 =>
                           REGISTERS_7_29_port, B2 => n152, ZN => n1190);
   U1179 : AOI22_X1 port map( A1 => REGISTERS_1_29_port, A2 => n203_port, B1 =>
                           REGISTERS_3_29_port, B2 => n186_port, ZN => n1189);
   U1180 : AOI22_X1 port map( A1 => REGISTERS_4_29_port, A2 => n237, B1 => 
                           REGISTERS_6_29_port, B2 => n220_port, ZN => n1188);
   U1181 : AOI22_X1 port map( A1 => REGISTERS_0_29_port, A2 => n271, B1 => 
                           REGISTERS_2_29_port, B2 => n254, ZN => n1187);
   U1182 : NAND4_X1 port map( A1 => n1190, A2 => n1189, A3 => n1188, A4 => 
                           n1187, ZN => n1196);
   U1183 : AOI22_X1 port map( A1 => REGISTERS_13_29_port, A2 => n169_port, B1 
                           => REGISTERS_15_29_port, B2 => n152, ZN => n1194);
   U1184 : AOI22_X1 port map( A1 => REGISTERS_9_29_port, A2 => n203_port, B1 =>
                           REGISTERS_11_29_port, B2 => n186_port, ZN => n1193);
   U1185 : AOI22_X1 port map( A1 => REGISTERS_12_29_port, A2 => n237, B1 => 
                           REGISTERS_14_29_port, B2 => n220_port, ZN => n1192);
   U1186 : AOI22_X1 port map( A1 => REGISTERS_8_29_port, A2 => n271, B1 => 
                           REGISTERS_10_29_port, B2 => n254, ZN => n1191);
   U1187 : NAND4_X1 port map( A1 => n1194, A2 => n1193, A3 => n1192, A4 => 
                           n1191, ZN => n1195);
   U1188 : AOI22_X1 port map( A1 => n1196, A2 => n1240, B1 => n1195, B2 => 
                           n1238, ZN => n1197);
   U1189 : OAI221_X1 port map( B1 => n1244, B2 => n1199, C1 => n1242, C2 => 
                           n1198, A => n1197, ZN => N158);
   U1190 : AOI22_X1 port map( A1 => REGISTERS_21_30_port, A2 => n170_port, B1 
                           => REGISTERS_23_30_port, B2 => n153, ZN => n1203);
   U1191 : AOI22_X1 port map( A1 => REGISTERS_17_30_port, A2 => n204_port, B1 
                           => REGISTERS_19_30_port, B2 => n187_port, ZN => 
                           n1202);
   U1192 : AOI22_X1 port map( A1 => REGISTERS_20_30_port, A2 => n238, B1 => 
                           REGISTERS_22_30_port, B2 => n221, ZN => n1201);
   U1193 : AOI22_X1 port map( A1 => REGISTERS_16_30_port, A2 => n272, B1 => 
                           REGISTERS_18_30_port, B2 => n255, ZN => n1200);
   U1194 : AND4_X1 port map( A1 => n1203, A2 => n1202, A3 => n1201, A4 => n1200
                           , ZN => n1220);
   U1195 : AOI22_X1 port map( A1 => REGISTERS_29_30_port, A2 => n170_port, B1 
                           => REGISTERS_31_30_port, B2 => n153, ZN => n1207);
   U1196 : AOI22_X1 port map( A1 => REGISTERS_25_30_port, A2 => n204_port, B1 
                           => REGISTERS_27_30_port, B2 => n187_port, ZN => 
                           n1206);
   U1197 : AOI22_X1 port map( A1 => REGISTERS_28_30_port, A2 => n238, B1 => 
                           REGISTERS_30_30_port, B2 => n221, ZN => n1205);
   U1198 : AOI22_X1 port map( A1 => REGISTERS_24_30_port, A2 => n272, B1 => 
                           REGISTERS_26_30_port, B2 => n255, ZN => n1204);
   U1199 : AND4_X1 port map( A1 => n1207, A2 => n1206, A3 => n1205, A4 => n1204
                           , ZN => n1219);
   U1200 : AOI22_X1 port map( A1 => REGISTERS_5_30_port, A2 => n170_port, B1 =>
                           REGISTERS_7_30_port, B2 => n153, ZN => n1211);
   U1201 : AOI22_X1 port map( A1 => REGISTERS_1_30_port, A2 => n204_port, B1 =>
                           REGISTERS_3_30_port, B2 => n187_port, ZN => n1210);
   U1202 : AOI22_X1 port map( A1 => REGISTERS_4_30_port, A2 => n238, B1 => 
                           REGISTERS_6_30_port, B2 => n221, ZN => n1209);
   U1203 : AOI22_X1 port map( A1 => REGISTERS_0_30_port, A2 => n272, B1 => 
                           REGISTERS_2_30_port, B2 => n255, ZN => n1208);
   U1204 : NAND4_X1 port map( A1 => n1211, A2 => n1210, A3 => n1209, A4 => 
                           n1208, ZN => n1217);
   U1205 : AOI22_X1 port map( A1 => REGISTERS_13_30_port, A2 => n170_port, B1 
                           => REGISTERS_15_30_port, B2 => n153, ZN => n1215);
   U1206 : AOI22_X1 port map( A1 => REGISTERS_9_30_port, A2 => n204_port, B1 =>
                           REGISTERS_11_30_port, B2 => n187_port, ZN => n1214);
   U1207 : AOI22_X1 port map( A1 => REGISTERS_12_30_port, A2 => n238, B1 => 
                           REGISTERS_14_30_port, B2 => n221, ZN => n1213);
   U1208 : AOI22_X1 port map( A1 => REGISTERS_8_30_port, A2 => n272, B1 => 
                           REGISTERS_10_30_port, B2 => n255, ZN => n1212);
   U1209 : NAND4_X1 port map( A1 => n1215, A2 => n1214, A3 => n1213, A4 => 
                           n1212, ZN => n1216);
   U1210 : AOI22_X1 port map( A1 => n1217, A2 => n1240, B1 => n1216, B2 => 
                           n1238, ZN => n1218);
   U1211 : OAI221_X1 port map( B1 => n1244, B2 => n1220, C1 => n1242, C2 => 
                           n1219, A => n1218, ZN => N157);
   U1212 : AOI22_X1 port map( A1 => REGISTERS_21_31_port, A2 => n170_port, B1 
                           => REGISTERS_23_31_port, B2 => n153, ZN => n1224);
   U1213 : AOI22_X1 port map( A1 => REGISTERS_17_31_port, A2 => n204_port, B1 
                           => REGISTERS_19_31_port, B2 => n187_port, ZN => 
                           n1223);
   U1214 : AOI22_X1 port map( A1 => REGISTERS_20_31_port, A2 => n238, B1 => 
                           REGISTERS_22_31_port, B2 => n221, ZN => n1222);
   U1215 : AOI22_X1 port map( A1 => REGISTERS_16_31_port, A2 => n272, B1 => 
                           REGISTERS_18_31_port, B2 => n255, ZN => n1221);
   U1216 : AND4_X1 port map( A1 => n1224, A2 => n1223, A3 => n1222, A4 => n1221
                           , ZN => n1245);
   U1217 : AOI22_X1 port map( A1 => REGISTERS_29_31_port, A2 => n170_port, B1 
                           => REGISTERS_31_31_port, B2 => n153, ZN => n1228);
   U1218 : AOI22_X1 port map( A1 => REGISTERS_25_31_port, A2 => n204_port, B1 
                           => REGISTERS_27_31_port, B2 => n187_port, ZN => 
                           n1227);
   U1219 : AOI22_X1 port map( A1 => REGISTERS_28_31_port, A2 => n238, B1 => 
                           REGISTERS_30_31_port, B2 => n221, ZN => n1226);
   U1220 : AOI22_X1 port map( A1 => REGISTERS_24_31_port, A2 => n272, B1 => 
                           REGISTERS_26_31_port, B2 => n255, ZN => n1225);
   U1221 : AND4_X1 port map( A1 => n1228, A2 => n1227, A3 => n1226, A4 => n1225
                           , ZN => n1243);
   U1222 : AOI22_X1 port map( A1 => REGISTERS_5_31_port, A2 => n170_port, B1 =>
                           REGISTERS_7_31_port, B2 => n153, ZN => n1232);
   U1223 : AOI22_X1 port map( A1 => REGISTERS_1_31_port, A2 => n204_port, B1 =>
                           REGISTERS_3_31_port, B2 => n187_port, ZN => n1231);
   U1224 : AOI22_X1 port map( A1 => REGISTERS_4_31_port, A2 => n238, B1 => 
                           REGISTERS_6_31_port, B2 => n221, ZN => n1230);
   U1225 : AOI22_X1 port map( A1 => REGISTERS_0_31_port, A2 => n272, B1 => 
                           REGISTERS_2_31_port, B2 => n255, ZN => n1229);
   U1226 : NAND4_X1 port map( A1 => n1232, A2 => n1231, A3 => n1230, A4 => 
                           n1229, ZN => n1239);
   U1227 : AOI22_X1 port map( A1 => REGISTERS_13_31_port, A2 => n170_port, B1 
                           => REGISTERS_15_31_port, B2 => n153, ZN => n1236);
   U1228 : AOI22_X1 port map( A1 => REGISTERS_9_31_port, A2 => n204_port, B1 =>
                           REGISTERS_11_31_port, B2 => n187_port, ZN => n1235);
   U1229 : AOI22_X1 port map( A1 => REGISTERS_12_31_port, A2 => n238, B1 => 
                           REGISTERS_14_31_port, B2 => n221, ZN => n1234);
   U1230 : AOI22_X1 port map( A1 => REGISTERS_8_31_port, A2 => n272, B1 => 
                           REGISTERS_10_31_port, B2 => n255, ZN => n1233);
   U1231 : NAND4_X1 port map( A1 => n1236, A2 => n1235, A3 => n1234, A4 => 
                           n1233, ZN => n1237);
   U1232 : AOI22_X1 port map( A1 => n1240, A2 => n1239, B1 => n1238, B2 => 
                           n1237, ZN => n1241);
   U1233 : OAI221_X1 port map( B1 => n1245, B2 => n1244, C1 => n1243, C2 => 
                           n1242, A => n1241, ZN => N156);
   U1234 : NOR2_X1 port map( A1 => n3084, A2 => ADD_RD2(1), ZN => n1250);
   U1235 : NOR2_X1 port map( A1 => n3084, A2 => n3083, ZN => n1251);
   U1236 : AOI22_X1 port map( A1 => REGISTERS_21_0_port, A2 => n296, B1 => 
                           REGISTERS_23_0_port, B2 => n279, ZN => n1257);
   U1237 : NOR2_X1 port map( A1 => ADD_RD2(1), A2 => ADD_RD2(2), ZN => n1252);
   U1238 : NOR2_X1 port map( A1 => n3083, A2 => ADD_RD2(2), ZN => n1253);
   U1239 : AOI22_X1 port map( A1 => REGISTERS_17_0_port, A2 => n330, B1 => 
                           REGISTERS_19_0_port, B2 => n313, ZN => n1256);
   U1240 : AOI22_X1 port map( A1 => REGISTERS_20_0_port, A2 => n364, B1 => 
                           REGISTERS_22_0_port, B2 => n347, ZN => n1255);
   U1241 : AOI22_X1 port map( A1 => REGISTERS_16_0_port, A2 => n398, B1 => 
                           REGISTERS_18_0_port, B2 => n381, ZN => n1254);
   U1242 : AND4_X1 port map( A1 => n1257, A2 => n1256, A3 => n1255, A4 => n1254
                           , ZN => n1274);
   U1243 : AOI22_X1 port map( A1 => REGISTERS_29_0_port, A2 => n296, B1 => 
                           REGISTERS_31_0_port, B2 => n279, ZN => n1261);
   U1244 : AOI22_X1 port map( A1 => REGISTERS_25_0_port, A2 => n330, B1 => 
                           REGISTERS_27_0_port, B2 => n313, ZN => n1260);
   U1245 : AOI22_X1 port map( A1 => REGISTERS_28_0_port, A2 => n364, B1 => 
                           REGISTERS_30_0_port, B2 => n347, ZN => n1259);
   U1246 : AOI22_X1 port map( A1 => REGISTERS_24_0_port, A2 => n398, B1 => 
                           REGISTERS_26_0_port, B2 => n381, ZN => n1258);
   U1247 : AND4_X1 port map( A1 => n1261, A2 => n1260, A3 => n1259, A4 => n1258
                           , ZN => n1273);
   U1248 : AOI22_X1 port map( A1 => REGISTERS_5_0_port, A2 => n296, B1 => 
                           REGISTERS_7_0_port, B2 => n279, ZN => n1265);
   U1249 : AOI22_X1 port map( A1 => REGISTERS_1_0_port, A2 => n330, B1 => 
                           REGISTERS_3_0_port, B2 => n313, ZN => n1264);
   U1250 : AOI22_X1 port map( A1 => REGISTERS_4_0_port, A2 => n364, B1 => 
                           REGISTERS_6_0_port, B2 => n347, ZN => n1263);
   U1251 : AOI22_X1 port map( A1 => REGISTERS_0_0_port, A2 => n398, B1 => 
                           REGISTERS_2_0_port, B2 => n381, ZN => n1262);
   U1252 : NAND4_X1 port map( A1 => n1265, A2 => n1264, A3 => n1263, A4 => 
                           n1262, ZN => n1271);
   U1253 : AOI22_X1 port map( A1 => REGISTERS_13_0_port, A2 => n296, B1 => 
                           REGISTERS_15_0_port, B2 => n279, ZN => n1269);
   U1254 : AOI22_X1 port map( A1 => REGISTERS_9_0_port, A2 => n330, B1 => 
                           REGISTERS_11_0_port, B2 => n313, ZN => n1268);
   U1255 : AOI22_X1 port map( A1 => REGISTERS_12_0_port, A2 => n364, B1 => 
                           REGISTERS_14_0_port, B2 => n347, ZN => n1267);
   U1256 : AOI22_X1 port map( A1 => REGISTERS_8_0_port, A2 => n398, B1 => 
                           REGISTERS_10_0_port, B2 => n381, ZN => n1266);
   U1257 : NAND4_X1 port map( A1 => n1269, A2 => n1268, A3 => n1267, A4 => 
                           n1266, ZN => n1270);
   U1258 : AOI22_X1 port map( A1 => n1271, A2 => n3076, B1 => n1270, B2 => 
                           n3074, ZN => n1272);
   U1259 : OAI221_X1 port map( B1 => n3080, B2 => n1274, C1 => n3078, C2 => 
                           n1273, A => n1272, ZN => N220);
   U1260 : AOI22_X1 port map( A1 => REGISTERS_21_1_port, A2 => n296, B1 => 
                           REGISTERS_23_1_port, B2 => n279, ZN => n1278);
   U1261 : AOI22_X1 port map( A1 => REGISTERS_17_1_port, A2 => n330, B1 => 
                           REGISTERS_19_1_port, B2 => n313, ZN => n1277);
   U1262 : AOI22_X1 port map( A1 => REGISTERS_20_1_port, A2 => n364, B1 => 
                           REGISTERS_22_1_port, B2 => n347, ZN => n1276);
   U1263 : AOI22_X1 port map( A1 => REGISTERS_16_1_port, A2 => n398, B1 => 
                           REGISTERS_18_1_port, B2 => n381, ZN => n1275);
   U1264 : AND4_X1 port map( A1 => n1278, A2 => n1277, A3 => n1276, A4 => n1275
                           , ZN => n1295);
   U1265 : AOI22_X1 port map( A1 => REGISTERS_29_1_port, A2 => n296, B1 => 
                           REGISTERS_31_1_port, B2 => n279, ZN => n1282);
   U1266 : AOI22_X1 port map( A1 => REGISTERS_25_1_port, A2 => n330, B1 => 
                           REGISTERS_27_1_port, B2 => n313, ZN => n1281);
   U1267 : AOI22_X1 port map( A1 => REGISTERS_28_1_port, A2 => n364, B1 => 
                           REGISTERS_30_1_port, B2 => n347, ZN => n1280);
   U1268 : AOI22_X1 port map( A1 => REGISTERS_24_1_port, A2 => n398, B1 => 
                           REGISTERS_26_1_port, B2 => n381, ZN => n1279);
   U1269 : AND4_X1 port map( A1 => n1282, A2 => n1281, A3 => n1280, A4 => n1279
                           , ZN => n1294);
   U1270 : AOI22_X1 port map( A1 => REGISTERS_5_1_port, A2 => n296, B1 => 
                           REGISTERS_7_1_port, B2 => n279, ZN => n1286);
   U1271 : AOI22_X1 port map( A1 => REGISTERS_1_1_port, A2 => n330, B1 => 
                           REGISTERS_3_1_port, B2 => n313, ZN => n1285);
   U1272 : AOI22_X1 port map( A1 => REGISTERS_4_1_port, A2 => n364, B1 => 
                           REGISTERS_6_1_port, B2 => n347, ZN => n1284);
   U1273 : AOI22_X1 port map( A1 => REGISTERS_0_1_port, A2 => n398, B1 => 
                           REGISTERS_2_1_port, B2 => n381, ZN => n1283);
   U1274 : NAND4_X1 port map( A1 => n1286, A2 => n1285, A3 => n1284, A4 => 
                           n1283, ZN => n1292);
   U1275 : AOI22_X1 port map( A1 => REGISTERS_13_1_port, A2 => n296, B1 => 
                           REGISTERS_15_1_port, B2 => n279, ZN => n1290);
   U1276 : AOI22_X1 port map( A1 => REGISTERS_9_1_port, A2 => n330, B1 => 
                           REGISTERS_11_1_port, B2 => n313, ZN => n1289);
   U1277 : AOI22_X1 port map( A1 => REGISTERS_12_1_port, A2 => n364, B1 => 
                           REGISTERS_14_1_port, B2 => n347, ZN => n1288);
   U1278 : AOI22_X1 port map( A1 => REGISTERS_8_1_port, A2 => n398, B1 => 
                           REGISTERS_10_1_port, B2 => n381, ZN => n1287);
   U1279 : NAND4_X1 port map( A1 => n1290, A2 => n1289, A3 => n1288, A4 => 
                           n1287, ZN => n1291);
   U1280 : AOI22_X1 port map( A1 => n1292, A2 => n3076, B1 => n1291, B2 => 
                           n3074, ZN => n1293);
   U1281 : OAI221_X1 port map( B1 => n3080, B2 => n1295, C1 => n3078, C2 => 
                           n1294, A => n1293, ZN => N219);
   U1282 : AOI22_X1 port map( A1 => REGISTERS_21_2_port, A2 => n296, B1 => 
                           REGISTERS_23_2_port, B2 => n279, ZN => n1299);
   U1283 : AOI22_X1 port map( A1 => REGISTERS_17_2_port, A2 => n330, B1 => 
                           REGISTERS_19_2_port, B2 => n313, ZN => n1298);
   U1284 : AOI22_X1 port map( A1 => REGISTERS_20_2_port, A2 => n364, B1 => 
                           REGISTERS_22_2_port, B2 => n347, ZN => n1297);
   U1285 : AOI22_X1 port map( A1 => REGISTERS_16_2_port, A2 => n398, B1 => 
                           REGISTERS_18_2_port, B2 => n381, ZN => n1296);
   U1286 : AND4_X1 port map( A1 => n1299, A2 => n1298, A3 => n1297, A4 => n1296
                           , ZN => n1316);
   U1287 : AOI22_X1 port map( A1 => REGISTERS_29_2_port, A2 => n296, B1 => 
                           REGISTERS_31_2_port, B2 => n279, ZN => n1303);
   U1288 : AOI22_X1 port map( A1 => REGISTERS_25_2_port, A2 => n330, B1 => 
                           REGISTERS_27_2_port, B2 => n313, ZN => n1302);
   U1289 : AOI22_X1 port map( A1 => REGISTERS_28_2_port, A2 => n364, B1 => 
                           REGISTERS_30_2_port, B2 => n347, ZN => n1301);
   U1290 : AOI22_X1 port map( A1 => REGISTERS_24_2_port, A2 => n398, B1 => 
                           REGISTERS_26_2_port, B2 => n381, ZN => n1300);
   U1291 : AND4_X1 port map( A1 => n1303, A2 => n1302, A3 => n1301, A4 => n1300
                           , ZN => n1315);
   U1292 : AOI22_X1 port map( A1 => REGISTERS_5_2_port, A2 => n296, B1 => 
                           REGISTERS_7_2_port, B2 => n279, ZN => n1307);
   U1293 : AOI22_X1 port map( A1 => REGISTERS_1_2_port, A2 => n330, B1 => 
                           REGISTERS_3_2_port, B2 => n313, ZN => n1306);
   U1294 : AOI22_X1 port map( A1 => REGISTERS_4_2_port, A2 => n364, B1 => 
                           REGISTERS_6_2_port, B2 => n347, ZN => n1305);
   U1295 : AOI22_X1 port map( A1 => REGISTERS_0_2_port, A2 => n398, B1 => 
                           REGISTERS_2_2_port, B2 => n381, ZN => n1304);
   U1296 : NAND4_X1 port map( A1 => n1307, A2 => n1306, A3 => n1305, A4 => 
                           n1304, ZN => n1313);
   U1297 : AOI22_X1 port map( A1 => REGISTERS_13_2_port, A2 => n296, B1 => 
                           REGISTERS_15_2_port, B2 => n279, ZN => n1311);
   U1298 : AOI22_X1 port map( A1 => REGISTERS_9_2_port, A2 => n330, B1 => 
                           REGISTERS_11_2_port, B2 => n313, ZN => n1310);
   U1299 : AOI22_X1 port map( A1 => REGISTERS_12_2_port, A2 => n364, B1 => 
                           REGISTERS_14_2_port, B2 => n347, ZN => n1309);
   U1300 : AOI22_X1 port map( A1 => REGISTERS_8_2_port, A2 => n398, B1 => 
                           REGISTERS_10_2_port, B2 => n381, ZN => n1308);
   U1301 : NAND4_X1 port map( A1 => n1311, A2 => n1310, A3 => n1309, A4 => 
                           n1308, ZN => n1312);
   U1302 : AOI22_X1 port map( A1 => n1313, A2 => n3076, B1 => n1312, B2 => 
                           n3074, ZN => n1314);
   U1303 : OAI221_X1 port map( B1 => n3080, B2 => n1316, C1 => n3078, C2 => 
                           n1315, A => n1314, ZN => N218);
   U1304 : AOI22_X1 port map( A1 => REGISTERS_21_3_port, A2 => n297, B1 => 
                           REGISTERS_23_3_port, B2 => n280, ZN => n1320);
   U1305 : AOI22_X1 port map( A1 => REGISTERS_17_3_port, A2 => n331, B1 => 
                           REGISTERS_19_3_port, B2 => n314, ZN => n1319);
   U1306 : AOI22_X1 port map( A1 => REGISTERS_20_3_port, A2 => n365, B1 => 
                           REGISTERS_22_3_port, B2 => n348, ZN => n1318);
   U1307 : AOI22_X1 port map( A1 => REGISTERS_16_3_port, A2 => n399, B1 => 
                           REGISTERS_18_3_port, B2 => n382, ZN => n1317);
   U1308 : AND4_X1 port map( A1 => n1320, A2 => n1319, A3 => n1318, A4 => n1317
                           , ZN => n1337);
   U1309 : AOI22_X1 port map( A1 => REGISTERS_29_3_port, A2 => n297, B1 => 
                           REGISTERS_31_3_port, B2 => n280, ZN => n1324);
   U1310 : AOI22_X1 port map( A1 => REGISTERS_25_3_port, A2 => n331, B1 => 
                           REGISTERS_27_3_port, B2 => n314, ZN => n1323);
   U1311 : AOI22_X1 port map( A1 => REGISTERS_28_3_port, A2 => n365, B1 => 
                           REGISTERS_30_3_port, B2 => n348, ZN => n1322);
   U1312 : AOI22_X1 port map( A1 => REGISTERS_24_3_port, A2 => n399, B1 => 
                           REGISTERS_26_3_port, B2 => n382, ZN => n1321);
   U1313 : AND4_X1 port map( A1 => n1324, A2 => n1323, A3 => n1322, A4 => n1321
                           , ZN => n1336);
   U1314 : AOI22_X1 port map( A1 => REGISTERS_5_3_port, A2 => n297, B1 => 
                           REGISTERS_7_3_port, B2 => n280, ZN => n1328);
   U1315 : AOI22_X1 port map( A1 => REGISTERS_1_3_port, A2 => n331, B1 => 
                           REGISTERS_3_3_port, B2 => n314, ZN => n1327);
   U1316 : AOI22_X1 port map( A1 => REGISTERS_4_3_port, A2 => n365, B1 => 
                           REGISTERS_6_3_port, B2 => n348, ZN => n1326);
   U1317 : AOI22_X1 port map( A1 => REGISTERS_0_3_port, A2 => n399, B1 => 
                           REGISTERS_2_3_port, B2 => n382, ZN => n1325);
   U1318 : NAND4_X1 port map( A1 => n1328, A2 => n1327, A3 => n1326, A4 => 
                           n1325, ZN => n1334);
   U1319 : AOI22_X1 port map( A1 => REGISTERS_13_3_port, A2 => n297, B1 => 
                           REGISTERS_15_3_port, B2 => n280, ZN => n1332);
   U1320 : AOI22_X1 port map( A1 => REGISTERS_9_3_port, A2 => n331, B1 => 
                           REGISTERS_11_3_port, B2 => n314, ZN => n1331);
   U1321 : AOI22_X1 port map( A1 => REGISTERS_12_3_port, A2 => n365, B1 => 
                           REGISTERS_14_3_port, B2 => n348, ZN => n1330);
   U1322 : AOI22_X1 port map( A1 => REGISTERS_8_3_port, A2 => n399, B1 => 
                           REGISTERS_10_3_port, B2 => n382, ZN => n1329);
   U1323 : NAND4_X1 port map( A1 => n1332, A2 => n1331, A3 => n1330, A4 => 
                           n1329, ZN => n1333);
   U1324 : AOI22_X1 port map( A1 => n1334, A2 => n3076, B1 => n1333, B2 => 
                           n3074, ZN => n1335);
   U1325 : OAI221_X1 port map( B1 => n3080, B2 => n1337, C1 => n3078, C2 => 
                           n1336, A => n1335, ZN => N217);
   U1326 : AOI22_X1 port map( A1 => REGISTERS_21_4_port, A2 => n297, B1 => 
                           REGISTERS_23_4_port, B2 => n280, ZN => n1341);
   U1327 : AOI22_X1 port map( A1 => REGISTERS_17_4_port, A2 => n331, B1 => 
                           REGISTERS_19_4_port, B2 => n314, ZN => n1340);
   U1328 : AOI22_X1 port map( A1 => REGISTERS_20_4_port, A2 => n365, B1 => 
                           REGISTERS_22_4_port, B2 => n348, ZN => n1339);
   U1329 : AOI22_X1 port map( A1 => REGISTERS_16_4_port, A2 => n399, B1 => 
                           REGISTERS_18_4_port, B2 => n382, ZN => n1338);
   U1330 : AND4_X1 port map( A1 => n1341, A2 => n1340, A3 => n1339, A4 => n1338
                           , ZN => n1358);
   U1331 : AOI22_X1 port map( A1 => REGISTERS_29_4_port, A2 => n297, B1 => 
                           REGISTERS_31_4_port, B2 => n280, ZN => n1345);
   U1332 : AOI22_X1 port map( A1 => REGISTERS_25_4_port, A2 => n331, B1 => 
                           REGISTERS_27_4_port, B2 => n314, ZN => n1344);
   U1333 : AOI22_X1 port map( A1 => REGISTERS_28_4_port, A2 => n365, B1 => 
                           REGISTERS_30_4_port, B2 => n348, ZN => n1343);
   U1334 : AOI22_X1 port map( A1 => REGISTERS_24_4_port, A2 => n399, B1 => 
                           REGISTERS_26_4_port, B2 => n382, ZN => n1342);
   U1335 : AND4_X1 port map( A1 => n1345, A2 => n1344, A3 => n1343, A4 => n1342
                           , ZN => n1357);
   U1336 : AOI22_X1 port map( A1 => REGISTERS_5_4_port, A2 => n297, B1 => 
                           REGISTERS_7_4_port, B2 => n280, ZN => n1349);
   U1337 : AOI22_X1 port map( A1 => REGISTERS_1_4_port, A2 => n331, B1 => 
                           REGISTERS_3_4_port, B2 => n314, ZN => n1348);
   U1338 : AOI22_X1 port map( A1 => REGISTERS_4_4_port, A2 => n365, B1 => 
                           REGISTERS_6_4_port, B2 => n348, ZN => n1347);
   U1339 : AOI22_X1 port map( A1 => REGISTERS_0_4_port, A2 => n399, B1 => 
                           REGISTERS_2_4_port, B2 => n382, ZN => n1346);
   U1340 : NAND4_X1 port map( A1 => n1349, A2 => n1348, A3 => n1347, A4 => 
                           n1346, ZN => n1355);
   U1341 : AOI22_X1 port map( A1 => REGISTERS_13_4_port, A2 => n297, B1 => 
                           REGISTERS_15_4_port, B2 => n280, ZN => n1353);
   U1342 : AOI22_X1 port map( A1 => REGISTERS_9_4_port, A2 => n331, B1 => 
                           REGISTERS_11_4_port, B2 => n314, ZN => n1352);
   U1343 : AOI22_X1 port map( A1 => REGISTERS_12_4_port, A2 => n365, B1 => 
                           REGISTERS_14_4_port, B2 => n348, ZN => n1351);
   U1344 : AOI22_X1 port map( A1 => REGISTERS_8_4_port, A2 => n399, B1 => 
                           REGISTERS_10_4_port, B2 => n382, ZN => n1350);
   U1345 : NAND4_X1 port map( A1 => n1353, A2 => n1352, A3 => n1351, A4 => 
                           n1350, ZN => n1354);
   U1346 : AOI22_X1 port map( A1 => n1355, A2 => n3076, B1 => n1354, B2 => 
                           n3074, ZN => n1356);
   U1347 : OAI221_X1 port map( B1 => n3080, B2 => n1358, C1 => n3078, C2 => 
                           n1357, A => n1356, ZN => N216);
   U1348 : AOI22_X1 port map( A1 => REGISTERS_21_5_port, A2 => n297, B1 => 
                           REGISTERS_23_5_port, B2 => n280, ZN => n1362);
   U1349 : AOI22_X1 port map( A1 => REGISTERS_17_5_port, A2 => n331, B1 => 
                           REGISTERS_19_5_port, B2 => n314, ZN => n1361);
   U1350 : AOI22_X1 port map( A1 => REGISTERS_20_5_port, A2 => n365, B1 => 
                           REGISTERS_22_5_port, B2 => n348, ZN => n1360);
   U1351 : AOI22_X1 port map( A1 => REGISTERS_16_5_port, A2 => n399, B1 => 
                           REGISTERS_18_5_port, B2 => n382, ZN => n1359);
   U1352 : AND4_X1 port map( A1 => n1362, A2 => n1361, A3 => n1360, A4 => n1359
                           , ZN => n1379);
   U1353 : AOI22_X1 port map( A1 => REGISTERS_29_5_port, A2 => n297, B1 => 
                           REGISTERS_31_5_port, B2 => n280, ZN => n1366);
   U1354 : AOI22_X1 port map( A1 => REGISTERS_25_5_port, A2 => n331, B1 => 
                           REGISTERS_27_5_port, B2 => n314, ZN => n1365);
   U1355 : AOI22_X1 port map( A1 => REGISTERS_28_5_port, A2 => n365, B1 => 
                           REGISTERS_30_5_port, B2 => n348, ZN => n1364);
   U1356 : AOI22_X1 port map( A1 => REGISTERS_24_5_port, A2 => n399, B1 => 
                           REGISTERS_26_5_port, B2 => n382, ZN => n1363);
   U1357 : AND4_X1 port map( A1 => n1366, A2 => n1365, A3 => n1364, A4 => n1363
                           , ZN => n1378);
   U1358 : AOI22_X1 port map( A1 => REGISTERS_5_5_port, A2 => n297, B1 => 
                           REGISTERS_7_5_port, B2 => n280, ZN => n1370);
   U1359 : AOI22_X1 port map( A1 => REGISTERS_1_5_port, A2 => n331, B1 => 
                           REGISTERS_3_5_port, B2 => n314, ZN => n1369);
   U1360 : AOI22_X1 port map( A1 => REGISTERS_4_5_port, A2 => n365, B1 => 
                           REGISTERS_6_5_port, B2 => n348, ZN => n1368);
   U1361 : AOI22_X1 port map( A1 => REGISTERS_0_5_port, A2 => n399, B1 => 
                           REGISTERS_2_5_port, B2 => n382, ZN => n1367);
   U1362 : NAND4_X1 port map( A1 => n1370, A2 => n1369, A3 => n1368, A4 => 
                           n1367, ZN => n1376);
   U1363 : AOI22_X1 port map( A1 => REGISTERS_13_5_port, A2 => n297, B1 => 
                           REGISTERS_15_5_port, B2 => n280, ZN => n1374);
   U1364 : AOI22_X1 port map( A1 => REGISTERS_9_5_port, A2 => n331, B1 => 
                           REGISTERS_11_5_port, B2 => n314, ZN => n1373);
   U1365 : AOI22_X1 port map( A1 => REGISTERS_12_5_port, A2 => n365, B1 => 
                           REGISTERS_14_5_port, B2 => n348, ZN => n1372);
   U1366 : AOI22_X1 port map( A1 => REGISTERS_8_5_port, A2 => n399, B1 => 
                           REGISTERS_10_5_port, B2 => n382, ZN => n1371);
   U1367 : NAND4_X1 port map( A1 => n1374, A2 => n1373, A3 => n1372, A4 => 
                           n1371, ZN => n1375);
   U1368 : AOI22_X1 port map( A1 => n1376, A2 => n3076, B1 => n1375, B2 => 
                           n3074, ZN => n1377);
   U1369 : OAI221_X1 port map( B1 => n3080, B2 => n1379, C1 => n3078, C2 => 
                           n1378, A => n1377, ZN => N215);
   U1370 : AOI22_X1 port map( A1 => REGISTERS_21_6_port, A2 => n298, B1 => 
                           REGISTERS_23_6_port, B2 => n281, ZN => n1383);
   U1371 : AOI22_X1 port map( A1 => REGISTERS_17_6_port, A2 => n332, B1 => 
                           REGISTERS_19_6_port, B2 => n315, ZN => n1382);
   U1372 : AOI22_X1 port map( A1 => REGISTERS_20_6_port, A2 => n366, B1 => 
                           REGISTERS_22_6_port, B2 => n349, ZN => n1381);
   U1373 : AOI22_X1 port map( A1 => REGISTERS_16_6_port, A2 => n400, B1 => 
                           REGISTERS_18_6_port, B2 => n383, ZN => n1380);
   U1374 : AND4_X1 port map( A1 => n1383, A2 => n1382, A3 => n1381, A4 => n1380
                           , ZN => n1402);
   U1375 : AOI22_X1 port map( A1 => REGISTERS_29_6_port, A2 => n298, B1 => 
                           REGISTERS_31_6_port, B2 => n281, ZN => n1387);
   U1376 : AOI22_X1 port map( A1 => REGISTERS_25_6_port, A2 => n332, B1 => 
                           REGISTERS_27_6_port, B2 => n315, ZN => n1386);
   U1377 : AOI22_X1 port map( A1 => REGISTERS_28_6_port, A2 => n366, B1 => 
                           REGISTERS_30_6_port, B2 => n349, ZN => n1385);
   U1378 : AOI22_X1 port map( A1 => REGISTERS_24_6_port, A2 => n400, B1 => 
                           REGISTERS_26_6_port, B2 => n383, ZN => n1384);
   U1379 : AND4_X1 port map( A1 => n1387, A2 => n1386, A3 => n1385, A4 => n1384
                           , ZN => n1400);
   U1380 : AOI22_X1 port map( A1 => REGISTERS_5_6_port, A2 => n298, B1 => 
                           REGISTERS_7_6_port, B2 => n281, ZN => n1391);
   U1381 : AOI22_X1 port map( A1 => REGISTERS_1_6_port, A2 => n332, B1 => 
                           REGISTERS_3_6_port, B2 => n315, ZN => n1390);
   U1382 : AOI22_X1 port map( A1 => REGISTERS_4_6_port, A2 => n366, B1 => 
                           REGISTERS_6_6_port, B2 => n349, ZN => n1389);
   U1383 : AOI22_X1 port map( A1 => REGISTERS_0_6_port, A2 => n400, B1 => 
                           REGISTERS_2_6_port, B2 => n383, ZN => n1388);
   U1384 : NAND4_X1 port map( A1 => n1391, A2 => n1390, A3 => n1389, A4 => 
                           n1388, ZN => n1397);
   U1385 : AOI22_X1 port map( A1 => REGISTERS_13_6_port, A2 => n298, B1 => 
                           REGISTERS_15_6_port, B2 => n281, ZN => n1395);
   U1386 : AOI22_X1 port map( A1 => REGISTERS_9_6_port, A2 => n332, B1 => 
                           REGISTERS_11_6_port, B2 => n315, ZN => n1394);
   U1387 : AOI22_X1 port map( A1 => REGISTERS_12_6_port, A2 => n366, B1 => 
                           REGISTERS_14_6_port, B2 => n349, ZN => n1393);
   U1388 : AOI22_X1 port map( A1 => REGISTERS_8_6_port, A2 => n400, B1 => 
                           REGISTERS_10_6_port, B2 => n383, ZN => n1392);
   U1389 : NAND4_X1 port map( A1 => n1395, A2 => n1394, A3 => n1393, A4 => 
                           n1392, ZN => n1396);
   U1390 : AOI22_X1 port map( A1 => n1397, A2 => n3076, B1 => n1396, B2 => 
                           n3074, ZN => n1398);
   U1391 : OAI221_X1 port map( B1 => n3080, B2 => n1402, C1 => n3078, C2 => 
                           n1400, A => n1398, ZN => N214);
   U1392 : AOI22_X1 port map( A1 => REGISTERS_21_7_port, A2 => n298, B1 => 
                           REGISTERS_23_7_port, B2 => n281, ZN => n1410);
   U1393 : AOI22_X1 port map( A1 => REGISTERS_17_7_port, A2 => n332, B1 => 
                           REGISTERS_19_7_port, B2 => n315, ZN => n1408);
   U1394 : AOI22_X1 port map( A1 => REGISTERS_20_7_port, A2 => n366, B1 => 
                           REGISTERS_22_7_port, B2 => n349, ZN => n1406);
   U1395 : AOI22_X1 port map( A1 => REGISTERS_16_7_port, A2 => n400, B1 => 
                           REGISTERS_18_7_port, B2 => n383, ZN => n1404);
   U1396 : AND4_X1 port map( A1 => n1410, A2 => n1408, A3 => n1406, A4 => n1404
                           , ZN => n1444);
   U1397 : AOI22_X1 port map( A1 => REGISTERS_29_7_port, A2 => n298, B1 => 
                           REGISTERS_31_7_port, B2 => n281, ZN => n1418);
   U1398 : AOI22_X1 port map( A1 => REGISTERS_25_7_port, A2 => n332, B1 => 
                           REGISTERS_27_7_port, B2 => n315, ZN => n1416);
   U1399 : AOI22_X1 port map( A1 => REGISTERS_28_7_port, A2 => n366, B1 => 
                           REGISTERS_30_7_port, B2 => n349, ZN => n1414);
   U1400 : AOI22_X1 port map( A1 => REGISTERS_24_7_port, A2 => n400, B1 => 
                           REGISTERS_26_7_port, B2 => n383, ZN => n1412);
   U1401 : AND4_X1 port map( A1 => n1418, A2 => n1416, A3 => n1414, A4 => n1412
                           , ZN => n1442);
   U1402 : AOI22_X1 port map( A1 => REGISTERS_5_7_port, A2 => n298, B1 => 
                           REGISTERS_7_7_port, B2 => n281, ZN => n1426);
   U1403 : AOI22_X1 port map( A1 => REGISTERS_1_7_port, A2 => n332, B1 => 
                           REGISTERS_3_7_port, B2 => n315, ZN => n1424);
   U1404 : AOI22_X1 port map( A1 => REGISTERS_4_7_port, A2 => n366, B1 => 
                           REGISTERS_6_7_port, B2 => n349, ZN => n1422);
   U1405 : AOI22_X1 port map( A1 => REGISTERS_0_7_port, A2 => n400, B1 => 
                           REGISTERS_2_7_port, B2 => n383, ZN => n1420);
   U1406 : NAND4_X1 port map( A1 => n1426, A2 => n1424, A3 => n1422, A4 => 
                           n1420, ZN => n1438);
   U1407 : AOI22_X1 port map( A1 => REGISTERS_13_7_port, A2 => n298, B1 => 
                           REGISTERS_15_7_port, B2 => n281, ZN => n1434);
   U1408 : AOI22_X1 port map( A1 => REGISTERS_9_7_port, A2 => n332, B1 => 
                           REGISTERS_11_7_port, B2 => n315, ZN => n1432);
   U1409 : AOI22_X1 port map( A1 => REGISTERS_12_7_port, A2 => n366, B1 => 
                           REGISTERS_14_7_port, B2 => n349, ZN => n1430);
   U1410 : AOI22_X1 port map( A1 => REGISTERS_8_7_port, A2 => n400, B1 => 
                           REGISTERS_10_7_port, B2 => n383, ZN => n1428);
   U1411 : NAND4_X1 port map( A1 => n1434, A2 => n1432, A3 => n1430, A4 => 
                           n1428, ZN => n1436);
   U1412 : AOI22_X1 port map( A1 => n1438, A2 => n3076, B1 => n1436, B2 => 
                           n3074, ZN => n1440);
   U1413 : OAI221_X1 port map( B1 => n3080, B2 => n1444, C1 => n3078, C2 => 
                           n1442, A => n1440, ZN => N213);
   U1414 : AOI22_X1 port map( A1 => REGISTERS_21_8_port, A2 => n298, B1 => 
                           REGISTERS_23_8_port, B2 => n281, ZN => n1452);
   U1415 : AOI22_X1 port map( A1 => REGISTERS_17_8_port, A2 => n332, B1 => 
                           REGISTERS_19_8_port, B2 => n315, ZN => n1450);
   U1416 : AOI22_X1 port map( A1 => REGISTERS_20_8_port, A2 => n366, B1 => 
                           REGISTERS_22_8_port, B2 => n349, ZN => n1448);
   U1417 : AOI22_X1 port map( A1 => REGISTERS_16_8_port, A2 => n400, B1 => 
                           REGISTERS_18_8_port, B2 => n383, ZN => n1446);
   U1418 : AND4_X1 port map( A1 => n1452, A2 => n1450, A3 => n1448, A4 => n1446
                           , ZN => n1506);
   U1419 : AOI22_X1 port map( A1 => REGISTERS_29_8_port, A2 => n298, B1 => 
                           REGISTERS_31_8_port, B2 => n281, ZN => n1460);
   U1420 : AOI22_X1 port map( A1 => REGISTERS_25_8_port, A2 => n332, B1 => 
                           REGISTERS_27_8_port, B2 => n315, ZN => n1458);
   U1421 : AOI22_X1 port map( A1 => REGISTERS_28_8_port, A2 => n366, B1 => 
                           REGISTERS_30_8_port, B2 => n349, ZN => n1456);
   U1422 : AOI22_X1 port map( A1 => REGISTERS_24_8_port, A2 => n400, B1 => 
                           REGISTERS_26_8_port, B2 => n383, ZN => n1454);
   U1423 : AND4_X1 port map( A1 => n1460, A2 => n1458, A3 => n1456, A4 => n1454
                           , ZN => n1505);
   U1424 : AOI22_X1 port map( A1 => REGISTERS_5_8_port, A2 => n298, B1 => 
                           REGISTERS_7_8_port, B2 => n281, ZN => n1497);
   U1425 : AOI22_X1 port map( A1 => REGISTERS_1_8_port, A2 => n332, B1 => 
                           REGISTERS_3_8_port, B2 => n315, ZN => n1496);
   U1426 : AOI22_X1 port map( A1 => REGISTERS_4_8_port, A2 => n366, B1 => 
                           REGISTERS_6_8_port, B2 => n349, ZN => n1495);
   U1427 : AOI22_X1 port map( A1 => REGISTERS_0_8_port, A2 => n400, B1 => 
                           REGISTERS_2_8_port, B2 => n383, ZN => n1462);
   U1428 : NAND4_X1 port map( A1 => n1497, A2 => n1496, A3 => n1495, A4 => 
                           n1462, ZN => n1503);
   U1429 : AOI22_X1 port map( A1 => REGISTERS_13_8_port, A2 => n298, B1 => 
                           REGISTERS_15_8_port, B2 => n281, ZN => n1501);
   U1430 : AOI22_X1 port map( A1 => REGISTERS_9_8_port, A2 => n332, B1 => 
                           REGISTERS_11_8_port, B2 => n315, ZN => n1500);
   U1431 : AOI22_X1 port map( A1 => REGISTERS_12_8_port, A2 => n366, B1 => 
                           REGISTERS_14_8_port, B2 => n349, ZN => n1499);
   U1432 : AOI22_X1 port map( A1 => REGISTERS_8_8_port, A2 => n400, B1 => 
                           REGISTERS_10_8_port, B2 => n383, ZN => n1498);
   U1433 : NAND4_X1 port map( A1 => n1501, A2 => n1500, A3 => n1499, A4 => 
                           n1498, ZN => n1502);
   U1434 : AOI22_X1 port map( A1 => n1503, A2 => n3076, B1 => n1502, B2 => 
                           n3074, ZN => n1504);
   U1435 : OAI221_X1 port map( B1 => n3080, B2 => n1506, C1 => n3078, C2 => 
                           n1505, A => n1504, ZN => N212);
   U1436 : AOI22_X1 port map( A1 => REGISTERS_21_9_port, A2 => n299, B1 => 
                           REGISTERS_23_9_port, B2 => n282, ZN => n1510);
   U1437 : AOI22_X1 port map( A1 => REGISTERS_17_9_port, A2 => n333, B1 => 
                           REGISTERS_19_9_port, B2 => n316, ZN => n1509);
   U1438 : AOI22_X1 port map( A1 => REGISTERS_20_9_port, A2 => n367, B1 => 
                           REGISTERS_22_9_port, B2 => n350, ZN => n1508);
   U1439 : AOI22_X1 port map( A1 => REGISTERS_16_9_port, A2 => n401, B1 => 
                           REGISTERS_18_9_port, B2 => n384, ZN => n1507);
   U1440 : AND4_X1 port map( A1 => n1510, A2 => n1509, A3 => n1508, A4 => n1507
                           , ZN => n2615);
   U1441 : AOI22_X1 port map( A1 => REGISTERS_29_9_port, A2 => n299, B1 => 
                           REGISTERS_31_9_port, B2 => n282, ZN => n1514);
   U1442 : AOI22_X1 port map( A1 => REGISTERS_25_9_port, A2 => n333, B1 => 
                           REGISTERS_27_9_port, B2 => n316, ZN => n1513);
   U1443 : AOI22_X1 port map( A1 => REGISTERS_28_9_port, A2 => n367, B1 => 
                           REGISTERS_30_9_port, B2 => n350, ZN => n1512);
   U1444 : AOI22_X1 port map( A1 => REGISTERS_24_9_port, A2 => n401, B1 => 
                           REGISTERS_26_9_port, B2 => n384, ZN => n1511);
   U1445 : AND4_X1 port map( A1 => n1514, A2 => n1513, A3 => n1512, A4 => n1511
                           , ZN => n1526);
   U1446 : AOI22_X1 port map( A1 => REGISTERS_5_9_port, A2 => n299, B1 => 
                           REGISTERS_7_9_port, B2 => n282, ZN => n1518);
   U1447 : AOI22_X1 port map( A1 => REGISTERS_1_9_port, A2 => n333, B1 => 
                           REGISTERS_3_9_port, B2 => n316, ZN => n1517);
   U1448 : AOI22_X1 port map( A1 => REGISTERS_4_9_port, A2 => n367, B1 => 
                           REGISTERS_6_9_port, B2 => n350, ZN => n1516);
   U1449 : AOI22_X1 port map( A1 => REGISTERS_0_9_port, A2 => n401, B1 => 
                           REGISTERS_2_9_port, B2 => n384, ZN => n1515);
   U1450 : NAND4_X1 port map( A1 => n1518, A2 => n1517, A3 => n1516, A4 => 
                           n1515, ZN => n1524);
   U1451 : AOI22_X1 port map( A1 => REGISTERS_13_9_port, A2 => n299, B1 => 
                           REGISTERS_15_9_port, B2 => n282, ZN => n1522);
   U1452 : AOI22_X1 port map( A1 => REGISTERS_9_9_port, A2 => n333, B1 => 
                           REGISTERS_11_9_port, B2 => n316, ZN => n1521);
   U1453 : AOI22_X1 port map( A1 => REGISTERS_12_9_port, A2 => n367, B1 => 
                           REGISTERS_14_9_port, B2 => n350, ZN => n1520);
   U1454 : AOI22_X1 port map( A1 => REGISTERS_8_9_port, A2 => n401, B1 => 
                           REGISTERS_10_9_port, B2 => n384, ZN => n1519);
   U1455 : NAND4_X1 port map( A1 => n1522, A2 => n1521, A3 => n1520, A4 => 
                           n1519, ZN => n1523);
   U1456 : AOI22_X1 port map( A1 => n1524, A2 => n3076, B1 => n1523, B2 => 
                           n3074, ZN => n1525);
   U1457 : OAI221_X1 port map( B1 => n3080, B2 => n2615, C1 => n3078, C2 => 
                           n1526, A => n1525, ZN => N211);
   U1458 : AOI22_X1 port map( A1 => REGISTERS_21_10_port, A2 => n299, B1 => 
                           REGISTERS_23_10_port, B2 => n282, ZN => n2619);
   U1459 : AOI22_X1 port map( A1 => REGISTERS_17_10_port, A2 => n333, B1 => 
                           REGISTERS_19_10_port, B2 => n316, ZN => n2618);
   U1460 : AOI22_X1 port map( A1 => REGISTERS_20_10_port, A2 => n367, B1 => 
                           REGISTERS_22_10_port, B2 => n350, ZN => n2617);
   U1461 : AOI22_X1 port map( A1 => REGISTERS_16_10_port, A2 => n401, B1 => 
                           REGISTERS_18_10_port, B2 => n384, ZN => n2616);
   U1462 : AND4_X1 port map( A1 => n2619, A2 => n2618, A3 => n2617, A4 => n2616
                           , ZN => n2636);
   U1463 : AOI22_X1 port map( A1 => REGISTERS_29_10_port, A2 => n299, B1 => 
                           REGISTERS_31_10_port, B2 => n282, ZN => n2623);
   U1464 : AOI22_X1 port map( A1 => REGISTERS_25_10_port, A2 => n333, B1 => 
                           REGISTERS_27_10_port, B2 => n316, ZN => n2622);
   U1465 : AOI22_X1 port map( A1 => REGISTERS_28_10_port, A2 => n367, B1 => 
                           REGISTERS_30_10_port, B2 => n350, ZN => n2621);
   U1466 : AOI22_X1 port map( A1 => REGISTERS_24_10_port, A2 => n401, B1 => 
                           REGISTERS_26_10_port, B2 => n384, ZN => n2620);
   U1467 : AND4_X1 port map( A1 => n2623, A2 => n2622, A3 => n2621, A4 => n2620
                           , ZN => n2635);
   U1468 : AOI22_X1 port map( A1 => REGISTERS_5_10_port, A2 => n299, B1 => 
                           REGISTERS_7_10_port, B2 => n282, ZN => n2627);
   U1469 : AOI22_X1 port map( A1 => REGISTERS_1_10_port, A2 => n333, B1 => 
                           REGISTERS_3_10_port, B2 => n316, ZN => n2626);
   U1470 : AOI22_X1 port map( A1 => REGISTERS_4_10_port, A2 => n367, B1 => 
                           REGISTERS_6_10_port, B2 => n350, ZN => n2625);
   U1471 : AOI22_X1 port map( A1 => REGISTERS_0_10_port, A2 => n401, B1 => 
                           REGISTERS_2_10_port, B2 => n384, ZN => n2624);
   U1472 : NAND4_X1 port map( A1 => n2627, A2 => n2626, A3 => n2625, A4 => 
                           n2624, ZN => n2633);
   U1473 : AOI22_X1 port map( A1 => REGISTERS_13_10_port, A2 => n299, B1 => 
                           REGISTERS_15_10_port, B2 => n282, ZN => n2631);
   U1474 : AOI22_X1 port map( A1 => REGISTERS_9_10_port, A2 => n333, B1 => 
                           REGISTERS_11_10_port, B2 => n316, ZN => n2630);
   U1475 : AOI22_X1 port map( A1 => REGISTERS_12_10_port, A2 => n367, B1 => 
                           REGISTERS_14_10_port, B2 => n350, ZN => n2629);
   U1476 : AOI22_X1 port map( A1 => REGISTERS_8_10_port, A2 => n401, B1 => 
                           REGISTERS_10_10_port, B2 => n384, ZN => n2628);
   U1477 : NAND4_X1 port map( A1 => n2631, A2 => n2630, A3 => n2629, A4 => 
                           n2628, ZN => n2632);
   U1478 : AOI22_X1 port map( A1 => n2633, A2 => n3076, B1 => n2632, B2 => 
                           n3074, ZN => n2634);
   U1479 : OAI221_X1 port map( B1 => n3080, B2 => n2636, C1 => n3078, C2 => 
                           n2635, A => n2634, ZN => N210);
   U1480 : AOI22_X1 port map( A1 => REGISTERS_21_11_port, A2 => n299, B1 => 
                           REGISTERS_23_11_port, B2 => n282, ZN => n2640);
   U1481 : AOI22_X1 port map( A1 => REGISTERS_17_11_port, A2 => n333, B1 => 
                           REGISTERS_19_11_port, B2 => n316, ZN => n2639);
   U1482 : AOI22_X1 port map( A1 => REGISTERS_20_11_port, A2 => n367, B1 => 
                           REGISTERS_22_11_port, B2 => n350, ZN => n2638);
   U1483 : AOI22_X1 port map( A1 => REGISTERS_16_11_port, A2 => n401, B1 => 
                           REGISTERS_18_11_port, B2 => n384, ZN => n2637);
   U1484 : AND4_X1 port map( A1 => n2640, A2 => n2639, A3 => n2638, A4 => n2637
                           , ZN => n2657);
   U1485 : AOI22_X1 port map( A1 => REGISTERS_29_11_port, A2 => n299, B1 => 
                           REGISTERS_31_11_port, B2 => n282, ZN => n2644);
   U1486 : AOI22_X1 port map( A1 => REGISTERS_25_11_port, A2 => n333, B1 => 
                           REGISTERS_27_11_port, B2 => n316, ZN => n2643);
   U1487 : AOI22_X1 port map( A1 => REGISTERS_28_11_port, A2 => n367, B1 => 
                           REGISTERS_30_11_port, B2 => n350, ZN => n2642);
   U1488 : AOI22_X1 port map( A1 => REGISTERS_24_11_port, A2 => n401, B1 => 
                           REGISTERS_26_11_port, B2 => n384, ZN => n2641);
   U1489 : AND4_X1 port map( A1 => n2644, A2 => n2643, A3 => n2642, A4 => n2641
                           , ZN => n2656);
   U1490 : AOI22_X1 port map( A1 => REGISTERS_5_11_port, A2 => n299, B1 => 
                           REGISTERS_7_11_port, B2 => n282, ZN => n2648);
   U1491 : AOI22_X1 port map( A1 => REGISTERS_1_11_port, A2 => n333, B1 => 
                           REGISTERS_3_11_port, B2 => n316, ZN => n2647);
   U1492 : AOI22_X1 port map( A1 => REGISTERS_4_11_port, A2 => n367, B1 => 
                           REGISTERS_6_11_port, B2 => n350, ZN => n2646);
   U1493 : AOI22_X1 port map( A1 => REGISTERS_0_11_port, A2 => n401, B1 => 
                           REGISTERS_2_11_port, B2 => n384, ZN => n2645);
   U1494 : NAND4_X1 port map( A1 => n2648, A2 => n2647, A3 => n2646, A4 => 
                           n2645, ZN => n2654);
   U1495 : AOI22_X1 port map( A1 => REGISTERS_13_11_port, A2 => n299, B1 => 
                           REGISTERS_15_11_port, B2 => n282, ZN => n2652);
   U1496 : AOI22_X1 port map( A1 => REGISTERS_9_11_port, A2 => n333, B1 => 
                           REGISTERS_11_11_port, B2 => n316, ZN => n2651);
   U1497 : AOI22_X1 port map( A1 => REGISTERS_12_11_port, A2 => n367, B1 => 
                           REGISTERS_14_11_port, B2 => n350, ZN => n2650);
   U1498 : AOI22_X1 port map( A1 => REGISTERS_8_11_port, A2 => n401, B1 => 
                           REGISTERS_10_11_port, B2 => n384, ZN => n2649);
   U1499 : NAND4_X1 port map( A1 => n2652, A2 => n2651, A3 => n2650, A4 => 
                           n2649, ZN => n2653);
   U1500 : AOI22_X1 port map( A1 => n2654, A2 => n3076, B1 => n2653, B2 => 
                           n3074, ZN => n2655);
   U1501 : OAI221_X1 port map( B1 => n3080, B2 => n2657, C1 => n3078, C2 => 
                           n2656, A => n2655, ZN => N209);
   U1502 : AOI22_X1 port map( A1 => REGISTERS_21_12_port, A2 => n300, B1 => 
                           REGISTERS_23_12_port, B2 => n283, ZN => n2661);
   U1503 : AOI22_X1 port map( A1 => REGISTERS_17_12_port, A2 => n334, B1 => 
                           REGISTERS_19_12_port, B2 => n317, ZN => n2660);
   U1504 : AOI22_X1 port map( A1 => REGISTERS_20_12_port, A2 => n368, B1 => 
                           REGISTERS_22_12_port, B2 => n351, ZN => n2659);
   U1505 : AOI22_X1 port map( A1 => REGISTERS_16_12_port, A2 => n402, B1 => 
                           REGISTERS_18_12_port, B2 => n385, ZN => n2658);
   U1506 : AND4_X1 port map( A1 => n2661, A2 => n2660, A3 => n2659, A4 => n2658
                           , ZN => n2678);
   U1507 : AOI22_X1 port map( A1 => REGISTERS_29_12_port, A2 => n300, B1 => 
                           REGISTERS_31_12_port, B2 => n283, ZN => n2665);
   U1508 : AOI22_X1 port map( A1 => REGISTERS_25_12_port, A2 => n334, B1 => 
                           REGISTERS_27_12_port, B2 => n317, ZN => n2664);
   U1509 : AOI22_X1 port map( A1 => REGISTERS_28_12_port, A2 => n368, B1 => 
                           REGISTERS_30_12_port, B2 => n351, ZN => n2663);
   U1510 : AOI22_X1 port map( A1 => REGISTERS_24_12_port, A2 => n402, B1 => 
                           REGISTERS_26_12_port, B2 => n385, ZN => n2662);
   U1511 : AND4_X1 port map( A1 => n2665, A2 => n2664, A3 => n2663, A4 => n2662
                           , ZN => n2677);
   U1512 : AOI22_X1 port map( A1 => REGISTERS_5_12_port, A2 => n300, B1 => 
                           REGISTERS_7_12_port, B2 => n283, ZN => n2669);
   U1513 : AOI22_X1 port map( A1 => REGISTERS_1_12_port, A2 => n334, B1 => 
                           REGISTERS_3_12_port, B2 => n317, ZN => n2668);
   U1514 : AOI22_X1 port map( A1 => REGISTERS_4_12_port, A2 => n368, B1 => 
                           REGISTERS_6_12_port, B2 => n351, ZN => n2667);
   U1515 : AOI22_X1 port map( A1 => REGISTERS_0_12_port, A2 => n402, B1 => 
                           REGISTERS_2_12_port, B2 => n385, ZN => n2666);
   U1516 : NAND4_X1 port map( A1 => n2669, A2 => n2668, A3 => n2667, A4 => 
                           n2666, ZN => n2675);
   U1517 : AOI22_X1 port map( A1 => REGISTERS_13_12_port, A2 => n300, B1 => 
                           REGISTERS_15_12_port, B2 => n283, ZN => n2673);
   U1518 : AOI22_X1 port map( A1 => REGISTERS_9_12_port, A2 => n334, B1 => 
                           REGISTERS_11_12_port, B2 => n317, ZN => n2672);
   U1519 : AOI22_X1 port map( A1 => REGISTERS_12_12_port, A2 => n368, B1 => 
                           REGISTERS_14_12_port, B2 => n351, ZN => n2671);
   U1520 : AOI22_X1 port map( A1 => REGISTERS_8_12_port, A2 => n402, B1 => 
                           REGISTERS_10_12_port, B2 => n385, ZN => n2670);
   U1521 : NAND4_X1 port map( A1 => n2673, A2 => n2672, A3 => n2671, A4 => 
                           n2670, ZN => n2674);
   U1522 : AOI22_X1 port map( A1 => n2675, A2 => n3076, B1 => n2674, B2 => 
                           n3074, ZN => n2676);
   U1523 : OAI221_X1 port map( B1 => n3080, B2 => n2678, C1 => n3078, C2 => 
                           n2677, A => n2676, ZN => N208);
   U1524 : AOI22_X1 port map( A1 => REGISTERS_21_13_port, A2 => n300, B1 => 
                           REGISTERS_23_13_port, B2 => n283, ZN => n2682);
   U1525 : AOI22_X1 port map( A1 => REGISTERS_17_13_port, A2 => n334, B1 => 
                           REGISTERS_19_13_port, B2 => n317, ZN => n2681);
   U1526 : AOI22_X1 port map( A1 => REGISTERS_20_13_port, A2 => n368, B1 => 
                           REGISTERS_22_13_port, B2 => n351, ZN => n2680);
   U1527 : AOI22_X1 port map( A1 => REGISTERS_16_13_port, A2 => n402, B1 => 
                           REGISTERS_18_13_port, B2 => n385, ZN => n2679);
   U1528 : AND4_X1 port map( A1 => n2682, A2 => n2681, A3 => n2680, A4 => n2679
                           , ZN => n2699);
   U1529 : AOI22_X1 port map( A1 => REGISTERS_29_13_port, A2 => n300, B1 => 
                           REGISTERS_31_13_port, B2 => n283, ZN => n2686);
   U1530 : AOI22_X1 port map( A1 => REGISTERS_25_13_port, A2 => n334, B1 => 
                           REGISTERS_27_13_port, B2 => n317, ZN => n2685);
   U1531 : AOI22_X1 port map( A1 => REGISTERS_28_13_port, A2 => n368, B1 => 
                           REGISTERS_30_13_port, B2 => n351, ZN => n2684);
   U1532 : AOI22_X1 port map( A1 => REGISTERS_24_13_port, A2 => n402, B1 => 
                           REGISTERS_26_13_port, B2 => n385, ZN => n2683);
   U1533 : AND4_X1 port map( A1 => n2686, A2 => n2685, A3 => n2684, A4 => n2683
                           , ZN => n2698);
   U1534 : AOI22_X1 port map( A1 => REGISTERS_5_13_port, A2 => n300, B1 => 
                           REGISTERS_7_13_port, B2 => n283, ZN => n2690);
   U1535 : AOI22_X1 port map( A1 => REGISTERS_1_13_port, A2 => n334, B1 => 
                           REGISTERS_3_13_port, B2 => n317, ZN => n2689);
   U1536 : AOI22_X1 port map( A1 => REGISTERS_4_13_port, A2 => n368, B1 => 
                           REGISTERS_6_13_port, B2 => n351, ZN => n2688);
   U1537 : AOI22_X1 port map( A1 => REGISTERS_0_13_port, A2 => n402, B1 => 
                           REGISTERS_2_13_port, B2 => n385, ZN => n2687);
   U1538 : NAND4_X1 port map( A1 => n2690, A2 => n2689, A3 => n2688, A4 => 
                           n2687, ZN => n2696);
   U1539 : AOI22_X1 port map( A1 => REGISTERS_13_13_port, A2 => n300, B1 => 
                           REGISTERS_15_13_port, B2 => n283, ZN => n2694);
   U1540 : AOI22_X1 port map( A1 => REGISTERS_9_13_port, A2 => n334, B1 => 
                           REGISTERS_11_13_port, B2 => n317, ZN => n2693);
   U1541 : AOI22_X1 port map( A1 => REGISTERS_12_13_port, A2 => n368, B1 => 
                           REGISTERS_14_13_port, B2 => n351, ZN => n2692);
   U1542 : AOI22_X1 port map( A1 => REGISTERS_8_13_port, A2 => n402, B1 => 
                           REGISTERS_10_13_port, B2 => n385, ZN => n2691);
   U1543 : NAND4_X1 port map( A1 => n2694, A2 => n2693, A3 => n2692, A4 => 
                           n2691, ZN => n2695);
   U1544 : AOI22_X1 port map( A1 => n2696, A2 => n3076, B1 => n2695, B2 => 
                           n3074, ZN => n2697);
   U1545 : OAI221_X1 port map( B1 => n3080, B2 => n2699, C1 => n3078, C2 => 
                           n2698, A => n2697, ZN => N207);
   U1546 : AOI22_X1 port map( A1 => REGISTERS_21_14_port, A2 => n300, B1 => 
                           REGISTERS_23_14_port, B2 => n283, ZN => n2703);
   U1547 : AOI22_X1 port map( A1 => REGISTERS_17_14_port, A2 => n334, B1 => 
                           REGISTERS_19_14_port, B2 => n317, ZN => n2702);
   U1548 : AOI22_X1 port map( A1 => REGISTERS_20_14_port, A2 => n368, B1 => 
                           REGISTERS_22_14_port, B2 => n351, ZN => n2701);
   U1549 : AOI22_X1 port map( A1 => REGISTERS_16_14_port, A2 => n402, B1 => 
                           REGISTERS_18_14_port, B2 => n385, ZN => n2700);
   U1550 : AND4_X1 port map( A1 => n2703, A2 => n2702, A3 => n2701, A4 => n2700
                           , ZN => n2720);
   U1551 : AOI22_X1 port map( A1 => REGISTERS_29_14_port, A2 => n300, B1 => 
                           REGISTERS_31_14_port, B2 => n283, ZN => n2707);
   U1552 : AOI22_X1 port map( A1 => REGISTERS_25_14_port, A2 => n334, B1 => 
                           REGISTERS_27_14_port, B2 => n317, ZN => n2706);
   U1553 : AOI22_X1 port map( A1 => REGISTERS_28_14_port, A2 => n368, B1 => 
                           REGISTERS_30_14_port, B2 => n351, ZN => n2705);
   U1554 : AOI22_X1 port map( A1 => REGISTERS_24_14_port, A2 => n402, B1 => 
                           REGISTERS_26_14_port, B2 => n385, ZN => n2704);
   U1555 : AND4_X1 port map( A1 => n2707, A2 => n2706, A3 => n2705, A4 => n2704
                           , ZN => n2719);
   U1556 : AOI22_X1 port map( A1 => REGISTERS_5_14_port, A2 => n300, B1 => 
                           REGISTERS_7_14_port, B2 => n283, ZN => n2711);
   U1557 : AOI22_X1 port map( A1 => REGISTERS_1_14_port, A2 => n334, B1 => 
                           REGISTERS_3_14_port, B2 => n317, ZN => n2710);
   U1558 : AOI22_X1 port map( A1 => REGISTERS_4_14_port, A2 => n368, B1 => 
                           REGISTERS_6_14_port, B2 => n351, ZN => n2709);
   U1559 : AOI22_X1 port map( A1 => REGISTERS_0_14_port, A2 => n402, B1 => 
                           REGISTERS_2_14_port, B2 => n385, ZN => n2708);
   U1560 : NAND4_X1 port map( A1 => n2711, A2 => n2710, A3 => n2709, A4 => 
                           n2708, ZN => n2717);
   U1561 : AOI22_X1 port map( A1 => REGISTERS_13_14_port, A2 => n300, B1 => 
                           REGISTERS_15_14_port, B2 => n283, ZN => n2715);
   U1562 : AOI22_X1 port map( A1 => REGISTERS_9_14_port, A2 => n334, B1 => 
                           REGISTERS_11_14_port, B2 => n317, ZN => n2714);
   U1563 : AOI22_X1 port map( A1 => REGISTERS_12_14_port, A2 => n368, B1 => 
                           REGISTERS_14_14_port, B2 => n351, ZN => n2713);
   U1564 : AOI22_X1 port map( A1 => REGISTERS_8_14_port, A2 => n402, B1 => 
                           REGISTERS_10_14_port, B2 => n385, ZN => n2712);
   U1565 : NAND4_X1 port map( A1 => n2715, A2 => n2714, A3 => n2713, A4 => 
                           n2712, ZN => n2716);
   U1566 : AOI22_X1 port map( A1 => n2717, A2 => n3076, B1 => n2716, B2 => 
                           n3074, ZN => n2718);
   U1567 : OAI221_X1 port map( B1 => n3080, B2 => n2720, C1 => n3078, C2 => 
                           n2719, A => n2718, ZN => N206);
   U1568 : AOI22_X1 port map( A1 => REGISTERS_21_15_port, A2 => n301, B1 => 
                           REGISTERS_23_15_port, B2 => n284, ZN => n2724);
   U1569 : AOI22_X1 port map( A1 => REGISTERS_17_15_port, A2 => n335, B1 => 
                           REGISTERS_19_15_port, B2 => n318, ZN => n2723);
   U1570 : AOI22_X1 port map( A1 => REGISTERS_20_15_port, A2 => n369, B1 => 
                           REGISTERS_22_15_port, B2 => n352, ZN => n2722);
   U1571 : AOI22_X1 port map( A1 => REGISTERS_16_15_port, A2 => n403, B1 => 
                           REGISTERS_18_15_port, B2 => n386, ZN => n2721);
   U1572 : AND4_X1 port map( A1 => n2724, A2 => n2723, A3 => n2722, A4 => n2721
                           , ZN => n2741);
   U1573 : AOI22_X1 port map( A1 => REGISTERS_29_15_port, A2 => n301, B1 => 
                           REGISTERS_31_15_port, B2 => n284, ZN => n2728);
   U1574 : AOI22_X1 port map( A1 => REGISTERS_25_15_port, A2 => n335, B1 => 
                           REGISTERS_27_15_port, B2 => n318, ZN => n2727);
   U1575 : AOI22_X1 port map( A1 => REGISTERS_28_15_port, A2 => n369, B1 => 
                           REGISTERS_30_15_port, B2 => n352, ZN => n2726);
   U1576 : AOI22_X1 port map( A1 => REGISTERS_24_15_port, A2 => n403, B1 => 
                           REGISTERS_26_15_port, B2 => n386, ZN => n2725);
   U1577 : AND4_X1 port map( A1 => n2728, A2 => n2727, A3 => n2726, A4 => n2725
                           , ZN => n2740);
   U1578 : AOI22_X1 port map( A1 => REGISTERS_5_15_port, A2 => n301, B1 => 
                           REGISTERS_7_15_port, B2 => n284, ZN => n2732);
   U1579 : AOI22_X1 port map( A1 => REGISTERS_1_15_port, A2 => n335, B1 => 
                           REGISTERS_3_15_port, B2 => n318, ZN => n2731);
   U1580 : AOI22_X1 port map( A1 => REGISTERS_4_15_port, A2 => n369, B1 => 
                           REGISTERS_6_15_port, B2 => n352, ZN => n2730);
   U1581 : AOI22_X1 port map( A1 => REGISTERS_0_15_port, A2 => n403, B1 => 
                           REGISTERS_2_15_port, B2 => n386, ZN => n2729);
   U1582 : NAND4_X1 port map( A1 => n2732, A2 => n2731, A3 => n2730, A4 => 
                           n2729, ZN => n2738);
   U1583 : AOI22_X1 port map( A1 => REGISTERS_13_15_port, A2 => n301, B1 => 
                           REGISTERS_15_15_port, B2 => n284, ZN => n2736);
   U1584 : AOI22_X1 port map( A1 => REGISTERS_9_15_port, A2 => n335, B1 => 
                           REGISTERS_11_15_port, B2 => n318, ZN => n2735);
   U1585 : AOI22_X1 port map( A1 => REGISTERS_12_15_port, A2 => n369, B1 => 
                           REGISTERS_14_15_port, B2 => n352, ZN => n2734);
   U1586 : AOI22_X1 port map( A1 => REGISTERS_8_15_port, A2 => n403, B1 => 
                           REGISTERS_10_15_port, B2 => n386, ZN => n2733);
   U1587 : NAND4_X1 port map( A1 => n2736, A2 => n2735, A3 => n2734, A4 => 
                           n2733, ZN => n2737);
   U1588 : AOI22_X1 port map( A1 => n2738, A2 => n3076, B1 => n2737, B2 => 
                           n3074, ZN => n2739);
   U1589 : OAI221_X1 port map( B1 => n3080, B2 => n2741, C1 => n3078, C2 => 
                           n2740, A => n2739, ZN => N205);
   U1590 : AOI22_X1 port map( A1 => REGISTERS_21_16_port, A2 => n301, B1 => 
                           REGISTERS_23_16_port, B2 => n284, ZN => n2745);
   U1591 : AOI22_X1 port map( A1 => REGISTERS_17_16_port, A2 => n335, B1 => 
                           REGISTERS_19_16_port, B2 => n318, ZN => n2744);
   U1592 : AOI22_X1 port map( A1 => REGISTERS_20_16_port, A2 => n369, B1 => 
                           REGISTERS_22_16_port, B2 => n352, ZN => n2743);
   U1593 : AOI22_X1 port map( A1 => REGISTERS_16_16_port, A2 => n403, B1 => 
                           REGISTERS_18_16_port, B2 => n386, ZN => n2742);
   U1594 : AND4_X1 port map( A1 => n2745, A2 => n2744, A3 => n2743, A4 => n2742
                           , ZN => n2762);
   U1595 : AOI22_X1 port map( A1 => REGISTERS_29_16_port, A2 => n301, B1 => 
                           REGISTERS_31_16_port, B2 => n284, ZN => n2749);
   U1596 : AOI22_X1 port map( A1 => REGISTERS_25_16_port, A2 => n335, B1 => 
                           REGISTERS_27_16_port, B2 => n318, ZN => n2748);
   U1597 : AOI22_X1 port map( A1 => REGISTERS_28_16_port, A2 => n369, B1 => 
                           REGISTERS_30_16_port, B2 => n352, ZN => n2747);
   U1598 : AOI22_X1 port map( A1 => REGISTERS_24_16_port, A2 => n403, B1 => 
                           REGISTERS_26_16_port, B2 => n386, ZN => n2746);
   U1599 : AND4_X1 port map( A1 => n2749, A2 => n2748, A3 => n2747, A4 => n2746
                           , ZN => n2761);
   U1600 : AOI22_X1 port map( A1 => REGISTERS_5_16_port, A2 => n301, B1 => 
                           REGISTERS_7_16_port, B2 => n284, ZN => n2753);
   U1601 : AOI22_X1 port map( A1 => REGISTERS_1_16_port, A2 => n335, B1 => 
                           REGISTERS_3_16_port, B2 => n318, ZN => n2752);
   U1602 : AOI22_X1 port map( A1 => REGISTERS_4_16_port, A2 => n369, B1 => 
                           REGISTERS_6_16_port, B2 => n352, ZN => n2751);
   U1603 : AOI22_X1 port map( A1 => REGISTERS_0_16_port, A2 => n403, B1 => 
                           REGISTERS_2_16_port, B2 => n386, ZN => n2750);
   U1604 : NAND4_X1 port map( A1 => n2753, A2 => n2752, A3 => n2751, A4 => 
                           n2750, ZN => n2759);
   U1605 : AOI22_X1 port map( A1 => REGISTERS_13_16_port, A2 => n301, B1 => 
                           REGISTERS_15_16_port, B2 => n284, ZN => n2757);
   U1606 : AOI22_X1 port map( A1 => REGISTERS_9_16_port, A2 => n335, B1 => 
                           REGISTERS_11_16_port, B2 => n318, ZN => n2756);
   U1607 : AOI22_X1 port map( A1 => REGISTERS_12_16_port, A2 => n369, B1 => 
                           REGISTERS_14_16_port, B2 => n352, ZN => n2755);
   U1608 : AOI22_X1 port map( A1 => REGISTERS_8_16_port, A2 => n403, B1 => 
                           REGISTERS_10_16_port, B2 => n386, ZN => n2754);
   U1609 : NAND4_X1 port map( A1 => n2757, A2 => n2756, A3 => n2755, A4 => 
                           n2754, ZN => n2758);
   U1610 : AOI22_X1 port map( A1 => n2759, A2 => n3076, B1 => n2758, B2 => 
                           n3074, ZN => n2760);
   U1611 : OAI221_X1 port map( B1 => n3080, B2 => n2762, C1 => n3078, C2 => 
                           n2761, A => n2760, ZN => N204);
   U1612 : AOI22_X1 port map( A1 => REGISTERS_21_17_port, A2 => n301, B1 => 
                           REGISTERS_23_17_port, B2 => n284, ZN => n2766);
   U1613 : AOI22_X1 port map( A1 => REGISTERS_17_17_port, A2 => n335, B1 => 
                           REGISTERS_19_17_port, B2 => n318, ZN => n2765);
   U1614 : AOI22_X1 port map( A1 => REGISTERS_20_17_port, A2 => n369, B1 => 
                           REGISTERS_22_17_port, B2 => n352, ZN => n2764);
   U1615 : AOI22_X1 port map( A1 => REGISTERS_16_17_port, A2 => n403, B1 => 
                           REGISTERS_18_17_port, B2 => n386, ZN => n2763);
   U1616 : AND4_X1 port map( A1 => n2766, A2 => n2765, A3 => n2764, A4 => n2763
                           , ZN => n2783);
   U1617 : AOI22_X1 port map( A1 => REGISTERS_29_17_port, A2 => n301, B1 => 
                           REGISTERS_31_17_port, B2 => n284, ZN => n2770);
   U1618 : AOI22_X1 port map( A1 => REGISTERS_25_17_port, A2 => n335, B1 => 
                           REGISTERS_27_17_port, B2 => n318, ZN => n2769);
   U1619 : AOI22_X1 port map( A1 => REGISTERS_28_17_port, A2 => n369, B1 => 
                           REGISTERS_30_17_port, B2 => n352, ZN => n2768);
   U1620 : AOI22_X1 port map( A1 => REGISTERS_24_17_port, A2 => n403, B1 => 
                           REGISTERS_26_17_port, B2 => n386, ZN => n2767);
   U1621 : AND4_X1 port map( A1 => n2770, A2 => n2769, A3 => n2768, A4 => n2767
                           , ZN => n2782);
   U1622 : AOI22_X1 port map( A1 => REGISTERS_5_17_port, A2 => n301, B1 => 
                           REGISTERS_7_17_port, B2 => n284, ZN => n2774);
   U1623 : AOI22_X1 port map( A1 => REGISTERS_1_17_port, A2 => n335, B1 => 
                           REGISTERS_3_17_port, B2 => n318, ZN => n2773);
   U1624 : AOI22_X1 port map( A1 => REGISTERS_4_17_port, A2 => n369, B1 => 
                           REGISTERS_6_17_port, B2 => n352, ZN => n2772);
   U1625 : AOI22_X1 port map( A1 => REGISTERS_0_17_port, A2 => n403, B1 => 
                           REGISTERS_2_17_port, B2 => n386, ZN => n2771);
   U1626 : NAND4_X1 port map( A1 => n2774, A2 => n2773, A3 => n2772, A4 => 
                           n2771, ZN => n2780);
   U1627 : AOI22_X1 port map( A1 => REGISTERS_13_17_port, A2 => n301, B1 => 
                           REGISTERS_15_17_port, B2 => n284, ZN => n2778);
   U1628 : AOI22_X1 port map( A1 => REGISTERS_9_17_port, A2 => n335, B1 => 
                           REGISTERS_11_17_port, B2 => n318, ZN => n2777);
   U1629 : AOI22_X1 port map( A1 => REGISTERS_12_17_port, A2 => n369, B1 => 
                           REGISTERS_14_17_port, B2 => n352, ZN => n2776);
   U1630 : AOI22_X1 port map( A1 => REGISTERS_8_17_port, A2 => n403, B1 => 
                           REGISTERS_10_17_port, B2 => n386, ZN => n2775);
   U1631 : NAND4_X1 port map( A1 => n2778, A2 => n2777, A3 => n2776, A4 => 
                           n2775, ZN => n2779);
   U1632 : AOI22_X1 port map( A1 => n2780, A2 => n3076, B1 => n2779, B2 => 
                           n3074, ZN => n2781);
   U1633 : OAI221_X1 port map( B1 => n3080, B2 => n2783, C1 => n3078, C2 => 
                           n2782, A => n2781, ZN => N203);
   U1634 : AOI22_X1 port map( A1 => REGISTERS_21_18_port, A2 => n302, B1 => 
                           REGISTERS_23_18_port, B2 => n285, ZN => n2787);
   U1635 : AOI22_X1 port map( A1 => REGISTERS_17_18_port, A2 => n336, B1 => 
                           REGISTERS_19_18_port, B2 => n319, ZN => n2786);
   U1636 : AOI22_X1 port map( A1 => REGISTERS_20_18_port, A2 => n370, B1 => 
                           REGISTERS_22_18_port, B2 => n353, ZN => n2785);
   U1637 : AOI22_X1 port map( A1 => REGISTERS_16_18_port, A2 => n404, B1 => 
                           REGISTERS_18_18_port, B2 => n387, ZN => n2784);
   U1638 : AND4_X1 port map( A1 => n2787, A2 => n2786, A3 => n2785, A4 => n2784
                           , ZN => n2804);
   U1639 : AOI22_X1 port map( A1 => REGISTERS_29_18_port, A2 => n302, B1 => 
                           REGISTERS_31_18_port, B2 => n285, ZN => n2791);
   U1640 : AOI22_X1 port map( A1 => REGISTERS_25_18_port, A2 => n336, B1 => 
                           REGISTERS_27_18_port, B2 => n319, ZN => n2790);
   U1641 : AOI22_X1 port map( A1 => REGISTERS_28_18_port, A2 => n370, B1 => 
                           REGISTERS_30_18_port, B2 => n353, ZN => n2789);
   U1642 : AOI22_X1 port map( A1 => REGISTERS_24_18_port, A2 => n404, B1 => 
                           REGISTERS_26_18_port, B2 => n387, ZN => n2788);
   U1643 : AND4_X1 port map( A1 => n2791, A2 => n2790, A3 => n2789, A4 => n2788
                           , ZN => n2803);
   U1644 : AOI22_X1 port map( A1 => REGISTERS_5_18_port, A2 => n302, B1 => 
                           REGISTERS_7_18_port, B2 => n285, ZN => n2795);
   U1645 : AOI22_X1 port map( A1 => REGISTERS_1_18_port, A2 => n336, B1 => 
                           REGISTERS_3_18_port, B2 => n319, ZN => n2794);
   U1646 : AOI22_X1 port map( A1 => REGISTERS_4_18_port, A2 => n370, B1 => 
                           REGISTERS_6_18_port, B2 => n353, ZN => n2793);
   U1647 : AOI22_X1 port map( A1 => REGISTERS_0_18_port, A2 => n404, B1 => 
                           REGISTERS_2_18_port, B2 => n387, ZN => n2792);
   U1648 : NAND4_X1 port map( A1 => n2795, A2 => n2794, A3 => n2793, A4 => 
                           n2792, ZN => n2801);
   U1649 : AOI22_X1 port map( A1 => REGISTERS_13_18_port, A2 => n302, B1 => 
                           REGISTERS_15_18_port, B2 => n285, ZN => n2799);
   U1650 : AOI22_X1 port map( A1 => REGISTERS_9_18_port, A2 => n336, B1 => 
                           REGISTERS_11_18_port, B2 => n319, ZN => n2798);
   U1651 : AOI22_X1 port map( A1 => REGISTERS_12_18_port, A2 => n370, B1 => 
                           REGISTERS_14_18_port, B2 => n353, ZN => n2797);
   U1652 : AOI22_X1 port map( A1 => REGISTERS_8_18_port, A2 => n404, B1 => 
                           REGISTERS_10_18_port, B2 => n387, ZN => n2796);
   U1653 : NAND4_X1 port map( A1 => n2799, A2 => n2798, A3 => n2797, A4 => 
                           n2796, ZN => n2800);
   U1654 : AOI22_X1 port map( A1 => n2801, A2 => n3076, B1 => n2800, B2 => 
                           n3074, ZN => n2802);
   U1655 : OAI221_X1 port map( B1 => n3080, B2 => n2804, C1 => n3078, C2 => 
                           n2803, A => n2802, ZN => N202);
   U1656 : AOI22_X1 port map( A1 => REGISTERS_21_19_port, A2 => n302, B1 => 
                           REGISTERS_23_19_port, B2 => n285, ZN => n2808);
   U1657 : AOI22_X1 port map( A1 => REGISTERS_17_19_port, A2 => n336, B1 => 
                           REGISTERS_19_19_port, B2 => n319, ZN => n2807);
   U1658 : AOI22_X1 port map( A1 => REGISTERS_20_19_port, A2 => n370, B1 => 
                           REGISTERS_22_19_port, B2 => n353, ZN => n2806);
   U1659 : AOI22_X1 port map( A1 => REGISTERS_16_19_port, A2 => n404, B1 => 
                           REGISTERS_18_19_port, B2 => n387, ZN => n2805);
   U1660 : AND4_X1 port map( A1 => n2808, A2 => n2807, A3 => n2806, A4 => n2805
                           , ZN => n2825);
   U1661 : AOI22_X1 port map( A1 => REGISTERS_29_19_port, A2 => n302, B1 => 
                           REGISTERS_31_19_port, B2 => n285, ZN => n2812);
   U1662 : AOI22_X1 port map( A1 => REGISTERS_25_19_port, A2 => n336, B1 => 
                           REGISTERS_27_19_port, B2 => n319, ZN => n2811);
   U1663 : AOI22_X1 port map( A1 => REGISTERS_28_19_port, A2 => n370, B1 => 
                           REGISTERS_30_19_port, B2 => n353, ZN => n2810);
   U1664 : AOI22_X1 port map( A1 => REGISTERS_24_19_port, A2 => n404, B1 => 
                           REGISTERS_26_19_port, B2 => n387, ZN => n2809);
   U1665 : AND4_X1 port map( A1 => n2812, A2 => n2811, A3 => n2810, A4 => n2809
                           , ZN => n2824);
   U1666 : AOI22_X1 port map( A1 => REGISTERS_5_19_port, A2 => n302, B1 => 
                           REGISTERS_7_19_port, B2 => n285, ZN => n2816);
   U1667 : AOI22_X1 port map( A1 => REGISTERS_1_19_port, A2 => n336, B1 => 
                           REGISTERS_3_19_port, B2 => n319, ZN => n2815);
   U1668 : AOI22_X1 port map( A1 => REGISTERS_4_19_port, A2 => n370, B1 => 
                           REGISTERS_6_19_port, B2 => n353, ZN => n2814);
   U1669 : AOI22_X1 port map( A1 => REGISTERS_0_19_port, A2 => n404, B1 => 
                           REGISTERS_2_19_port, B2 => n387, ZN => n2813);
   U1670 : NAND4_X1 port map( A1 => n2816, A2 => n2815, A3 => n2814, A4 => 
                           n2813, ZN => n2822);
   U1671 : AOI22_X1 port map( A1 => REGISTERS_13_19_port, A2 => n302, B1 => 
                           REGISTERS_15_19_port, B2 => n285, ZN => n2820);
   U1672 : AOI22_X1 port map( A1 => REGISTERS_9_19_port, A2 => n336, B1 => 
                           REGISTERS_11_19_port, B2 => n319, ZN => n2819);
   U1673 : AOI22_X1 port map( A1 => REGISTERS_12_19_port, A2 => n370, B1 => 
                           REGISTERS_14_19_port, B2 => n353, ZN => n2818);
   U1674 : AOI22_X1 port map( A1 => REGISTERS_8_19_port, A2 => n404, B1 => 
                           REGISTERS_10_19_port, B2 => n387, ZN => n2817);
   U1675 : NAND4_X1 port map( A1 => n2820, A2 => n2819, A3 => n2818, A4 => 
                           n2817, ZN => n2821);
   U1676 : AOI22_X1 port map( A1 => n2822, A2 => n3076, B1 => n2821, B2 => 
                           n3074, ZN => n2823);
   U1677 : OAI221_X1 port map( B1 => n3080, B2 => n2825, C1 => n3078, C2 => 
                           n2824, A => n2823, ZN => N201);
   U1678 : AOI22_X1 port map( A1 => REGISTERS_21_20_port, A2 => n302, B1 => 
                           REGISTERS_23_20_port, B2 => n285, ZN => n2829);
   U1679 : AOI22_X1 port map( A1 => REGISTERS_17_20_port, A2 => n336, B1 => 
                           REGISTERS_19_20_port, B2 => n319, ZN => n2828);
   U1680 : AOI22_X1 port map( A1 => REGISTERS_20_20_port, A2 => n370, B1 => 
                           REGISTERS_22_20_port, B2 => n353, ZN => n2827);
   U1681 : AOI22_X1 port map( A1 => REGISTERS_16_20_port, A2 => n404, B1 => 
                           REGISTERS_18_20_port, B2 => n387, ZN => n2826);
   U1682 : AND4_X1 port map( A1 => n2829, A2 => n2828, A3 => n2827, A4 => n2826
                           , ZN => n2846);
   U1683 : AOI22_X1 port map( A1 => REGISTERS_29_20_port, A2 => n302, B1 => 
                           REGISTERS_31_20_port, B2 => n285, ZN => n2833);
   U1684 : AOI22_X1 port map( A1 => REGISTERS_25_20_port, A2 => n336, B1 => 
                           REGISTERS_27_20_port, B2 => n319, ZN => n2832);
   U1685 : AOI22_X1 port map( A1 => REGISTERS_28_20_port, A2 => n370, B1 => 
                           REGISTERS_30_20_port, B2 => n353, ZN => n2831);
   U1686 : AOI22_X1 port map( A1 => REGISTERS_24_20_port, A2 => n404, B1 => 
                           REGISTERS_26_20_port, B2 => n387, ZN => n2830);
   U1687 : AND4_X1 port map( A1 => n2833, A2 => n2832, A3 => n2831, A4 => n2830
                           , ZN => n2845);
   U1688 : AOI22_X1 port map( A1 => REGISTERS_5_20_port, A2 => n302, B1 => 
                           REGISTERS_7_20_port, B2 => n285, ZN => n2837);
   U1689 : AOI22_X1 port map( A1 => REGISTERS_1_20_port, A2 => n336, B1 => 
                           REGISTERS_3_20_port, B2 => n319, ZN => n2836);
   U1690 : AOI22_X1 port map( A1 => REGISTERS_4_20_port, A2 => n370, B1 => 
                           REGISTERS_6_20_port, B2 => n353, ZN => n2835);
   U1691 : AOI22_X1 port map( A1 => REGISTERS_0_20_port, A2 => n404, B1 => 
                           REGISTERS_2_20_port, B2 => n387, ZN => n2834);
   U1692 : NAND4_X1 port map( A1 => n2837, A2 => n2836, A3 => n2835, A4 => 
                           n2834, ZN => n2843);
   U1693 : AOI22_X1 port map( A1 => REGISTERS_13_20_port, A2 => n302, B1 => 
                           REGISTERS_15_20_port, B2 => n285, ZN => n2841);
   U1694 : AOI22_X1 port map( A1 => REGISTERS_9_20_port, A2 => n336, B1 => 
                           REGISTERS_11_20_port, B2 => n319, ZN => n2840);
   U1695 : AOI22_X1 port map( A1 => REGISTERS_12_20_port, A2 => n370, B1 => 
                           REGISTERS_14_20_port, B2 => n353, ZN => n2839);
   U1696 : AOI22_X1 port map( A1 => REGISTERS_8_20_port, A2 => n404, B1 => 
                           REGISTERS_10_20_port, B2 => n387, ZN => n2838);
   U1697 : NAND4_X1 port map( A1 => n2841, A2 => n2840, A3 => n2839, A4 => 
                           n2838, ZN => n2842);
   U1698 : AOI22_X1 port map( A1 => n2843, A2 => n3076, B1 => n2842, B2 => 
                           n3074, ZN => n2844);
   U1699 : OAI221_X1 port map( B1 => n3080, B2 => n2846, C1 => n3078, C2 => 
                           n2845, A => n2844, ZN => N200);
   U1700 : AOI22_X1 port map( A1 => REGISTERS_21_21_port, A2 => n303, B1 => 
                           REGISTERS_23_21_port, B2 => n286, ZN => n2850);
   U1701 : AOI22_X1 port map( A1 => REGISTERS_17_21_port, A2 => n337, B1 => 
                           REGISTERS_19_21_port, B2 => n320, ZN => n2849);
   U1702 : AOI22_X1 port map( A1 => REGISTERS_20_21_port, A2 => n371, B1 => 
                           REGISTERS_22_21_port, B2 => n354, ZN => n2848);
   U1703 : AOI22_X1 port map( A1 => REGISTERS_16_21_port, A2 => n405, B1 => 
                           REGISTERS_18_21_port, B2 => n388, ZN => n2847);
   U1704 : AND4_X1 port map( A1 => n2850, A2 => n2849, A3 => n2848, A4 => n2847
                           , ZN => n2867);
   U1705 : AOI22_X1 port map( A1 => REGISTERS_29_21_port, A2 => n303, B1 => 
                           REGISTERS_31_21_port, B2 => n286, ZN => n2854);
   U1706 : AOI22_X1 port map( A1 => REGISTERS_25_21_port, A2 => n337, B1 => 
                           REGISTERS_27_21_port, B2 => n320, ZN => n2853);
   U1707 : AOI22_X1 port map( A1 => REGISTERS_28_21_port, A2 => n371, B1 => 
                           REGISTERS_30_21_port, B2 => n354, ZN => n2852);
   U1708 : AOI22_X1 port map( A1 => REGISTERS_24_21_port, A2 => n405, B1 => 
                           REGISTERS_26_21_port, B2 => n388, ZN => n2851);
   U1709 : AND4_X1 port map( A1 => n2854, A2 => n2853, A3 => n2852, A4 => n2851
                           , ZN => n2866);
   U1710 : AOI22_X1 port map( A1 => REGISTERS_5_21_port, A2 => n303, B1 => 
                           REGISTERS_7_21_port, B2 => n286, ZN => n2858);
   U1711 : AOI22_X1 port map( A1 => REGISTERS_1_21_port, A2 => n337, B1 => 
                           REGISTERS_3_21_port, B2 => n320, ZN => n2857);
   U1712 : AOI22_X1 port map( A1 => REGISTERS_4_21_port, A2 => n371, B1 => 
                           REGISTERS_6_21_port, B2 => n354, ZN => n2856);
   U1713 : AOI22_X1 port map( A1 => REGISTERS_0_21_port, A2 => n405, B1 => 
                           REGISTERS_2_21_port, B2 => n388, ZN => n2855);
   U1714 : NAND4_X1 port map( A1 => n2858, A2 => n2857, A3 => n2856, A4 => 
                           n2855, ZN => n2864);
   U1715 : AOI22_X1 port map( A1 => REGISTERS_13_21_port, A2 => n303, B1 => 
                           REGISTERS_15_21_port, B2 => n286, ZN => n2862);
   U1716 : AOI22_X1 port map( A1 => REGISTERS_9_21_port, A2 => n337, B1 => 
                           REGISTERS_11_21_port, B2 => n320, ZN => n2861);
   U1717 : AOI22_X1 port map( A1 => REGISTERS_12_21_port, A2 => n371, B1 => 
                           REGISTERS_14_21_port, B2 => n354, ZN => n2860);
   U1718 : AOI22_X1 port map( A1 => REGISTERS_8_21_port, A2 => n405, B1 => 
                           REGISTERS_10_21_port, B2 => n388, ZN => n2859);
   U1719 : NAND4_X1 port map( A1 => n2862, A2 => n2861, A3 => n2860, A4 => 
                           n2859, ZN => n2863);
   U1720 : AOI22_X1 port map( A1 => n2864, A2 => n3076, B1 => n2863, B2 => 
                           n3074, ZN => n2865);
   U1721 : OAI221_X1 port map( B1 => n3080, B2 => n2867, C1 => n3078, C2 => 
                           n2866, A => n2865, ZN => N199);
   U1722 : AOI22_X1 port map( A1 => REGISTERS_21_22_port, A2 => n303, B1 => 
                           REGISTERS_23_22_port, B2 => n286, ZN => n2871);
   U1723 : AOI22_X1 port map( A1 => REGISTERS_17_22_port, A2 => n337, B1 => 
                           REGISTERS_19_22_port, B2 => n320, ZN => n2870);
   U1724 : AOI22_X1 port map( A1 => REGISTERS_20_22_port, A2 => n371, B1 => 
                           REGISTERS_22_22_port, B2 => n354, ZN => n2869);
   U1725 : AOI22_X1 port map( A1 => REGISTERS_16_22_port, A2 => n405, B1 => 
                           REGISTERS_18_22_port, B2 => n388, ZN => n2868);
   U1726 : AND4_X1 port map( A1 => n2871, A2 => n2870, A3 => n2869, A4 => n2868
                           , ZN => n2888);
   U1727 : AOI22_X1 port map( A1 => REGISTERS_29_22_port, A2 => n303, B1 => 
                           REGISTERS_31_22_port, B2 => n286, ZN => n2875);
   U1728 : AOI22_X1 port map( A1 => REGISTERS_25_22_port, A2 => n337, B1 => 
                           REGISTERS_27_22_port, B2 => n320, ZN => n2874);
   U1729 : AOI22_X1 port map( A1 => REGISTERS_28_22_port, A2 => n371, B1 => 
                           REGISTERS_30_22_port, B2 => n354, ZN => n2873);
   U1730 : AOI22_X1 port map( A1 => REGISTERS_24_22_port, A2 => n405, B1 => 
                           REGISTERS_26_22_port, B2 => n388, ZN => n2872);
   U1731 : AND4_X1 port map( A1 => n2875, A2 => n2874, A3 => n2873, A4 => n2872
                           , ZN => n2887);
   U1732 : AOI22_X1 port map( A1 => REGISTERS_5_22_port, A2 => n303, B1 => 
                           REGISTERS_7_22_port, B2 => n286, ZN => n2879);
   U1733 : AOI22_X1 port map( A1 => REGISTERS_1_22_port, A2 => n337, B1 => 
                           REGISTERS_3_22_port, B2 => n320, ZN => n2878);
   U1734 : AOI22_X1 port map( A1 => REGISTERS_4_22_port, A2 => n371, B1 => 
                           REGISTERS_6_22_port, B2 => n354, ZN => n2877);
   U1735 : AOI22_X1 port map( A1 => REGISTERS_0_22_port, A2 => n405, B1 => 
                           REGISTERS_2_22_port, B2 => n388, ZN => n2876);
   U1736 : NAND4_X1 port map( A1 => n2879, A2 => n2878, A3 => n2877, A4 => 
                           n2876, ZN => n2885);
   U1737 : AOI22_X1 port map( A1 => REGISTERS_13_22_port, A2 => n303, B1 => 
                           REGISTERS_15_22_port, B2 => n286, ZN => n2883);
   U1738 : AOI22_X1 port map( A1 => REGISTERS_9_22_port, A2 => n337, B1 => 
                           REGISTERS_11_22_port, B2 => n320, ZN => n2882);
   U1739 : AOI22_X1 port map( A1 => REGISTERS_12_22_port, A2 => n371, B1 => 
                           REGISTERS_14_22_port, B2 => n354, ZN => n2881);
   U1740 : AOI22_X1 port map( A1 => REGISTERS_8_22_port, A2 => n405, B1 => 
                           REGISTERS_10_22_port, B2 => n388, ZN => n2880);
   U1741 : NAND4_X1 port map( A1 => n2883, A2 => n2882, A3 => n2881, A4 => 
                           n2880, ZN => n2884);
   U1742 : AOI22_X1 port map( A1 => n2885, A2 => n3076, B1 => n2884, B2 => 
                           n3074, ZN => n2886);
   U1743 : OAI221_X1 port map( B1 => n3080, B2 => n2888, C1 => n3078, C2 => 
                           n2887, A => n2886, ZN => N198);
   U1744 : AOI22_X1 port map( A1 => REGISTERS_21_23_port, A2 => n303, B1 => 
                           REGISTERS_23_23_port, B2 => n286, ZN => n2892);
   U1745 : AOI22_X1 port map( A1 => REGISTERS_17_23_port, A2 => n337, B1 => 
                           REGISTERS_19_23_port, B2 => n320, ZN => n2891);
   U1746 : AOI22_X1 port map( A1 => REGISTERS_20_23_port, A2 => n371, B1 => 
                           REGISTERS_22_23_port, B2 => n354, ZN => n2890);
   U1747 : AOI22_X1 port map( A1 => REGISTERS_16_23_port, A2 => n405, B1 => 
                           REGISTERS_18_23_port, B2 => n388, ZN => n2889);
   U1748 : AND4_X1 port map( A1 => n2892, A2 => n2891, A3 => n2890, A4 => n2889
                           , ZN => n2909);
   U1749 : AOI22_X1 port map( A1 => REGISTERS_29_23_port, A2 => n303, B1 => 
                           REGISTERS_31_23_port, B2 => n286, ZN => n2896);
   U1750 : AOI22_X1 port map( A1 => REGISTERS_25_23_port, A2 => n337, B1 => 
                           REGISTERS_27_23_port, B2 => n320, ZN => n2895);
   U1751 : AOI22_X1 port map( A1 => REGISTERS_28_23_port, A2 => n371, B1 => 
                           REGISTERS_30_23_port, B2 => n354, ZN => n2894);
   U1752 : AOI22_X1 port map( A1 => REGISTERS_24_23_port, A2 => n405, B1 => 
                           REGISTERS_26_23_port, B2 => n388, ZN => n2893);
   U1753 : AND4_X1 port map( A1 => n2896, A2 => n2895, A3 => n2894, A4 => n2893
                           , ZN => n2908);
   U1754 : AOI22_X1 port map( A1 => REGISTERS_5_23_port, A2 => n303, B1 => 
                           REGISTERS_7_23_port, B2 => n286, ZN => n2900);
   U1755 : AOI22_X1 port map( A1 => REGISTERS_1_23_port, A2 => n337, B1 => 
                           REGISTERS_3_23_port, B2 => n320, ZN => n2899);
   U1756 : AOI22_X1 port map( A1 => REGISTERS_4_23_port, A2 => n371, B1 => 
                           REGISTERS_6_23_port, B2 => n354, ZN => n2898);
   U1757 : AOI22_X1 port map( A1 => REGISTERS_0_23_port, A2 => n405, B1 => 
                           REGISTERS_2_23_port, B2 => n388, ZN => n2897);
   U1758 : NAND4_X1 port map( A1 => n2900, A2 => n2899, A3 => n2898, A4 => 
                           n2897, ZN => n2906);
   U1759 : AOI22_X1 port map( A1 => REGISTERS_13_23_port, A2 => n303, B1 => 
                           REGISTERS_15_23_port, B2 => n286, ZN => n2904);
   U1760 : AOI22_X1 port map( A1 => REGISTERS_9_23_port, A2 => n337, B1 => 
                           REGISTERS_11_23_port, B2 => n320, ZN => n2903);
   U1761 : AOI22_X1 port map( A1 => REGISTERS_12_23_port, A2 => n371, B1 => 
                           REGISTERS_14_23_port, B2 => n354, ZN => n2902);
   U1762 : AOI22_X1 port map( A1 => REGISTERS_8_23_port, A2 => n405, B1 => 
                           REGISTERS_10_23_port, B2 => n388, ZN => n2901);
   U1763 : NAND4_X1 port map( A1 => n2904, A2 => n2903, A3 => n2902, A4 => 
                           n2901, ZN => n2905);
   U1764 : AOI22_X1 port map( A1 => n2906, A2 => n3076, B1 => n2905, B2 => 
                           n3074, ZN => n2907);
   U1765 : OAI221_X1 port map( B1 => n3080, B2 => n2909, C1 => n3078, C2 => 
                           n2908, A => n2907, ZN => N197);
   U1766 : AOI22_X1 port map( A1 => REGISTERS_21_24_port, A2 => n304, B1 => 
                           REGISTERS_23_24_port, B2 => n287, ZN => n2913);
   U1767 : AOI22_X1 port map( A1 => REGISTERS_17_24_port, A2 => n338, B1 => 
                           REGISTERS_19_24_port, B2 => n321, ZN => n2912);
   U1768 : AOI22_X1 port map( A1 => REGISTERS_20_24_port, A2 => n372, B1 => 
                           REGISTERS_22_24_port, B2 => n355, ZN => n2911);
   U1769 : AOI22_X1 port map( A1 => REGISTERS_16_24_port, A2 => n406, B1 => 
                           REGISTERS_18_24_port, B2 => n389, ZN => n2910);
   U1770 : AND4_X1 port map( A1 => n2913, A2 => n2912, A3 => n2911, A4 => n2910
                           , ZN => n2930);
   U1771 : AOI22_X1 port map( A1 => REGISTERS_29_24_port, A2 => n304, B1 => 
                           REGISTERS_31_24_port, B2 => n287, ZN => n2917);
   U1772 : AOI22_X1 port map( A1 => REGISTERS_25_24_port, A2 => n338, B1 => 
                           REGISTERS_27_24_port, B2 => n321, ZN => n2916);
   U1773 : AOI22_X1 port map( A1 => REGISTERS_28_24_port, A2 => n372, B1 => 
                           REGISTERS_30_24_port, B2 => n355, ZN => n2915);
   U1774 : AOI22_X1 port map( A1 => REGISTERS_24_24_port, A2 => n406, B1 => 
                           REGISTERS_26_24_port, B2 => n389, ZN => n2914);
   U1775 : AND4_X1 port map( A1 => n2917, A2 => n2916, A3 => n2915, A4 => n2914
                           , ZN => n2929);
   U1776 : AOI22_X1 port map( A1 => REGISTERS_5_24_port, A2 => n304, B1 => 
                           REGISTERS_7_24_port, B2 => n287, ZN => n2921);
   U1777 : AOI22_X1 port map( A1 => REGISTERS_1_24_port, A2 => n338, B1 => 
                           REGISTERS_3_24_port, B2 => n321, ZN => n2920);
   U1778 : AOI22_X1 port map( A1 => REGISTERS_4_24_port, A2 => n372, B1 => 
                           REGISTERS_6_24_port, B2 => n355, ZN => n2919);
   U1779 : AOI22_X1 port map( A1 => REGISTERS_0_24_port, A2 => n406, B1 => 
                           REGISTERS_2_24_port, B2 => n389, ZN => n2918);
   U1780 : NAND4_X1 port map( A1 => n2921, A2 => n2920, A3 => n2919, A4 => 
                           n2918, ZN => n2927);
   U1781 : AOI22_X1 port map( A1 => REGISTERS_13_24_port, A2 => n304, B1 => 
                           REGISTERS_15_24_port, B2 => n287, ZN => n2925);
   U1782 : AOI22_X1 port map( A1 => REGISTERS_9_24_port, A2 => n338, B1 => 
                           REGISTERS_11_24_port, B2 => n321, ZN => n2924);
   U1783 : AOI22_X1 port map( A1 => REGISTERS_12_24_port, A2 => n372, B1 => 
                           REGISTERS_14_24_port, B2 => n355, ZN => n2923);
   U1784 : AOI22_X1 port map( A1 => REGISTERS_8_24_port, A2 => n406, B1 => 
                           REGISTERS_10_24_port, B2 => n389, ZN => n2922);
   U1785 : NAND4_X1 port map( A1 => n2925, A2 => n2924, A3 => n2923, A4 => 
                           n2922, ZN => n2926);
   U1786 : AOI22_X1 port map( A1 => n2927, A2 => n3076, B1 => n2926, B2 => 
                           n3074, ZN => n2928);
   U1787 : OAI221_X1 port map( B1 => n3080, B2 => n2930, C1 => n3078, C2 => 
                           n2929, A => n2928, ZN => N196);
   U1788 : AOI22_X1 port map( A1 => REGISTERS_21_25_port, A2 => n304, B1 => 
                           REGISTERS_23_25_port, B2 => n287, ZN => n2934);
   U1789 : AOI22_X1 port map( A1 => REGISTERS_17_25_port, A2 => n338, B1 => 
                           REGISTERS_19_25_port, B2 => n321, ZN => n2933);
   U1790 : AOI22_X1 port map( A1 => REGISTERS_20_25_port, A2 => n372, B1 => 
                           REGISTERS_22_25_port, B2 => n355, ZN => n2932);
   U1791 : AOI22_X1 port map( A1 => REGISTERS_16_25_port, A2 => n406, B1 => 
                           REGISTERS_18_25_port, B2 => n389, ZN => n2931);
   U1792 : AND4_X1 port map( A1 => n2934, A2 => n2933, A3 => n2932, A4 => n2931
                           , ZN => n2951);
   U1793 : AOI22_X1 port map( A1 => REGISTERS_29_25_port, A2 => n304, B1 => 
                           REGISTERS_31_25_port, B2 => n287, ZN => n2938);
   U1794 : AOI22_X1 port map( A1 => REGISTERS_25_25_port, A2 => n338, B1 => 
                           REGISTERS_27_25_port, B2 => n321, ZN => n2937);
   U1795 : AOI22_X1 port map( A1 => REGISTERS_28_25_port, A2 => n372, B1 => 
                           REGISTERS_30_25_port, B2 => n355, ZN => n2936);
   U1796 : AOI22_X1 port map( A1 => REGISTERS_24_25_port, A2 => n406, B1 => 
                           REGISTERS_26_25_port, B2 => n389, ZN => n2935);
   U1797 : AND4_X1 port map( A1 => n2938, A2 => n2937, A3 => n2936, A4 => n2935
                           , ZN => n2950);
   U1798 : AOI22_X1 port map( A1 => REGISTERS_5_25_port, A2 => n304, B1 => 
                           REGISTERS_7_25_port, B2 => n287, ZN => n2942);
   U1799 : AOI22_X1 port map( A1 => REGISTERS_1_25_port, A2 => n338, B1 => 
                           REGISTERS_3_25_port, B2 => n321, ZN => n2941);
   U1800 : AOI22_X1 port map( A1 => REGISTERS_4_25_port, A2 => n372, B1 => 
                           REGISTERS_6_25_port, B2 => n355, ZN => n2940);
   U1801 : AOI22_X1 port map( A1 => REGISTERS_0_25_port, A2 => n406, B1 => 
                           REGISTERS_2_25_port, B2 => n389, ZN => n2939);
   U1802 : NAND4_X1 port map( A1 => n2942, A2 => n2941, A3 => n2940, A4 => 
                           n2939, ZN => n2948);
   U1803 : AOI22_X1 port map( A1 => REGISTERS_13_25_port, A2 => n304, B1 => 
                           REGISTERS_15_25_port, B2 => n287, ZN => n2946);
   U1804 : AOI22_X1 port map( A1 => REGISTERS_9_25_port, A2 => n338, B1 => 
                           REGISTERS_11_25_port, B2 => n321, ZN => n2945);
   U1805 : AOI22_X1 port map( A1 => REGISTERS_12_25_port, A2 => n372, B1 => 
                           REGISTERS_14_25_port, B2 => n355, ZN => n2944);
   U1806 : AOI22_X1 port map( A1 => REGISTERS_8_25_port, A2 => n406, B1 => 
                           REGISTERS_10_25_port, B2 => n389, ZN => n2943);
   U1807 : NAND4_X1 port map( A1 => n2946, A2 => n2945, A3 => n2944, A4 => 
                           n2943, ZN => n2947);
   U1808 : AOI22_X1 port map( A1 => n2948, A2 => n3076, B1 => n2947, B2 => 
                           n3074, ZN => n2949);
   U1809 : OAI221_X1 port map( B1 => n3080, B2 => n2951, C1 => n3078, C2 => 
                           n2950, A => n2949, ZN => N195);
   U1810 : AOI22_X1 port map( A1 => REGISTERS_21_26_port, A2 => n304, B1 => 
                           REGISTERS_23_26_port, B2 => n287, ZN => n2955);
   U1811 : AOI22_X1 port map( A1 => REGISTERS_17_26_port, A2 => n338, B1 => 
                           REGISTERS_19_26_port, B2 => n321, ZN => n2954);
   U1812 : AOI22_X1 port map( A1 => REGISTERS_20_26_port, A2 => n372, B1 => 
                           REGISTERS_22_26_port, B2 => n355, ZN => n2953);
   U1813 : AOI22_X1 port map( A1 => REGISTERS_16_26_port, A2 => n406, B1 => 
                           REGISTERS_18_26_port, B2 => n389, ZN => n2952);
   U1814 : AND4_X1 port map( A1 => n2955, A2 => n2954, A3 => n2953, A4 => n2952
                           , ZN => n2972);
   U1815 : AOI22_X1 port map( A1 => REGISTERS_29_26_port, A2 => n304, B1 => 
                           REGISTERS_31_26_port, B2 => n287, ZN => n2959);
   U1816 : AOI22_X1 port map( A1 => REGISTERS_25_26_port, A2 => n338, B1 => 
                           REGISTERS_27_26_port, B2 => n321, ZN => n2958);
   U1817 : AOI22_X1 port map( A1 => REGISTERS_28_26_port, A2 => n372, B1 => 
                           REGISTERS_30_26_port, B2 => n355, ZN => n2957);
   U1818 : AOI22_X1 port map( A1 => REGISTERS_24_26_port, A2 => n406, B1 => 
                           REGISTERS_26_26_port, B2 => n389, ZN => n2956);
   U1819 : AND4_X1 port map( A1 => n2959, A2 => n2958, A3 => n2957, A4 => n2956
                           , ZN => n2971);
   U1820 : AOI22_X1 port map( A1 => REGISTERS_5_26_port, A2 => n304, B1 => 
                           REGISTERS_7_26_port, B2 => n287, ZN => n2963);
   U1821 : AOI22_X1 port map( A1 => REGISTERS_1_26_port, A2 => n338, B1 => 
                           REGISTERS_3_26_port, B2 => n321, ZN => n2962);
   U1822 : AOI22_X1 port map( A1 => REGISTERS_4_26_port, A2 => n372, B1 => 
                           REGISTERS_6_26_port, B2 => n355, ZN => n2961);
   U1823 : AOI22_X1 port map( A1 => REGISTERS_0_26_port, A2 => n406, B1 => 
                           REGISTERS_2_26_port, B2 => n389, ZN => n2960);
   U1824 : NAND4_X1 port map( A1 => n2963, A2 => n2962, A3 => n2961, A4 => 
                           n2960, ZN => n2969);
   U1825 : AOI22_X1 port map( A1 => REGISTERS_13_26_port, A2 => n304, B1 => 
                           REGISTERS_15_26_port, B2 => n287, ZN => n2967);
   U1826 : AOI22_X1 port map( A1 => REGISTERS_9_26_port, A2 => n338, B1 => 
                           REGISTERS_11_26_port, B2 => n321, ZN => n2966);
   U1827 : AOI22_X1 port map( A1 => REGISTERS_12_26_port, A2 => n372, B1 => 
                           REGISTERS_14_26_port, B2 => n355, ZN => n2965);
   U1828 : AOI22_X1 port map( A1 => REGISTERS_8_26_port, A2 => n406, B1 => 
                           REGISTERS_10_26_port, B2 => n389, ZN => n2964);
   U1829 : NAND4_X1 port map( A1 => n2967, A2 => n2966, A3 => n2965, A4 => 
                           n2964, ZN => n2968);
   U1830 : AOI22_X1 port map( A1 => n2969, A2 => n3076, B1 => n2968, B2 => 
                           n3074, ZN => n2970);
   U1831 : OAI221_X1 port map( B1 => n3080, B2 => n2972, C1 => n3078, C2 => 
                           n2971, A => n2970, ZN => N194);
   U1832 : AOI22_X1 port map( A1 => REGISTERS_21_27_port, A2 => n305, B1 => 
                           REGISTERS_23_27_port, B2 => n288, ZN => n2976);
   U1833 : AOI22_X1 port map( A1 => REGISTERS_17_27_port, A2 => n339, B1 => 
                           REGISTERS_19_27_port, B2 => n322, ZN => n2975);
   U1834 : AOI22_X1 port map( A1 => REGISTERS_20_27_port, A2 => n373, B1 => 
                           REGISTERS_22_27_port, B2 => n356, ZN => n2974);
   U1835 : AOI22_X1 port map( A1 => REGISTERS_16_27_port, A2 => n407, B1 => 
                           REGISTERS_18_27_port, B2 => n390, ZN => n2973);
   U1836 : AND4_X1 port map( A1 => n2976, A2 => n2975, A3 => n2974, A4 => n2973
                           , ZN => n2993);
   U1837 : AOI22_X1 port map( A1 => REGISTERS_29_27_port, A2 => n305, B1 => 
                           REGISTERS_31_27_port, B2 => n288, ZN => n2980);
   U1838 : AOI22_X1 port map( A1 => REGISTERS_25_27_port, A2 => n339, B1 => 
                           REGISTERS_27_27_port, B2 => n322, ZN => n2979);
   U1839 : AOI22_X1 port map( A1 => REGISTERS_28_27_port, A2 => n373, B1 => 
                           REGISTERS_30_27_port, B2 => n356, ZN => n2978);
   U1840 : AOI22_X1 port map( A1 => REGISTERS_24_27_port, A2 => n407, B1 => 
                           REGISTERS_26_27_port, B2 => n390, ZN => n2977);
   U1841 : AND4_X1 port map( A1 => n2980, A2 => n2979, A3 => n2978, A4 => n2977
                           , ZN => n2992);
   U1842 : AOI22_X1 port map( A1 => REGISTERS_5_27_port, A2 => n305, B1 => 
                           REGISTERS_7_27_port, B2 => n288, ZN => n2984);
   U1843 : AOI22_X1 port map( A1 => REGISTERS_1_27_port, A2 => n339, B1 => 
                           REGISTERS_3_27_port, B2 => n322, ZN => n2983);
   U1844 : AOI22_X1 port map( A1 => REGISTERS_4_27_port, A2 => n373, B1 => 
                           REGISTERS_6_27_port, B2 => n356, ZN => n2982);
   U1845 : AOI22_X1 port map( A1 => REGISTERS_0_27_port, A2 => n407, B1 => 
                           REGISTERS_2_27_port, B2 => n390, ZN => n2981);
   U1846 : NAND4_X1 port map( A1 => n2984, A2 => n2983, A3 => n2982, A4 => 
                           n2981, ZN => n2990);
   U1847 : AOI22_X1 port map( A1 => REGISTERS_13_27_port, A2 => n305, B1 => 
                           REGISTERS_15_27_port, B2 => n288, ZN => n2988);
   U1848 : AOI22_X1 port map( A1 => REGISTERS_9_27_port, A2 => n339, B1 => 
                           REGISTERS_11_27_port, B2 => n322, ZN => n2987);
   U1849 : AOI22_X1 port map( A1 => REGISTERS_12_27_port, A2 => n373, B1 => 
                           REGISTERS_14_27_port, B2 => n356, ZN => n2986);
   U1850 : AOI22_X1 port map( A1 => REGISTERS_8_27_port, A2 => n407, B1 => 
                           REGISTERS_10_27_port, B2 => n390, ZN => n2985);
   U1851 : NAND4_X1 port map( A1 => n2988, A2 => n2987, A3 => n2986, A4 => 
                           n2985, ZN => n2989);
   U1852 : AOI22_X1 port map( A1 => n2990, A2 => n3076, B1 => n2989, B2 => 
                           n3074, ZN => n2991);
   U1853 : OAI221_X1 port map( B1 => n3080, B2 => n2993, C1 => n3078, C2 => 
                           n2992, A => n2991, ZN => N193);
   U1854 : AOI22_X1 port map( A1 => REGISTERS_21_28_port, A2 => n305, B1 => 
                           REGISTERS_23_28_port, B2 => n288, ZN => n2997);
   U1855 : AOI22_X1 port map( A1 => REGISTERS_17_28_port, A2 => n339, B1 => 
                           REGISTERS_19_28_port, B2 => n322, ZN => n2996);
   U1856 : AOI22_X1 port map( A1 => REGISTERS_20_28_port, A2 => n373, B1 => 
                           REGISTERS_22_28_port, B2 => n356, ZN => n2995);
   U1857 : AOI22_X1 port map( A1 => REGISTERS_16_28_port, A2 => n407, B1 => 
                           REGISTERS_18_28_port, B2 => n390, ZN => n2994);
   U1858 : AND4_X1 port map( A1 => n2997, A2 => n2996, A3 => n2995, A4 => n2994
                           , ZN => n3014);
   U1859 : AOI22_X1 port map( A1 => REGISTERS_29_28_port, A2 => n305, B1 => 
                           REGISTERS_31_28_port, B2 => n288, ZN => n3001);
   U1860 : AOI22_X1 port map( A1 => REGISTERS_25_28_port, A2 => n339, B1 => 
                           REGISTERS_27_28_port, B2 => n322, ZN => n3000);
   U1861 : AOI22_X1 port map( A1 => REGISTERS_28_28_port, A2 => n373, B1 => 
                           REGISTERS_30_28_port, B2 => n356, ZN => n2999);
   U1862 : AOI22_X1 port map( A1 => REGISTERS_24_28_port, A2 => n407, B1 => 
                           REGISTERS_26_28_port, B2 => n390, ZN => n2998);
   U1863 : AND4_X1 port map( A1 => n3001, A2 => n3000, A3 => n2999, A4 => n2998
                           , ZN => n3013);
   U1864 : AOI22_X1 port map( A1 => REGISTERS_5_28_port, A2 => n305, B1 => 
                           REGISTERS_7_28_port, B2 => n288, ZN => n3005);
   U1865 : AOI22_X1 port map( A1 => REGISTERS_1_28_port, A2 => n339, B1 => 
                           REGISTERS_3_28_port, B2 => n322, ZN => n3004);
   U1866 : AOI22_X1 port map( A1 => REGISTERS_4_28_port, A2 => n373, B1 => 
                           REGISTERS_6_28_port, B2 => n356, ZN => n3003);
   U1867 : AOI22_X1 port map( A1 => REGISTERS_0_28_port, A2 => n407, B1 => 
                           REGISTERS_2_28_port, B2 => n390, ZN => n3002);
   U1868 : NAND4_X1 port map( A1 => n3005, A2 => n3004, A3 => n3003, A4 => 
                           n3002, ZN => n3011);
   U1869 : AOI22_X1 port map( A1 => REGISTERS_13_28_port, A2 => n305, B1 => 
                           REGISTERS_15_28_port, B2 => n288, ZN => n3009);
   U1870 : AOI22_X1 port map( A1 => REGISTERS_9_28_port, A2 => n339, B1 => 
                           REGISTERS_11_28_port, B2 => n322, ZN => n3008);
   U1871 : AOI22_X1 port map( A1 => REGISTERS_12_28_port, A2 => n373, B1 => 
                           REGISTERS_14_28_port, B2 => n356, ZN => n3007);
   U1872 : AOI22_X1 port map( A1 => REGISTERS_8_28_port, A2 => n407, B1 => 
                           REGISTERS_10_28_port, B2 => n390, ZN => n3006);
   U1873 : NAND4_X1 port map( A1 => n3009, A2 => n3008, A3 => n3007, A4 => 
                           n3006, ZN => n3010);
   U1874 : AOI22_X1 port map( A1 => n3011, A2 => n3076, B1 => n3010, B2 => 
                           n3074, ZN => n3012);
   U1875 : OAI221_X1 port map( B1 => n3080, B2 => n3014, C1 => n3078, C2 => 
                           n3013, A => n3012, ZN => N192);
   U1876 : AOI22_X1 port map( A1 => REGISTERS_21_29_port, A2 => n305, B1 => 
                           REGISTERS_23_29_port, B2 => n288, ZN => n3018);
   U1877 : AOI22_X1 port map( A1 => REGISTERS_17_29_port, A2 => n339, B1 => 
                           REGISTERS_19_29_port, B2 => n322, ZN => n3017);
   U1878 : AOI22_X1 port map( A1 => REGISTERS_20_29_port, A2 => n373, B1 => 
                           REGISTERS_22_29_port, B2 => n356, ZN => n3016);
   U1879 : AOI22_X1 port map( A1 => REGISTERS_16_29_port, A2 => n407, B1 => 
                           REGISTERS_18_29_port, B2 => n390, ZN => n3015);
   U1880 : AND4_X1 port map( A1 => n3018, A2 => n3017, A3 => n3016, A4 => n3015
                           , ZN => n3035);
   U1881 : AOI22_X1 port map( A1 => REGISTERS_29_29_port, A2 => n305, B1 => 
                           REGISTERS_31_29_port, B2 => n288, ZN => n3022);
   U1882 : AOI22_X1 port map( A1 => REGISTERS_25_29_port, A2 => n339, B1 => 
                           REGISTERS_27_29_port, B2 => n322, ZN => n3021);
   U1883 : AOI22_X1 port map( A1 => REGISTERS_28_29_port, A2 => n373, B1 => 
                           REGISTERS_30_29_port, B2 => n356, ZN => n3020);
   U1884 : AOI22_X1 port map( A1 => REGISTERS_24_29_port, A2 => n407, B1 => 
                           REGISTERS_26_29_port, B2 => n390, ZN => n3019);
   U1885 : AND4_X1 port map( A1 => n3022, A2 => n3021, A3 => n3020, A4 => n3019
                           , ZN => n3034);
   U1886 : AOI22_X1 port map( A1 => REGISTERS_5_29_port, A2 => n305, B1 => 
                           REGISTERS_7_29_port, B2 => n288, ZN => n3026);
   U1887 : AOI22_X1 port map( A1 => REGISTERS_1_29_port, A2 => n339, B1 => 
                           REGISTERS_3_29_port, B2 => n322, ZN => n3025);
   U1888 : AOI22_X1 port map( A1 => REGISTERS_4_29_port, A2 => n373, B1 => 
                           REGISTERS_6_29_port, B2 => n356, ZN => n3024);
   U1889 : AOI22_X1 port map( A1 => REGISTERS_0_29_port, A2 => n407, B1 => 
                           REGISTERS_2_29_port, B2 => n390, ZN => n3023);
   U1890 : NAND4_X1 port map( A1 => n3026, A2 => n3025, A3 => n3024, A4 => 
                           n3023, ZN => n3032);
   U1891 : AOI22_X1 port map( A1 => REGISTERS_13_29_port, A2 => n305, B1 => 
                           REGISTERS_15_29_port, B2 => n288, ZN => n3030);
   U1892 : AOI22_X1 port map( A1 => REGISTERS_9_29_port, A2 => n339, B1 => 
                           REGISTERS_11_29_port, B2 => n322, ZN => n3029);
   U1893 : AOI22_X1 port map( A1 => REGISTERS_12_29_port, A2 => n373, B1 => 
                           REGISTERS_14_29_port, B2 => n356, ZN => n3028);
   U1894 : AOI22_X1 port map( A1 => REGISTERS_8_29_port, A2 => n407, B1 => 
                           REGISTERS_10_29_port, B2 => n390, ZN => n3027);
   U1895 : NAND4_X1 port map( A1 => n3030, A2 => n3029, A3 => n3028, A4 => 
                           n3027, ZN => n3031);
   U1896 : AOI22_X1 port map( A1 => n3032, A2 => n3076, B1 => n3031, B2 => 
                           n3074, ZN => n3033);
   U1897 : OAI221_X1 port map( B1 => n3080, B2 => n3035, C1 => n3078, C2 => 
                           n3034, A => n3033, ZN => N191);
   U1898 : AOI22_X1 port map( A1 => REGISTERS_21_30_port, A2 => n306, B1 => 
                           REGISTERS_23_30_port, B2 => n289, ZN => n3039);
   U1899 : AOI22_X1 port map( A1 => REGISTERS_17_30_port, A2 => n340, B1 => 
                           REGISTERS_19_30_port, B2 => n323, ZN => n3038);
   U1900 : AOI22_X1 port map( A1 => REGISTERS_20_30_port, A2 => n374, B1 => 
                           REGISTERS_22_30_port, B2 => n357, ZN => n3037);
   U1901 : AOI22_X1 port map( A1 => REGISTERS_16_30_port, A2 => n408, B1 => 
                           REGISTERS_18_30_port, B2 => n391, ZN => n3036);
   U1902 : AND4_X1 port map( A1 => n3039, A2 => n3038, A3 => n3037, A4 => n3036
                           , ZN => n3056);
   U1903 : AOI22_X1 port map( A1 => REGISTERS_29_30_port, A2 => n306, B1 => 
                           REGISTERS_31_30_port, B2 => n289, ZN => n3043);
   U1904 : AOI22_X1 port map( A1 => REGISTERS_25_30_port, A2 => n340, B1 => 
                           REGISTERS_27_30_port, B2 => n323, ZN => n3042);
   U1905 : AOI22_X1 port map( A1 => REGISTERS_28_30_port, A2 => n374, B1 => 
                           REGISTERS_30_30_port, B2 => n357, ZN => n3041);
   U1906 : AOI22_X1 port map( A1 => REGISTERS_24_30_port, A2 => n408, B1 => 
                           REGISTERS_26_30_port, B2 => n391, ZN => n3040);
   U1907 : AND4_X1 port map( A1 => n3043, A2 => n3042, A3 => n3041, A4 => n3040
                           , ZN => n3055);
   U1908 : AOI22_X1 port map( A1 => REGISTERS_5_30_port, A2 => n306, B1 => 
                           REGISTERS_7_30_port, B2 => n289, ZN => n3047);
   U1909 : AOI22_X1 port map( A1 => REGISTERS_1_30_port, A2 => n340, B1 => 
                           REGISTERS_3_30_port, B2 => n323, ZN => n3046);
   U1910 : AOI22_X1 port map( A1 => REGISTERS_4_30_port, A2 => n374, B1 => 
                           REGISTERS_6_30_port, B2 => n357, ZN => n3045);
   U1911 : AOI22_X1 port map( A1 => REGISTERS_0_30_port, A2 => n408, B1 => 
                           REGISTERS_2_30_port, B2 => n391, ZN => n3044);
   U1912 : NAND4_X1 port map( A1 => n3047, A2 => n3046, A3 => n3045, A4 => 
                           n3044, ZN => n3053);
   U1913 : AOI22_X1 port map( A1 => REGISTERS_13_30_port, A2 => n306, B1 => 
                           REGISTERS_15_30_port, B2 => n289, ZN => n3051);
   U1914 : AOI22_X1 port map( A1 => REGISTERS_9_30_port, A2 => n340, B1 => 
                           REGISTERS_11_30_port, B2 => n323, ZN => n3050);
   U1915 : AOI22_X1 port map( A1 => REGISTERS_12_30_port, A2 => n374, B1 => 
                           REGISTERS_14_30_port, B2 => n357, ZN => n3049);
   U1916 : AOI22_X1 port map( A1 => REGISTERS_8_30_port, A2 => n408, B1 => 
                           REGISTERS_10_30_port, B2 => n391, ZN => n3048);
   U1917 : NAND4_X1 port map( A1 => n3051, A2 => n3050, A3 => n3049, A4 => 
                           n3048, ZN => n3052);
   U1918 : AOI22_X1 port map( A1 => n3053, A2 => n3076, B1 => n3052, B2 => 
                           n3074, ZN => n3054);
   U1919 : OAI221_X1 port map( B1 => n3080, B2 => n3056, C1 => n3078, C2 => 
                           n3055, A => n3054, ZN => N190);
   U1920 : AOI22_X1 port map( A1 => REGISTERS_21_31_port, A2 => n306, B1 => 
                           REGISTERS_23_31_port, B2 => n289, ZN => n3060);
   U1921 : AOI22_X1 port map( A1 => REGISTERS_17_31_port, A2 => n340, B1 => 
                           REGISTERS_19_31_port, B2 => n323, ZN => n3059);
   U1922 : AOI22_X1 port map( A1 => REGISTERS_20_31_port, A2 => n374, B1 => 
                           REGISTERS_22_31_port, B2 => n357, ZN => n3058);
   U1923 : AOI22_X1 port map( A1 => REGISTERS_16_31_port, A2 => n408, B1 => 
                           REGISTERS_18_31_port, B2 => n391, ZN => n3057);
   U1924 : AND4_X1 port map( A1 => n3060, A2 => n3059, A3 => n3058, A4 => n3057
                           , ZN => n3081);
   U1925 : AOI22_X1 port map( A1 => REGISTERS_29_31_port, A2 => n306, B1 => 
                           REGISTERS_31_31_port, B2 => n289, ZN => n3064);
   U1926 : AOI22_X1 port map( A1 => REGISTERS_25_31_port, A2 => n340, B1 => 
                           REGISTERS_27_31_port, B2 => n323, ZN => n3063);
   U1927 : AOI22_X1 port map( A1 => REGISTERS_28_31_port, A2 => n374, B1 => 
                           REGISTERS_30_31_port, B2 => n357, ZN => n3062);
   U1928 : AOI22_X1 port map( A1 => REGISTERS_24_31_port, A2 => n408, B1 => 
                           REGISTERS_26_31_port, B2 => n391, ZN => n3061);
   U1929 : AND4_X1 port map( A1 => n3064, A2 => n3063, A3 => n3062, A4 => n3061
                           , ZN => n3079);
   U1930 : AOI22_X1 port map( A1 => REGISTERS_5_31_port, A2 => n306, B1 => 
                           REGISTERS_7_31_port, B2 => n289, ZN => n3068);
   U1931 : AOI22_X1 port map( A1 => REGISTERS_1_31_port, A2 => n340, B1 => 
                           REGISTERS_3_31_port, B2 => n323, ZN => n3067);
   U1932 : AOI22_X1 port map( A1 => REGISTERS_4_31_port, A2 => n374, B1 => 
                           REGISTERS_6_31_port, B2 => n357, ZN => n3066);
   U1933 : AOI22_X1 port map( A1 => REGISTERS_0_31_port, A2 => n408, B1 => 
                           REGISTERS_2_31_port, B2 => n391, ZN => n3065);
   U1934 : NAND4_X1 port map( A1 => n3068, A2 => n3067, A3 => n3066, A4 => 
                           n3065, ZN => n3075);
   U1935 : AOI22_X1 port map( A1 => REGISTERS_13_31_port, A2 => n306, B1 => 
                           REGISTERS_15_31_port, B2 => n289, ZN => n3072);
   U1936 : AOI22_X1 port map( A1 => REGISTERS_9_31_port, A2 => n340, B1 => 
                           REGISTERS_11_31_port, B2 => n323, ZN => n3071);
   U1937 : AOI22_X1 port map( A1 => REGISTERS_12_31_port, A2 => n374, B1 => 
                           REGISTERS_14_31_port, B2 => n357, ZN => n3070);
   U1938 : AOI22_X1 port map( A1 => REGISTERS_8_31_port, A2 => n408, B1 => 
                           REGISTERS_10_31_port, B2 => n391, ZN => n3069);
   U1939 : NAND4_X1 port map( A1 => n3072, A2 => n3071, A3 => n3070, A4 => 
                           n3069, ZN => n3073);
   U1940 : AOI22_X1 port map( A1 => n3076, A2 => n3075, B1 => n3074, B2 => 
                           n3073, ZN => n3077);
   U1941 : OAI221_X1 port map( B1 => n3081, B2 => n3080, C1 => n3079, C2 => 
                           n3078, A => n3077, ZN => N189);
   U1942 : OAI21_X1 port map( B1 => n3086, B2 => n17, A => n3087, ZN => n2614);
   U1943 : OAI21_X1 port map( B1 => n3086, B2 => n18, A => n3087, ZN => n2613);
   U1944 : OAI21_X1 port map( B1 => n3086, B2 => n19, A => n3087, ZN => n2612);
   U1945 : OAI21_X1 port map( B1 => n3086, B2 => n20, A => n3087, ZN => n2611);
   U1946 : OAI21_X1 port map( B1 => n3086, B2 => n21, A => n3087, ZN => n2610);
   U1947 : OAI21_X1 port map( B1 => n3086, B2 => n22, A => n3087, ZN => n2609);
   U1948 : OAI21_X1 port map( B1 => n3086, B2 => n23, A => n3087, ZN => n2608);
   U1949 : OAI21_X1 port map( B1 => n3086, B2 => n24, A => n3087, ZN => n2607);
   U1950 : OAI21_X1 port map( B1 => n3086, B2 => n25, A => n3087, ZN => n2606);
   U1951 : OAI21_X1 port map( B1 => n3086, B2 => n26, A => n3087, ZN => n2605);
   U1952 : OAI21_X1 port map( B1 => n3086, B2 => n27, A => n3087, ZN => n2604);
   U1953 : OAI21_X1 port map( B1 => n3086, B2 => n28, A => n3087, ZN => n2603);
   U1954 : OAI21_X1 port map( B1 => n3086, B2 => n29, A => n3087, ZN => n2602);
   U1955 : OAI21_X1 port map( B1 => n3086, B2 => n30, A => n3087, ZN => n2601);
   U1956 : OAI21_X1 port map( B1 => n3086, B2 => n31, A => n3087, ZN => n2600);
   U1957 : OAI21_X1 port map( B1 => n3086, B2 => n32, A => n3087, ZN => n2599);
   U1958 : OAI21_X1 port map( B1 => n3086, B2 => n33, A => n3087, ZN => n2598);
   U1959 : OAI21_X1 port map( B1 => n3086, B2 => n34, A => n3087, ZN => n2597);
   U1960 : OAI21_X1 port map( B1 => n3086, B2 => n35, A => n3087, ZN => n2596);
   U1961 : OAI21_X1 port map( B1 => n3086, B2 => n36, A => n3087, ZN => n2595);
   U1962 : OAI21_X1 port map( B1 => n3086, B2 => n37, A => n3087, ZN => n2594);
   U1963 : OAI21_X1 port map( B1 => n3086, B2 => n38, A => n3087, ZN => n2593);
   U1964 : OAI21_X1 port map( B1 => n3086, B2 => n39, A => n3087, ZN => n2592);
   U1965 : OAI21_X1 port map( B1 => n3086, B2 => n40, A => n3087, ZN => n2591);
   U1966 : OAI21_X1 port map( B1 => n3086, B2 => n41, A => n3087, ZN => n2590);
   U1967 : OAI21_X1 port map( B1 => n3086, B2 => n42, A => n3087, ZN => n2589);
   U1968 : OAI21_X1 port map( B1 => n3086, B2 => n43, A => n3087, ZN => n2588);
   U1969 : OAI21_X1 port map( B1 => n3086, B2 => n44, A => n3087, ZN => n2587);
   U1970 : OAI21_X1 port map( B1 => n3086, B2 => n45, A => n3087, ZN => n2586);
   U1971 : OAI21_X1 port map( B1 => n3086, B2 => n46, A => n3087, ZN => n2585);
   U1972 : OAI21_X1 port map( B1 => n3086, B2 => n47, A => n3087, ZN => n2584);
   U1973 : OAI21_X1 port map( B1 => n3086, B2 => n48, A => n3087, ZN => n2583);
   U1974 : MUX2_X1 port map( A => REGISTERS_0_31_port, B => n3089, S => n3090, 
                           Z => n2582);
   U1975 : MUX2_X1 port map( A => REGISTERS_0_30_port, B => n3091, S => n3090, 
                           Z => n2581);
   U1976 : MUX2_X1 port map( A => REGISTERS_0_29_port, B => n3092, S => n3090, 
                           Z => n2580);
   U1977 : MUX2_X1 port map( A => REGISTERS_0_28_port, B => n3093, S => n3090, 
                           Z => n2579);
   U1978 : MUX2_X1 port map( A => REGISTERS_0_27_port, B => n3094, S => n3090, 
                           Z => n2578);
   U1979 : MUX2_X1 port map( A => REGISTERS_0_26_port, B => n3095, S => n3090, 
                           Z => n2577);
   U1980 : MUX2_X1 port map( A => REGISTERS_0_25_port, B => n3096, S => n3090, 
                           Z => n2576);
   U1981 : MUX2_X1 port map( A => REGISTERS_0_24_port, B => n3097, S => n3090, 
                           Z => n2575);
   U1982 : MUX2_X1 port map( A => REGISTERS_0_23_port, B => n3098, S => n3090, 
                           Z => n2574);
   U1983 : MUX2_X1 port map( A => REGISTERS_0_22_port, B => n3099, S => n3090, 
                           Z => n2573);
   U1984 : MUX2_X1 port map( A => REGISTERS_0_21_port, B => n3100, S => n3090, 
                           Z => n2572);
   U1985 : MUX2_X1 port map( A => REGISTERS_0_20_port, B => n3101, S => n3090, 
                           Z => n2571);
   U1986 : MUX2_X1 port map( A => REGISTERS_0_19_port, B => n3102, S => n3090, 
                           Z => n2570);
   U1987 : MUX2_X1 port map( A => REGISTERS_0_18_port, B => n3103, S => n3090, 
                           Z => n2569);
   U1988 : MUX2_X1 port map( A => REGISTERS_0_17_port, B => n3104, S => n3090, 
                           Z => n2568);
   U1989 : MUX2_X1 port map( A => REGISTERS_0_16_port, B => n3105, S => n3090, 
                           Z => n2567);
   U1990 : MUX2_X1 port map( A => REGISTERS_0_15_port, B => n3106, S => n3090, 
                           Z => n2566);
   U1991 : MUX2_X1 port map( A => REGISTERS_0_14_port, B => n3107, S => n3090, 
                           Z => n2565);
   U1992 : MUX2_X1 port map( A => REGISTERS_0_13_port, B => n3108, S => n3090, 
                           Z => n2564);
   U1993 : MUX2_X1 port map( A => REGISTERS_0_12_port, B => n3109, S => n3090, 
                           Z => n2563);
   U1994 : MUX2_X1 port map( A => REGISTERS_0_11_port, B => n3110, S => n3090, 
                           Z => n2562);
   U1995 : MUX2_X1 port map( A => REGISTERS_0_10_port, B => n3111, S => n3090, 
                           Z => n2561);
   U1996 : MUX2_X1 port map( A => REGISTERS_0_9_port, B => n3112, S => n3090, Z
                           => n2560);
   U1997 : MUX2_X1 port map( A => REGISTERS_0_8_port, B => n3113, S => n3090, Z
                           => n2559);
   U1998 : MUX2_X1 port map( A => REGISTERS_0_7_port, B => n3114, S => n3090, Z
                           => n2558);
   U1999 : MUX2_X1 port map( A => REGISTERS_0_6_port, B => n3115, S => n3090, Z
                           => n2557);
   U2000 : MUX2_X1 port map( A => REGISTERS_0_5_port, B => n3116, S => n3090, Z
                           => n2556);
   U2001 : MUX2_X1 port map( A => REGISTERS_0_4_port, B => n3117, S => n3090, Z
                           => n2555);
   U2002 : MUX2_X1 port map( A => REGISTERS_0_3_port, B => n3118, S => n3090, Z
                           => n2554);
   U2003 : MUX2_X1 port map( A => REGISTERS_0_2_port, B => n3119, S => n3090, Z
                           => n2553);
   U2004 : MUX2_X1 port map( A => REGISTERS_0_1_port, B => n3120, S => n3090, Z
                           => n2552);
   U2005 : MUX2_X1 port map( A => REGISTERS_0_0_port, B => n3121, S => n3090, Z
                           => n2551);
   U2006 : MUX2_X1 port map( A => REGISTERS_1_31_port, B => n3089, S => n140, Z
                           => n2550);
   U2007 : MUX2_X1 port map( A => REGISTERS_1_30_port, B => n3091, S => n140, Z
                           => n2549);
   U2008 : MUX2_X1 port map( A => REGISTERS_1_29_port, B => n3092, S => n140, Z
                           => n2548);
   U2009 : MUX2_X1 port map( A => REGISTERS_1_28_port, B => n3093, S => n140, Z
                           => n2547);
   U2010 : MUX2_X1 port map( A => REGISTERS_1_27_port, B => n3094, S => n140, Z
                           => n2546);
   U2011 : MUX2_X1 port map( A => REGISTERS_1_26_port, B => n3095, S => n140, Z
                           => n2545);
   U2012 : MUX2_X1 port map( A => REGISTERS_1_25_port, B => n3096, S => n140, Z
                           => n2544);
   U2013 : MUX2_X1 port map( A => REGISTERS_1_24_port, B => n3097, S => n140, Z
                           => n2543);
   U2014 : MUX2_X1 port map( A => REGISTERS_1_23_port, B => n3098, S => n140, Z
                           => n2542);
   U2015 : MUX2_X1 port map( A => REGISTERS_1_22_port, B => n3099, S => n140, Z
                           => n2541);
   U2016 : MUX2_X1 port map( A => REGISTERS_1_21_port, B => n3100, S => n140, Z
                           => n2540);
   U2017 : MUX2_X1 port map( A => REGISTERS_1_20_port, B => n3101, S => n140, Z
                           => n2539);
   U2018 : MUX2_X1 port map( A => REGISTERS_1_19_port, B => n3102, S => n140, Z
                           => n2538);
   U2019 : MUX2_X1 port map( A => REGISTERS_1_18_port, B => n3103, S => n140, Z
                           => n2537);
   U2020 : MUX2_X1 port map( A => REGISTERS_1_17_port, B => n3104, S => n140, Z
                           => n2536);
   U2021 : MUX2_X1 port map( A => REGISTERS_1_16_port, B => n3105, S => n140, Z
                           => n2535);
   U2022 : MUX2_X1 port map( A => REGISTERS_1_15_port, B => n3106, S => n140, Z
                           => n2534);
   U2023 : MUX2_X1 port map( A => REGISTERS_1_14_port, B => n3107, S => n140, Z
                           => n2533);
   U2024 : MUX2_X1 port map( A => REGISTERS_1_13_port, B => n3108, S => n140, Z
                           => n2532);
   U2025 : MUX2_X1 port map( A => REGISTERS_1_12_port, B => n3109, S => n140, Z
                           => n2531);
   U2026 : MUX2_X1 port map( A => REGISTERS_1_11_port, B => n3110, S => n140, Z
                           => n2530);
   U2027 : MUX2_X1 port map( A => REGISTERS_1_10_port, B => n3111, S => n140, Z
                           => n2529);
   U2028 : MUX2_X1 port map( A => REGISTERS_1_9_port, B => n3112, S => n140, Z 
                           => n2528);
   U2029 : MUX2_X1 port map( A => REGISTERS_1_8_port, B => n3113, S => n140, Z 
                           => n2527);
   U2030 : MUX2_X1 port map( A => REGISTERS_1_7_port, B => n3114, S => n140, Z 
                           => n2526);
   U2031 : MUX2_X1 port map( A => REGISTERS_1_6_port, B => n3115, S => n140, Z 
                           => n2525);
   U2032 : MUX2_X1 port map( A => REGISTERS_1_5_port, B => n3116, S => n140, Z 
                           => n2524);
   U2033 : MUX2_X1 port map( A => REGISTERS_1_4_port, B => n3117, S => n140, Z 
                           => n2523);
   U2034 : MUX2_X1 port map( A => REGISTERS_1_3_port, B => n3118, S => n140, Z 
                           => n2522);
   U2035 : MUX2_X1 port map( A => REGISTERS_1_2_port, B => n3119, S => n140, Z 
                           => n2521);
   U2036 : MUX2_X1 port map( A => REGISTERS_1_1_port, B => n3120, S => n140, Z 
                           => n2520);
   U2037 : MUX2_X1 port map( A => REGISTERS_1_0_port, B => n3121, S => n140, Z 
                           => n2519);
   U2038 : OAI21_X1 port map( B1 => n3122, B2 => n3126, A => n3124, ZN => n3125
                           );
   U2039 : MUX2_X1 port map( A => REGISTERS_2_31_port, B => n3089, S => n142, Z
                           => n2518);
   U2040 : MUX2_X1 port map( A => REGISTERS_2_30_port, B => n3091, S => n142, Z
                           => n2517);
   U2041 : MUX2_X1 port map( A => REGISTERS_2_29_port, B => n3092, S => n142, Z
                           => n2516);
   U2042 : MUX2_X1 port map( A => REGISTERS_2_28_port, B => n3093, S => n142, Z
                           => n2515);
   U2043 : MUX2_X1 port map( A => REGISTERS_2_27_port, B => n3094, S => n142, Z
                           => n2514);
   U2044 : MUX2_X1 port map( A => REGISTERS_2_26_port, B => n3095, S => n142, Z
                           => n2513);
   U2045 : MUX2_X1 port map( A => REGISTERS_2_25_port, B => n3096, S => n142, Z
                           => n2512);
   U2046 : MUX2_X1 port map( A => REGISTERS_2_24_port, B => n3097, S => n142, Z
                           => n2511);
   U2047 : MUX2_X1 port map( A => REGISTERS_2_23_port, B => n3098, S => n142, Z
                           => n2510);
   U2048 : MUX2_X1 port map( A => REGISTERS_2_22_port, B => n3099, S => n142, Z
                           => n2509);
   U2049 : MUX2_X1 port map( A => REGISTERS_2_21_port, B => n3100, S => n142, Z
                           => n2508);
   U2050 : MUX2_X1 port map( A => REGISTERS_2_20_port, B => n3101, S => n142, Z
                           => n2507);
   U2051 : MUX2_X1 port map( A => REGISTERS_2_19_port, B => n3102, S => n142, Z
                           => n2506);
   U2052 : MUX2_X1 port map( A => REGISTERS_2_18_port, B => n3103, S => n142, Z
                           => n2505);
   U2053 : MUX2_X1 port map( A => REGISTERS_2_17_port, B => n3104, S => n142, Z
                           => n2504);
   U2054 : MUX2_X1 port map( A => REGISTERS_2_16_port, B => n3105, S => n142, Z
                           => n2503);
   U2055 : MUX2_X1 port map( A => REGISTERS_2_15_port, B => n3106, S => n142, Z
                           => n2502);
   U2056 : MUX2_X1 port map( A => REGISTERS_2_14_port, B => n3107, S => n142, Z
                           => n2501);
   U2057 : MUX2_X1 port map( A => REGISTERS_2_13_port, B => n3108, S => n142, Z
                           => n2500);
   U2058 : MUX2_X1 port map( A => REGISTERS_2_12_port, B => n3109, S => n142, Z
                           => n2499);
   U2059 : MUX2_X1 port map( A => REGISTERS_2_11_port, B => n3110, S => n142, Z
                           => n2498);
   U2060 : MUX2_X1 port map( A => REGISTERS_2_10_port, B => n3111, S => n142, Z
                           => n2497);
   U2061 : MUX2_X1 port map( A => REGISTERS_2_9_port, B => n3112, S => n142, Z 
                           => n2496);
   U2062 : MUX2_X1 port map( A => REGISTERS_2_8_port, B => n3113, S => n142, Z 
                           => n2495);
   U2063 : MUX2_X1 port map( A => REGISTERS_2_7_port, B => n3114, S => n142, Z 
                           => n2494);
   U2064 : MUX2_X1 port map( A => REGISTERS_2_6_port, B => n3115, S => n142, Z 
                           => n2493);
   U2065 : MUX2_X1 port map( A => REGISTERS_2_5_port, B => n3116, S => n142, Z 
                           => n2492);
   U2066 : MUX2_X1 port map( A => REGISTERS_2_4_port, B => n3117, S => n142, Z 
                           => n2491);
   U2067 : MUX2_X1 port map( A => REGISTERS_2_3_port, B => n3118, S => n142, Z 
                           => n2490);
   U2068 : MUX2_X1 port map( A => REGISTERS_2_2_port, B => n3119, S => n142, Z 
                           => n2489);
   U2069 : MUX2_X1 port map( A => REGISTERS_2_1_port, B => n3120, S => n142, Z 
                           => n2488);
   U2070 : MUX2_X1 port map( A => REGISTERS_2_0_port, B => n3121, S => n142, Z 
                           => n2487);
   U2071 : OAI21_X1 port map( B1 => n3122, B2 => n3128, A => n3124, ZN => n3127
                           );
   U2072 : MUX2_X1 port map( A => REGISTERS_3_31_port, B => n3089, S => n136, Z
                           => n2486);
   U2073 : MUX2_X1 port map( A => REGISTERS_3_30_port, B => n3091, S => n136, Z
                           => n2485);
   U2074 : MUX2_X1 port map( A => REGISTERS_3_29_port, B => n3092, S => n136, Z
                           => n2484);
   U2075 : MUX2_X1 port map( A => REGISTERS_3_28_port, B => n3093, S => n136, Z
                           => n2483);
   U2076 : MUX2_X1 port map( A => REGISTERS_3_27_port, B => n3094, S => n136, Z
                           => n2482);
   U2077 : MUX2_X1 port map( A => REGISTERS_3_26_port, B => n3095, S => n136, Z
                           => n2481);
   U2078 : MUX2_X1 port map( A => REGISTERS_3_25_port, B => n3096, S => n136, Z
                           => n2480);
   U2079 : MUX2_X1 port map( A => REGISTERS_3_24_port, B => n3097, S => n136, Z
                           => n2479);
   U2080 : MUX2_X1 port map( A => REGISTERS_3_23_port, B => n3098, S => n136, Z
                           => n2478);
   U2081 : MUX2_X1 port map( A => REGISTERS_3_22_port, B => n3099, S => n136, Z
                           => n2477);
   U2082 : MUX2_X1 port map( A => REGISTERS_3_21_port, B => n3100, S => n136, Z
                           => n2476);
   U2083 : MUX2_X1 port map( A => REGISTERS_3_20_port, B => n3101, S => n136, Z
                           => n2475);
   U2084 : MUX2_X1 port map( A => REGISTERS_3_19_port, B => n3102, S => n136, Z
                           => n2474);
   U2085 : MUX2_X1 port map( A => REGISTERS_3_18_port, B => n3103, S => n136, Z
                           => n2473);
   U2086 : MUX2_X1 port map( A => REGISTERS_3_17_port, B => n3104, S => n136, Z
                           => n2472);
   U2087 : MUX2_X1 port map( A => REGISTERS_3_16_port, B => n3105, S => n136, Z
                           => n2471);
   U2088 : MUX2_X1 port map( A => REGISTERS_3_15_port, B => n3106, S => n136, Z
                           => n2470);
   U2089 : MUX2_X1 port map( A => REGISTERS_3_14_port, B => n3107, S => n136, Z
                           => n2469);
   U2090 : MUX2_X1 port map( A => REGISTERS_3_13_port, B => n3108, S => n136, Z
                           => n2468);
   U2091 : MUX2_X1 port map( A => REGISTERS_3_12_port, B => n3109, S => n136, Z
                           => n2467);
   U2092 : MUX2_X1 port map( A => REGISTERS_3_11_port, B => n3110, S => n136, Z
                           => n2466);
   U2093 : MUX2_X1 port map( A => REGISTERS_3_10_port, B => n3111, S => n136, Z
                           => n2465);
   U2094 : MUX2_X1 port map( A => REGISTERS_3_9_port, B => n3112, S => n136, Z 
                           => n2464);
   U2095 : MUX2_X1 port map( A => REGISTERS_3_8_port, B => n3113, S => n136, Z 
                           => n2463);
   U2096 : MUX2_X1 port map( A => REGISTERS_3_7_port, B => n3114, S => n136, Z 
                           => n2462);
   U2097 : MUX2_X1 port map( A => REGISTERS_3_6_port, B => n3115, S => n136, Z 
                           => n2461);
   U2098 : MUX2_X1 port map( A => REGISTERS_3_5_port, B => n3116, S => n136, Z 
                           => n2460);
   U2099 : MUX2_X1 port map( A => REGISTERS_3_4_port, B => n3117, S => n136, Z 
                           => n2459);
   U2100 : MUX2_X1 port map( A => REGISTERS_3_3_port, B => n3118, S => n136, Z 
                           => n2458);
   U2101 : MUX2_X1 port map( A => REGISTERS_3_2_port, B => n3119, S => n136, Z 
                           => n2457);
   U2102 : MUX2_X1 port map( A => REGISTERS_3_1_port, B => n3120, S => n136, Z 
                           => n2456);
   U2103 : MUX2_X1 port map( A => REGISTERS_3_0_port, B => n3121, S => n136, Z 
                           => n2455);
   U2104 : OAI21_X1 port map( B1 => n3122, B2 => n3130, A => n3124, ZN => n3129
                           );
   U2105 : MUX2_X1 port map( A => REGISTERS_4_31_port, B => n3089, S => n138, Z
                           => n2454);
   U2106 : MUX2_X1 port map( A => REGISTERS_4_30_port, B => n3091, S => n138, Z
                           => n2453);
   U2107 : MUX2_X1 port map( A => REGISTERS_4_29_port, B => n3092, S => n138, Z
                           => n2452);
   U2108 : MUX2_X1 port map( A => REGISTERS_4_28_port, B => n3093, S => n138, Z
                           => n2451);
   U2109 : MUX2_X1 port map( A => REGISTERS_4_27_port, B => n3094, S => n138, Z
                           => n2450);
   U2110 : MUX2_X1 port map( A => REGISTERS_4_26_port, B => n3095, S => n138, Z
                           => n2449);
   U2111 : MUX2_X1 port map( A => REGISTERS_4_25_port, B => n3096, S => n138, Z
                           => n2448);
   U2112 : MUX2_X1 port map( A => REGISTERS_4_24_port, B => n3097, S => n138, Z
                           => n2447);
   U2113 : MUX2_X1 port map( A => REGISTERS_4_23_port, B => n3098, S => n138, Z
                           => n2446);
   U2114 : MUX2_X1 port map( A => REGISTERS_4_22_port, B => n3099, S => n138, Z
                           => n2445);
   U2115 : MUX2_X1 port map( A => REGISTERS_4_21_port, B => n3100, S => n138, Z
                           => n2444);
   U2116 : MUX2_X1 port map( A => REGISTERS_4_20_port, B => n3101, S => n138, Z
                           => n2443);
   U2117 : MUX2_X1 port map( A => REGISTERS_4_19_port, B => n3102, S => n138, Z
                           => n2442);
   U2118 : MUX2_X1 port map( A => REGISTERS_4_18_port, B => n3103, S => n138, Z
                           => n2441);
   U2119 : MUX2_X1 port map( A => REGISTERS_4_17_port, B => n3104, S => n138, Z
                           => n2440);
   U2120 : MUX2_X1 port map( A => REGISTERS_4_16_port, B => n3105, S => n138, Z
                           => n2439);
   U2121 : MUX2_X1 port map( A => REGISTERS_4_15_port, B => n3106, S => n138, Z
                           => n2438);
   U2122 : MUX2_X1 port map( A => REGISTERS_4_14_port, B => n3107, S => n138, Z
                           => n2437);
   U2123 : MUX2_X1 port map( A => REGISTERS_4_13_port, B => n3108, S => n138, Z
                           => n2436);
   U2124 : MUX2_X1 port map( A => REGISTERS_4_12_port, B => n3109, S => n138, Z
                           => n2435);
   U2125 : MUX2_X1 port map( A => REGISTERS_4_11_port, B => n3110, S => n138, Z
                           => n2434);
   U2126 : MUX2_X1 port map( A => REGISTERS_4_10_port, B => n3111, S => n138, Z
                           => n2433);
   U2127 : MUX2_X1 port map( A => REGISTERS_4_9_port, B => n3112, S => n138, Z 
                           => n2432);
   U2128 : MUX2_X1 port map( A => REGISTERS_4_8_port, B => n3113, S => n138, Z 
                           => n2431);
   U2129 : MUX2_X1 port map( A => REGISTERS_4_7_port, B => n3114, S => n138, Z 
                           => n2430);
   U2130 : MUX2_X1 port map( A => REGISTERS_4_6_port, B => n3115, S => n138, Z 
                           => n2429);
   U2131 : MUX2_X1 port map( A => REGISTERS_4_5_port, B => n3116, S => n138, Z 
                           => n2428);
   U2132 : MUX2_X1 port map( A => REGISTERS_4_4_port, B => n3117, S => n138, Z 
                           => n2427);
   U2133 : MUX2_X1 port map( A => REGISTERS_4_3_port, B => n3118, S => n138, Z 
                           => n2426);
   U2134 : MUX2_X1 port map( A => REGISTERS_4_2_port, B => n3119, S => n138, Z 
                           => n2425);
   U2135 : MUX2_X1 port map( A => REGISTERS_4_1_port, B => n3120, S => n138, Z 
                           => n2424);
   U2136 : MUX2_X1 port map( A => REGISTERS_4_0_port, B => n3121, S => n138, Z 
                           => n2423);
   U2137 : OAI21_X1 port map( B1 => n3122, B2 => n3132, A => n3124, ZN => n3131
                           );
   U2138 : MUX2_X1 port map( A => REGISTERS_5_31_port, B => n3089, S => n132, Z
                           => n2422);
   U2139 : MUX2_X1 port map( A => REGISTERS_5_30_port, B => n3091, S => n132, Z
                           => n2421);
   U2140 : MUX2_X1 port map( A => REGISTERS_5_29_port, B => n3092, S => n132, Z
                           => n2420);
   U2141 : MUX2_X1 port map( A => REGISTERS_5_28_port, B => n3093, S => n132, Z
                           => n2419);
   U2142 : MUX2_X1 port map( A => REGISTERS_5_27_port, B => n3094, S => n132, Z
                           => n2418);
   U2143 : MUX2_X1 port map( A => REGISTERS_5_26_port, B => n3095, S => n132, Z
                           => n2417);
   U2144 : MUX2_X1 port map( A => REGISTERS_5_25_port, B => n3096, S => n132, Z
                           => n2416);
   U2145 : MUX2_X1 port map( A => REGISTERS_5_24_port, B => n3097, S => n132, Z
                           => n2415);
   U2146 : MUX2_X1 port map( A => REGISTERS_5_23_port, B => n3098, S => n132, Z
                           => n2414);
   U2147 : MUX2_X1 port map( A => REGISTERS_5_22_port, B => n3099, S => n132, Z
                           => n2413);
   U2148 : MUX2_X1 port map( A => REGISTERS_5_21_port, B => n3100, S => n132, Z
                           => n2412);
   U2149 : MUX2_X1 port map( A => REGISTERS_5_20_port, B => n3101, S => n132, Z
                           => n2411);
   U2150 : MUX2_X1 port map( A => REGISTERS_5_19_port, B => n3102, S => n132, Z
                           => n2410);
   U2151 : MUX2_X1 port map( A => REGISTERS_5_18_port, B => n3103, S => n132, Z
                           => n2409);
   U2152 : MUX2_X1 port map( A => REGISTERS_5_17_port, B => n3104, S => n132, Z
                           => n2408);
   U2153 : MUX2_X1 port map( A => REGISTERS_5_16_port, B => n3105, S => n132, Z
                           => n2407);
   U2154 : MUX2_X1 port map( A => REGISTERS_5_15_port, B => n3106, S => n132, Z
                           => n2406);
   U2155 : MUX2_X1 port map( A => REGISTERS_5_14_port, B => n3107, S => n132, Z
                           => n2405);
   U2156 : MUX2_X1 port map( A => REGISTERS_5_13_port, B => n3108, S => n132, Z
                           => n2404);
   U2157 : MUX2_X1 port map( A => REGISTERS_5_12_port, B => n3109, S => n132, Z
                           => n2403);
   U2158 : MUX2_X1 port map( A => REGISTERS_5_11_port, B => n3110, S => n132, Z
                           => n2402);
   U2159 : MUX2_X1 port map( A => REGISTERS_5_10_port, B => n3111, S => n132, Z
                           => n2401);
   U2160 : MUX2_X1 port map( A => REGISTERS_5_9_port, B => n3112, S => n132, Z 
                           => n2400);
   U2161 : MUX2_X1 port map( A => REGISTERS_5_8_port, B => n3113, S => n132, Z 
                           => n2399);
   U2162 : MUX2_X1 port map( A => REGISTERS_5_7_port, B => n3114, S => n132, Z 
                           => n2398);
   U2163 : MUX2_X1 port map( A => REGISTERS_5_6_port, B => n3115, S => n132, Z 
                           => n2397);
   U2164 : MUX2_X1 port map( A => REGISTERS_5_5_port, B => n3116, S => n132, Z 
                           => n2396);
   U2165 : MUX2_X1 port map( A => REGISTERS_5_4_port, B => n3117, S => n132, Z 
                           => n2395);
   U2166 : MUX2_X1 port map( A => REGISTERS_5_3_port, B => n3118, S => n132, Z 
                           => n2394);
   U2167 : MUX2_X1 port map( A => REGISTERS_5_2_port, B => n3119, S => n132, Z 
                           => n2393);
   U2168 : MUX2_X1 port map( A => REGISTERS_5_1_port, B => n3120, S => n132, Z 
                           => n2392);
   U2169 : MUX2_X1 port map( A => REGISTERS_5_0_port, B => n3121, S => n132, Z 
                           => n2391);
   U2170 : OAI21_X1 port map( B1 => n3122, B2 => n3134, A => n3124, ZN => n3133
                           );
   U2171 : MUX2_X1 port map( A => REGISTERS_6_31_port, B => n3089, S => n134, Z
                           => n2390);
   U2172 : MUX2_X1 port map( A => REGISTERS_6_30_port, B => n3091, S => n134, Z
                           => n2389);
   U2173 : MUX2_X1 port map( A => REGISTERS_6_29_port, B => n3092, S => n134, Z
                           => n2388);
   U2174 : MUX2_X1 port map( A => REGISTERS_6_28_port, B => n3093, S => n134, Z
                           => n2387);
   U2175 : MUX2_X1 port map( A => REGISTERS_6_27_port, B => n3094, S => n134, Z
                           => n2386);
   U2176 : MUX2_X1 port map( A => REGISTERS_6_26_port, B => n3095, S => n134, Z
                           => n2385);
   U2177 : MUX2_X1 port map( A => REGISTERS_6_25_port, B => n3096, S => n134, Z
                           => n2384);
   U2178 : MUX2_X1 port map( A => REGISTERS_6_24_port, B => n3097, S => n134, Z
                           => n2383);
   U2179 : MUX2_X1 port map( A => REGISTERS_6_23_port, B => n3098, S => n134, Z
                           => n2382);
   U2180 : MUX2_X1 port map( A => REGISTERS_6_22_port, B => n3099, S => n134, Z
                           => n2381);
   U2181 : MUX2_X1 port map( A => REGISTERS_6_21_port, B => n3100, S => n134, Z
                           => n2380);
   U2182 : MUX2_X1 port map( A => REGISTERS_6_20_port, B => n3101, S => n134, Z
                           => n2379);
   U2183 : MUX2_X1 port map( A => REGISTERS_6_19_port, B => n3102, S => n134, Z
                           => n2378);
   U2184 : MUX2_X1 port map( A => REGISTERS_6_18_port, B => n3103, S => n134, Z
                           => n2377);
   U2185 : MUX2_X1 port map( A => REGISTERS_6_17_port, B => n3104, S => n134, Z
                           => n2376);
   U2186 : MUX2_X1 port map( A => REGISTERS_6_16_port, B => n3105, S => n134, Z
                           => n2375);
   U2187 : MUX2_X1 port map( A => REGISTERS_6_15_port, B => n3106, S => n134, Z
                           => n2374);
   U2188 : MUX2_X1 port map( A => REGISTERS_6_14_port, B => n3107, S => n134, Z
                           => n2373);
   U2189 : MUX2_X1 port map( A => REGISTERS_6_13_port, B => n3108, S => n134, Z
                           => n2372);
   U2190 : MUX2_X1 port map( A => REGISTERS_6_12_port, B => n3109, S => n134, Z
                           => n2371);
   U2191 : MUX2_X1 port map( A => REGISTERS_6_11_port, B => n3110, S => n134, Z
                           => n2370);
   U2192 : MUX2_X1 port map( A => REGISTERS_6_10_port, B => n3111, S => n134, Z
                           => n2369);
   U2193 : MUX2_X1 port map( A => REGISTERS_6_9_port, B => n3112, S => n134, Z 
                           => n2368);
   U2194 : MUX2_X1 port map( A => REGISTERS_6_8_port, B => n3113, S => n134, Z 
                           => n2367);
   U2195 : MUX2_X1 port map( A => REGISTERS_6_7_port, B => n3114, S => n134, Z 
                           => n2366);
   U2196 : MUX2_X1 port map( A => REGISTERS_6_6_port, B => n3115, S => n134, Z 
                           => n2365);
   U2197 : MUX2_X1 port map( A => REGISTERS_6_5_port, B => n3116, S => n134, Z 
                           => n2364);
   U2198 : MUX2_X1 port map( A => REGISTERS_6_4_port, B => n3117, S => n134, Z 
                           => n2363);
   U2199 : MUX2_X1 port map( A => REGISTERS_6_3_port, B => n3118, S => n134, Z 
                           => n2362);
   U2200 : MUX2_X1 port map( A => REGISTERS_6_2_port, B => n3119, S => n134, Z 
                           => n2361);
   U2201 : MUX2_X1 port map( A => REGISTERS_6_1_port, B => n3120, S => n134, Z 
                           => n2360);
   U2202 : MUX2_X1 port map( A => REGISTERS_6_0_port, B => n3121, S => n134, Z 
                           => n2359);
   U2203 : OAI21_X1 port map( B1 => n3122, B2 => n3136, A => n3124, ZN => n3135
                           );
   U2204 : MUX2_X1 port map( A => REGISTERS_7_31_port, B => n3089, S => n128, Z
                           => n2358);
   U2205 : MUX2_X1 port map( A => REGISTERS_7_30_port, B => n3091, S => n128, Z
                           => n2357);
   U2206 : MUX2_X1 port map( A => REGISTERS_7_29_port, B => n3092, S => n128, Z
                           => n2356);
   U2207 : MUX2_X1 port map( A => REGISTERS_7_28_port, B => n3093, S => n128, Z
                           => n2355);
   U2208 : MUX2_X1 port map( A => REGISTERS_7_27_port, B => n3094, S => n128, Z
                           => n2354);
   U2209 : MUX2_X1 port map( A => REGISTERS_7_26_port, B => n3095, S => n128, Z
                           => n2353);
   U2210 : MUX2_X1 port map( A => REGISTERS_7_25_port, B => n3096, S => n128, Z
                           => n2352);
   U2211 : MUX2_X1 port map( A => REGISTERS_7_24_port, B => n3097, S => n128, Z
                           => n2351);
   U2212 : MUX2_X1 port map( A => REGISTERS_7_23_port, B => n3098, S => n128, Z
                           => n2350);
   U2213 : MUX2_X1 port map( A => REGISTERS_7_22_port, B => n3099, S => n128, Z
                           => n2349);
   U2214 : MUX2_X1 port map( A => REGISTERS_7_21_port, B => n3100, S => n128, Z
                           => n2348);
   U2215 : MUX2_X1 port map( A => REGISTERS_7_20_port, B => n3101, S => n128, Z
                           => n2347);
   U2216 : MUX2_X1 port map( A => REGISTERS_7_19_port, B => n3102, S => n128, Z
                           => n2346);
   U2217 : MUX2_X1 port map( A => REGISTERS_7_18_port, B => n3103, S => n128, Z
                           => n2345);
   U2218 : MUX2_X1 port map( A => REGISTERS_7_17_port, B => n3104, S => n128, Z
                           => n2344);
   U2219 : MUX2_X1 port map( A => REGISTERS_7_16_port, B => n3105, S => n128, Z
                           => n2343);
   U2220 : MUX2_X1 port map( A => REGISTERS_7_15_port, B => n3106, S => n128, Z
                           => n2342);
   U2221 : MUX2_X1 port map( A => REGISTERS_7_14_port, B => n3107, S => n128, Z
                           => n2341);
   U2222 : MUX2_X1 port map( A => REGISTERS_7_13_port, B => n3108, S => n128, Z
                           => n2340);
   U2223 : MUX2_X1 port map( A => REGISTERS_7_12_port, B => n3109, S => n128, Z
                           => n2339);
   U2224 : MUX2_X1 port map( A => REGISTERS_7_11_port, B => n3110, S => n128, Z
                           => n2338);
   U2225 : MUX2_X1 port map( A => REGISTERS_7_10_port, B => n3111, S => n128, Z
                           => n2337);
   U2226 : MUX2_X1 port map( A => REGISTERS_7_9_port, B => n3112, S => n128, Z 
                           => n2336);
   U2227 : MUX2_X1 port map( A => REGISTERS_7_8_port, B => n3113, S => n128, Z 
                           => n2335);
   U2228 : MUX2_X1 port map( A => REGISTERS_7_7_port, B => n3114, S => n128, Z 
                           => n2334);
   U2229 : MUX2_X1 port map( A => REGISTERS_7_6_port, B => n3115, S => n128, Z 
                           => n2333);
   U2230 : MUX2_X1 port map( A => REGISTERS_7_5_port, B => n3116, S => n128, Z 
                           => n2332);
   U2231 : MUX2_X1 port map( A => REGISTERS_7_4_port, B => n3117, S => n128, Z 
                           => n2331);
   U2232 : MUX2_X1 port map( A => REGISTERS_7_3_port, B => n3118, S => n128, Z 
                           => n2330);
   U2233 : MUX2_X1 port map( A => REGISTERS_7_2_port, B => n3119, S => n128, Z 
                           => n2329);
   U2234 : MUX2_X1 port map( A => REGISTERS_7_1_port, B => n3120, S => n128, Z 
                           => n2328);
   U2235 : MUX2_X1 port map( A => REGISTERS_7_0_port, B => n3121, S => n128, Z 
                           => n2327);
   U2236 : OAI21_X1 port map( B1 => n3122, B2 => n3138, A => n3124, ZN => n3137
                           );
   U2237 : NAND3_X1 port map( A1 => n3139, A2 => n3140, A3 => n3141, ZN => 
                           n3122);
   U2238 : MUX2_X1 port map( A => REGISTERS_8_31_port, B => n3089, S => n130, Z
                           => n2326);
   U2239 : MUX2_X1 port map( A => REGISTERS_8_30_port, B => n3091, S => n130, Z
                           => n2325);
   U2240 : MUX2_X1 port map( A => REGISTERS_8_29_port, B => n3092, S => n130, Z
                           => n2324);
   U2241 : MUX2_X1 port map( A => REGISTERS_8_28_port, B => n3093, S => n130, Z
                           => n2323);
   U2242 : MUX2_X1 port map( A => REGISTERS_8_27_port, B => n3094, S => n130, Z
                           => n2322);
   U2243 : MUX2_X1 port map( A => REGISTERS_8_26_port, B => n3095, S => n130, Z
                           => n2321);
   U2244 : MUX2_X1 port map( A => REGISTERS_8_25_port, B => n3096, S => n130, Z
                           => n2320);
   U2245 : MUX2_X1 port map( A => REGISTERS_8_24_port, B => n3097, S => n130, Z
                           => n2319);
   U2246 : MUX2_X1 port map( A => REGISTERS_8_23_port, B => n3098, S => n130, Z
                           => n2318);
   U2247 : MUX2_X1 port map( A => REGISTERS_8_22_port, B => n3099, S => n130, Z
                           => n2317);
   U2248 : MUX2_X1 port map( A => REGISTERS_8_21_port, B => n3100, S => n130, Z
                           => n2316);
   U2249 : MUX2_X1 port map( A => REGISTERS_8_20_port, B => n3101, S => n130, Z
                           => n2315);
   U2250 : MUX2_X1 port map( A => REGISTERS_8_19_port, B => n3102, S => n130, Z
                           => n2314);
   U2251 : MUX2_X1 port map( A => REGISTERS_8_18_port, B => n3103, S => n130, Z
                           => n2313);
   U2252 : MUX2_X1 port map( A => REGISTERS_8_17_port, B => n3104, S => n130, Z
                           => n2312);
   U2253 : MUX2_X1 port map( A => REGISTERS_8_16_port, B => n3105, S => n130, Z
                           => n2311);
   U2254 : MUX2_X1 port map( A => REGISTERS_8_15_port, B => n3106, S => n130, Z
                           => n2310);
   U2255 : MUX2_X1 port map( A => REGISTERS_8_14_port, B => n3107, S => n130, Z
                           => n2309);
   U2256 : MUX2_X1 port map( A => REGISTERS_8_13_port, B => n3108, S => n130, Z
                           => n2308);
   U2257 : MUX2_X1 port map( A => REGISTERS_8_12_port, B => n3109, S => n130, Z
                           => n2307);
   U2258 : MUX2_X1 port map( A => REGISTERS_8_11_port, B => n3110, S => n130, Z
                           => n2306);
   U2259 : MUX2_X1 port map( A => REGISTERS_8_10_port, B => n3111, S => n130, Z
                           => n2305);
   U2260 : MUX2_X1 port map( A => REGISTERS_8_9_port, B => n3112, S => n130, Z 
                           => n2304);
   U2261 : MUX2_X1 port map( A => REGISTERS_8_8_port, B => n3113, S => n130, Z 
                           => n2303);
   U2262 : MUX2_X1 port map( A => REGISTERS_8_7_port, B => n3114, S => n130, Z 
                           => n2302);
   U2263 : MUX2_X1 port map( A => REGISTERS_8_6_port, B => n3115, S => n130, Z 
                           => n2301);
   U2264 : MUX2_X1 port map( A => REGISTERS_8_5_port, B => n3116, S => n130, Z 
                           => n2300);
   U2265 : MUX2_X1 port map( A => REGISTERS_8_4_port, B => n3117, S => n130, Z 
                           => n2299);
   U2266 : MUX2_X1 port map( A => REGISTERS_8_3_port, B => n3118, S => n130, Z 
                           => n2298);
   U2267 : MUX2_X1 port map( A => REGISTERS_8_2_port, B => n3119, S => n130, Z 
                           => n2297);
   U2268 : MUX2_X1 port map( A => REGISTERS_8_1_port, B => n3120, S => n130, Z 
                           => n2296);
   U2269 : MUX2_X1 port map( A => REGISTERS_8_0_port, B => n3121, S => n130, Z 
                           => n2295);
   U2270 : OAI21_X1 port map( B1 => n3123, B2 => n3143, A => n3124, ZN => n3142
                           );
   U2271 : MUX2_X1 port map( A => REGISTERS_9_31_port, B => n3089, S => n124, Z
                           => n2294);
   U2272 : MUX2_X1 port map( A => REGISTERS_9_30_port, B => n3091, S => n124, Z
                           => n2293);
   U2273 : MUX2_X1 port map( A => REGISTERS_9_29_port, B => n3092, S => n124, Z
                           => n2292);
   U2274 : MUX2_X1 port map( A => REGISTERS_9_28_port, B => n3093, S => n124, Z
                           => n2291);
   U2275 : MUX2_X1 port map( A => REGISTERS_9_27_port, B => n3094, S => n124, Z
                           => n2290);
   U2276 : MUX2_X1 port map( A => REGISTERS_9_26_port, B => n3095, S => n124, Z
                           => n2289);
   U2277 : MUX2_X1 port map( A => REGISTERS_9_25_port, B => n3096, S => n124, Z
                           => n2288);
   U2278 : MUX2_X1 port map( A => REGISTERS_9_24_port, B => n3097, S => n124, Z
                           => n2287);
   U2279 : MUX2_X1 port map( A => REGISTERS_9_23_port, B => n3098, S => n124, Z
                           => n2286);
   U2280 : MUX2_X1 port map( A => REGISTERS_9_22_port, B => n3099, S => n124, Z
                           => n2285);
   U2281 : MUX2_X1 port map( A => REGISTERS_9_21_port, B => n3100, S => n124, Z
                           => n2284);
   U2282 : MUX2_X1 port map( A => REGISTERS_9_20_port, B => n3101, S => n124, Z
                           => n2283);
   U2283 : MUX2_X1 port map( A => REGISTERS_9_19_port, B => n3102, S => n124, Z
                           => n2282);
   U2284 : MUX2_X1 port map( A => REGISTERS_9_18_port, B => n3103, S => n124, Z
                           => n2281);
   U2285 : MUX2_X1 port map( A => REGISTERS_9_17_port, B => n3104, S => n124, Z
                           => n2280);
   U2286 : MUX2_X1 port map( A => REGISTERS_9_16_port, B => n3105, S => n124, Z
                           => n2279);
   U2287 : MUX2_X1 port map( A => REGISTERS_9_15_port, B => n3106, S => n124, Z
                           => n2278);
   U2288 : MUX2_X1 port map( A => REGISTERS_9_14_port, B => n3107, S => n124, Z
                           => n2277);
   U2289 : MUX2_X1 port map( A => REGISTERS_9_13_port, B => n3108, S => n124, Z
                           => n2276);
   U2290 : MUX2_X1 port map( A => REGISTERS_9_12_port, B => n3109, S => n124, Z
                           => n2275);
   U2291 : MUX2_X1 port map( A => REGISTERS_9_11_port, B => n3110, S => n124, Z
                           => n2274);
   U2292 : MUX2_X1 port map( A => REGISTERS_9_10_port, B => n3111, S => n124, Z
                           => n2273);
   U2293 : MUX2_X1 port map( A => REGISTERS_9_9_port, B => n3112, S => n124, Z 
                           => n2272);
   U2294 : MUX2_X1 port map( A => REGISTERS_9_8_port, B => n3113, S => n124, Z 
                           => n2271);
   U2295 : MUX2_X1 port map( A => REGISTERS_9_7_port, B => n3114, S => n124, Z 
                           => n2270);
   U2296 : MUX2_X1 port map( A => REGISTERS_9_6_port, B => n3115, S => n124, Z 
                           => n2269);
   U2297 : MUX2_X1 port map( A => REGISTERS_9_5_port, B => n3116, S => n124, Z 
                           => n2268);
   U2298 : MUX2_X1 port map( A => REGISTERS_9_4_port, B => n3117, S => n124, Z 
                           => n2267);
   U2299 : MUX2_X1 port map( A => REGISTERS_9_3_port, B => n3118, S => n124, Z 
                           => n2266);
   U2300 : MUX2_X1 port map( A => REGISTERS_9_2_port, B => n3119, S => n124, Z 
                           => n2265);
   U2301 : MUX2_X1 port map( A => REGISTERS_9_1_port, B => n3120, S => n124, Z 
                           => n2264);
   U2302 : MUX2_X1 port map( A => REGISTERS_9_0_port, B => n3121, S => n124, Z 
                           => n2263);
   U2303 : OAI21_X1 port map( B1 => n3126, B2 => n3143, A => n3124, ZN => n3144
                           );
   U2304 : MUX2_X1 port map( A => REGISTERS_10_31_port, B => n3089, S => n126, 
                           Z => n2262);
   U2305 : MUX2_X1 port map( A => REGISTERS_10_30_port, B => n3091, S => n126, 
                           Z => n2261);
   U2306 : MUX2_X1 port map( A => REGISTERS_10_29_port, B => n3092, S => n126, 
                           Z => n2260);
   U2307 : MUX2_X1 port map( A => REGISTERS_10_28_port, B => n3093, S => n126, 
                           Z => n2259);
   U2308 : MUX2_X1 port map( A => REGISTERS_10_27_port, B => n3094, S => n126, 
                           Z => n2258);
   U2309 : MUX2_X1 port map( A => REGISTERS_10_26_port, B => n3095, S => n126, 
                           Z => n2257);
   U2310 : MUX2_X1 port map( A => REGISTERS_10_25_port, B => n3096, S => n126, 
                           Z => n2256);
   U2311 : MUX2_X1 port map( A => REGISTERS_10_24_port, B => n3097, S => n126, 
                           Z => n2255);
   U2312 : MUX2_X1 port map( A => REGISTERS_10_23_port, B => n3098, S => n126, 
                           Z => n2254);
   U2313 : MUX2_X1 port map( A => REGISTERS_10_22_port, B => n3099, S => n126, 
                           Z => n2253);
   U2314 : MUX2_X1 port map( A => REGISTERS_10_21_port, B => n3100, S => n126, 
                           Z => n2252);
   U2315 : MUX2_X1 port map( A => REGISTERS_10_20_port, B => n3101, S => n126, 
                           Z => n2251);
   U2316 : MUX2_X1 port map( A => REGISTERS_10_19_port, B => n3102, S => n126, 
                           Z => n2250);
   U2317 : MUX2_X1 port map( A => REGISTERS_10_18_port, B => n3103, S => n126, 
                           Z => n2249);
   U2318 : MUX2_X1 port map( A => REGISTERS_10_17_port, B => n3104, S => n126, 
                           Z => n2248);
   U2319 : MUX2_X1 port map( A => REGISTERS_10_16_port, B => n3105, S => n126, 
                           Z => n2247);
   U2320 : MUX2_X1 port map( A => REGISTERS_10_15_port, B => n3106, S => n126, 
                           Z => n2246);
   U2321 : MUX2_X1 port map( A => REGISTERS_10_14_port, B => n3107, S => n126, 
                           Z => n2245);
   U2322 : MUX2_X1 port map( A => REGISTERS_10_13_port, B => n3108, S => n126, 
                           Z => n2244);
   U2323 : MUX2_X1 port map( A => REGISTERS_10_12_port, B => n3109, S => n126, 
                           Z => n2243);
   U2324 : MUX2_X1 port map( A => REGISTERS_10_11_port, B => n3110, S => n126, 
                           Z => n2242);
   U2325 : MUX2_X1 port map( A => REGISTERS_10_10_port, B => n3111, S => n126, 
                           Z => n2241);
   U2326 : MUX2_X1 port map( A => REGISTERS_10_9_port, B => n3112, S => n126, Z
                           => n2240);
   U2327 : MUX2_X1 port map( A => REGISTERS_10_8_port, B => n3113, S => n126, Z
                           => n2239);
   U2328 : MUX2_X1 port map( A => REGISTERS_10_7_port, B => n3114, S => n126, Z
                           => n2238);
   U2329 : MUX2_X1 port map( A => REGISTERS_10_6_port, B => n3115, S => n126, Z
                           => n2237);
   U2330 : MUX2_X1 port map( A => REGISTERS_10_5_port, B => n3116, S => n126, Z
                           => n2236);
   U2331 : MUX2_X1 port map( A => REGISTERS_10_4_port, B => n3117, S => n126, Z
                           => n2235);
   U2332 : MUX2_X1 port map( A => REGISTERS_10_3_port, B => n3118, S => n126, Z
                           => n2234);
   U2333 : MUX2_X1 port map( A => REGISTERS_10_2_port, B => n3119, S => n126, Z
                           => n2233);
   U2334 : MUX2_X1 port map( A => REGISTERS_10_1_port, B => n3120, S => n126, Z
                           => n2232);
   U2335 : MUX2_X1 port map( A => REGISTERS_10_0_port, B => n3121, S => n126, Z
                           => n2231);
   U2336 : OAI21_X1 port map( B1 => n3128, B2 => n3143, A => n3124, ZN => n3145
                           );
   U2337 : MUX2_X1 port map( A => REGISTERS_11_31_port, B => n3089, S => n120, 
                           Z => n2230);
   U2338 : MUX2_X1 port map( A => REGISTERS_11_30_port, B => n3091, S => n120, 
                           Z => n2229);
   U2339 : MUX2_X1 port map( A => REGISTERS_11_29_port, B => n3092, S => n120, 
                           Z => n2228);
   U2340 : MUX2_X1 port map( A => REGISTERS_11_28_port, B => n3093, S => n120, 
                           Z => n2227);
   U2341 : MUX2_X1 port map( A => REGISTERS_11_27_port, B => n3094, S => n120, 
                           Z => n2226);
   U2342 : MUX2_X1 port map( A => REGISTERS_11_26_port, B => n3095, S => n120, 
                           Z => n2225);
   U2343 : MUX2_X1 port map( A => REGISTERS_11_25_port, B => n3096, S => n120, 
                           Z => n2224);
   U2344 : MUX2_X1 port map( A => REGISTERS_11_24_port, B => n3097, S => n120, 
                           Z => n2223);
   U2345 : MUX2_X1 port map( A => REGISTERS_11_23_port, B => n3098, S => n120, 
                           Z => n2222);
   U2346 : MUX2_X1 port map( A => REGISTERS_11_22_port, B => n3099, S => n120, 
                           Z => n2221);
   U2347 : MUX2_X1 port map( A => REGISTERS_11_21_port, B => n3100, S => n120, 
                           Z => n2220);
   U2348 : MUX2_X1 port map( A => REGISTERS_11_20_port, B => n3101, S => n120, 
                           Z => n2219);
   U2349 : MUX2_X1 port map( A => REGISTERS_11_19_port, B => n3102, S => n120, 
                           Z => n2218);
   U2350 : MUX2_X1 port map( A => REGISTERS_11_18_port, B => n3103, S => n120, 
                           Z => n2217);
   U2351 : MUX2_X1 port map( A => REGISTERS_11_17_port, B => n3104, S => n120, 
                           Z => n2216);
   U2352 : MUX2_X1 port map( A => REGISTERS_11_16_port, B => n3105, S => n120, 
                           Z => n2215);
   U2353 : MUX2_X1 port map( A => REGISTERS_11_15_port, B => n3106, S => n120, 
                           Z => n2214);
   U2354 : MUX2_X1 port map( A => REGISTERS_11_14_port, B => n3107, S => n120, 
                           Z => n2213);
   U2355 : MUX2_X1 port map( A => REGISTERS_11_13_port, B => n3108, S => n120, 
                           Z => n2212);
   U2356 : MUX2_X1 port map( A => REGISTERS_11_12_port, B => n3109, S => n120, 
                           Z => n2211);
   U2357 : MUX2_X1 port map( A => REGISTERS_11_11_port, B => n3110, S => n120, 
                           Z => n2210);
   U2358 : MUX2_X1 port map( A => REGISTERS_11_10_port, B => n3111, S => n120, 
                           Z => n2209);
   U2359 : MUX2_X1 port map( A => REGISTERS_11_9_port, B => n3112, S => n120, Z
                           => n2208);
   U2360 : MUX2_X1 port map( A => REGISTERS_11_8_port, B => n3113, S => n120, Z
                           => n2207);
   U2361 : MUX2_X1 port map( A => REGISTERS_11_7_port, B => n3114, S => n120, Z
                           => n2206);
   U2362 : MUX2_X1 port map( A => REGISTERS_11_6_port, B => n3115, S => n120, Z
                           => n2205);
   U2363 : MUX2_X1 port map( A => REGISTERS_11_5_port, B => n3116, S => n120, Z
                           => n2204);
   U2364 : MUX2_X1 port map( A => REGISTERS_11_4_port, B => n3117, S => n120, Z
                           => n2203);
   U2365 : MUX2_X1 port map( A => REGISTERS_11_3_port, B => n3118, S => n120, Z
                           => n2202);
   U2366 : MUX2_X1 port map( A => REGISTERS_11_2_port, B => n3119, S => n120, Z
                           => n2201);
   U2367 : MUX2_X1 port map( A => REGISTERS_11_1_port, B => n3120, S => n120, Z
                           => n2200);
   U2368 : MUX2_X1 port map( A => REGISTERS_11_0_port, B => n3121, S => n120, Z
                           => n2199);
   U2369 : OAI21_X1 port map( B1 => n3130, B2 => n3143, A => n3124, ZN => n3146
                           );
   U2370 : MUX2_X1 port map( A => REGISTERS_12_31_port, B => n3089, S => n122, 
                           Z => n2198);
   U2371 : MUX2_X1 port map( A => REGISTERS_12_30_port, B => n3091, S => n122, 
                           Z => n2197);
   U2372 : MUX2_X1 port map( A => REGISTERS_12_29_port, B => n3092, S => n122, 
                           Z => n2196);
   U2373 : MUX2_X1 port map( A => REGISTERS_12_28_port, B => n3093, S => n122, 
                           Z => n2195);
   U2374 : MUX2_X1 port map( A => REGISTERS_12_27_port, B => n3094, S => n122, 
                           Z => n2194);
   U2375 : MUX2_X1 port map( A => REGISTERS_12_26_port, B => n3095, S => n122, 
                           Z => n2193);
   U2376 : MUX2_X1 port map( A => REGISTERS_12_25_port, B => n3096, S => n122, 
                           Z => n2192);
   U2377 : MUX2_X1 port map( A => REGISTERS_12_24_port, B => n3097, S => n122, 
                           Z => n2191);
   U2378 : MUX2_X1 port map( A => REGISTERS_12_23_port, B => n3098, S => n122, 
                           Z => n2190);
   U2379 : MUX2_X1 port map( A => REGISTERS_12_22_port, B => n3099, S => n122, 
                           Z => n2189);
   U2380 : MUX2_X1 port map( A => REGISTERS_12_21_port, B => n3100, S => n122, 
                           Z => n2188);
   U2381 : MUX2_X1 port map( A => REGISTERS_12_20_port, B => n3101, S => n122, 
                           Z => n2187);
   U2382 : MUX2_X1 port map( A => REGISTERS_12_19_port, B => n3102, S => n122, 
                           Z => n2186);
   U2383 : MUX2_X1 port map( A => REGISTERS_12_18_port, B => n3103, S => n122, 
                           Z => n2185);
   U2384 : MUX2_X1 port map( A => REGISTERS_12_17_port, B => n3104, S => n122, 
                           Z => n2184);
   U2385 : MUX2_X1 port map( A => REGISTERS_12_16_port, B => n3105, S => n122, 
                           Z => n2183);
   U2386 : MUX2_X1 port map( A => REGISTERS_12_15_port, B => n3106, S => n122, 
                           Z => n2182);
   U2387 : MUX2_X1 port map( A => REGISTERS_12_14_port, B => n3107, S => n122, 
                           Z => n2181);
   U2388 : MUX2_X1 port map( A => REGISTERS_12_13_port, B => n3108, S => n122, 
                           Z => n2180);
   U2389 : MUX2_X1 port map( A => REGISTERS_12_12_port, B => n3109, S => n122, 
                           Z => n2179);
   U2390 : MUX2_X1 port map( A => REGISTERS_12_11_port, B => n3110, S => n122, 
                           Z => n2178);
   U2391 : MUX2_X1 port map( A => REGISTERS_12_10_port, B => n3111, S => n122, 
                           Z => n2177);
   U2392 : MUX2_X1 port map( A => REGISTERS_12_9_port, B => n3112, S => n122, Z
                           => n2176);
   U2393 : MUX2_X1 port map( A => REGISTERS_12_8_port, B => n3113, S => n122, Z
                           => n2175);
   U2394 : MUX2_X1 port map( A => REGISTERS_12_7_port, B => n3114, S => n122, Z
                           => n2174);
   U2395 : MUX2_X1 port map( A => REGISTERS_12_6_port, B => n3115, S => n122, Z
                           => n2173);
   U2396 : MUX2_X1 port map( A => REGISTERS_12_5_port, B => n3116, S => n122, Z
                           => n2172);
   U2397 : MUX2_X1 port map( A => REGISTERS_12_4_port, B => n3117, S => n122, Z
                           => n2171);
   U2398 : MUX2_X1 port map( A => REGISTERS_12_3_port, B => n3118, S => n122, Z
                           => n2170);
   U2399 : MUX2_X1 port map( A => REGISTERS_12_2_port, B => n3119, S => n122, Z
                           => n2169);
   U2400 : MUX2_X1 port map( A => REGISTERS_12_1_port, B => n3120, S => n122, Z
                           => n2168);
   U2401 : MUX2_X1 port map( A => REGISTERS_12_0_port, B => n3121, S => n122, Z
                           => n2167);
   U2402 : OAI21_X1 port map( B1 => n3132, B2 => n3143, A => n3124, ZN => n3147
                           );
   U2403 : MUX2_X1 port map( A => REGISTERS_13_31_port, B => n3089, S => n116, 
                           Z => n2166);
   U2404 : MUX2_X1 port map( A => REGISTERS_13_30_port, B => n3091, S => n116, 
                           Z => n2165);
   U2405 : MUX2_X1 port map( A => REGISTERS_13_29_port, B => n3092, S => n116, 
                           Z => n2164);
   U2406 : MUX2_X1 port map( A => REGISTERS_13_28_port, B => n3093, S => n116, 
                           Z => n2163);
   U2407 : MUX2_X1 port map( A => REGISTERS_13_27_port, B => n3094, S => n116, 
                           Z => n2162);
   U2408 : MUX2_X1 port map( A => REGISTERS_13_26_port, B => n3095, S => n116, 
                           Z => n2161);
   U2409 : MUX2_X1 port map( A => REGISTERS_13_25_port, B => n3096, S => n116, 
                           Z => n2160);
   U2410 : MUX2_X1 port map( A => REGISTERS_13_24_port, B => n3097, S => n116, 
                           Z => n2159);
   U2411 : MUX2_X1 port map( A => REGISTERS_13_23_port, B => n3098, S => n116, 
                           Z => n2158);
   U2412 : MUX2_X1 port map( A => REGISTERS_13_22_port, B => n3099, S => n116, 
                           Z => n2157);
   U2413 : MUX2_X1 port map( A => REGISTERS_13_21_port, B => n3100, S => n116, 
                           Z => n2156);
   U2414 : MUX2_X1 port map( A => REGISTERS_13_20_port, B => n3101, S => n116, 
                           Z => n2155);
   U2415 : MUX2_X1 port map( A => REGISTERS_13_19_port, B => n3102, S => n116, 
                           Z => n2154);
   U2416 : MUX2_X1 port map( A => REGISTERS_13_18_port, B => n3103, S => n116, 
                           Z => n2153);
   U2417 : MUX2_X1 port map( A => REGISTERS_13_17_port, B => n3104, S => n116, 
                           Z => n2152);
   U2418 : MUX2_X1 port map( A => REGISTERS_13_16_port, B => n3105, S => n116, 
                           Z => n2151);
   U2419 : MUX2_X1 port map( A => REGISTERS_13_15_port, B => n3106, S => n116, 
                           Z => n2150);
   U2420 : MUX2_X1 port map( A => REGISTERS_13_14_port, B => n3107, S => n116, 
                           Z => n2149);
   U2421 : MUX2_X1 port map( A => REGISTERS_13_13_port, B => n3108, S => n116, 
                           Z => n2148);
   U2422 : MUX2_X1 port map( A => REGISTERS_13_12_port, B => n3109, S => n116, 
                           Z => n2147);
   U2423 : MUX2_X1 port map( A => REGISTERS_13_11_port, B => n3110, S => n116, 
                           Z => n2146);
   U2424 : MUX2_X1 port map( A => REGISTERS_13_10_port, B => n3111, S => n116, 
                           Z => n2145);
   U2425 : MUX2_X1 port map( A => REGISTERS_13_9_port, B => n3112, S => n116, Z
                           => n2144);
   U2426 : MUX2_X1 port map( A => REGISTERS_13_8_port, B => n3113, S => n116, Z
                           => n2143);
   U2427 : MUX2_X1 port map( A => REGISTERS_13_7_port, B => n3114, S => n116, Z
                           => n2142);
   U2428 : MUX2_X1 port map( A => REGISTERS_13_6_port, B => n3115, S => n116, Z
                           => n2141);
   U2429 : MUX2_X1 port map( A => REGISTERS_13_5_port, B => n3116, S => n116, Z
                           => n2140);
   U2430 : MUX2_X1 port map( A => REGISTERS_13_4_port, B => n3117, S => n116, Z
                           => n2139);
   U2431 : MUX2_X1 port map( A => REGISTERS_13_3_port, B => n3118, S => n116, Z
                           => n2138);
   U2432 : MUX2_X1 port map( A => REGISTERS_13_2_port, B => n3119, S => n116, Z
                           => n2137);
   U2433 : MUX2_X1 port map( A => REGISTERS_13_1_port, B => n3120, S => n116, Z
                           => n2136);
   U2434 : MUX2_X1 port map( A => REGISTERS_13_0_port, B => n3121, S => n116, Z
                           => n2135);
   U2435 : OAI21_X1 port map( B1 => n3134, B2 => n3143, A => n3124, ZN => n3148
                           );
   U2436 : MUX2_X1 port map( A => REGISTERS_14_31_port, B => n3089, S => n118, 
                           Z => n2134);
   U2437 : MUX2_X1 port map( A => REGISTERS_14_30_port, B => n3091, S => n118, 
                           Z => n2133);
   U2438 : MUX2_X1 port map( A => REGISTERS_14_29_port, B => n3092, S => n118, 
                           Z => n2132);
   U2439 : MUX2_X1 port map( A => REGISTERS_14_28_port, B => n3093, S => n118, 
                           Z => n2131);
   U2440 : MUX2_X1 port map( A => REGISTERS_14_27_port, B => n3094, S => n118, 
                           Z => n2130);
   U2441 : MUX2_X1 port map( A => REGISTERS_14_26_port, B => n3095, S => n118, 
                           Z => n2129);
   U2442 : MUX2_X1 port map( A => REGISTERS_14_25_port, B => n3096, S => n118, 
                           Z => n2128);
   U2443 : MUX2_X1 port map( A => REGISTERS_14_24_port, B => n3097, S => n118, 
                           Z => n2127);
   U2444 : MUX2_X1 port map( A => REGISTERS_14_23_port, B => n3098, S => n118, 
                           Z => n2126);
   U2445 : MUX2_X1 port map( A => REGISTERS_14_22_port, B => n3099, S => n118, 
                           Z => n2125);
   U2446 : MUX2_X1 port map( A => REGISTERS_14_21_port, B => n3100, S => n118, 
                           Z => n2124);
   U2447 : MUX2_X1 port map( A => REGISTERS_14_20_port, B => n3101, S => n118, 
                           Z => n2123);
   U2448 : MUX2_X1 port map( A => REGISTERS_14_19_port, B => n3102, S => n118, 
                           Z => n2122);
   U2449 : MUX2_X1 port map( A => REGISTERS_14_18_port, B => n3103, S => n118, 
                           Z => n2121);
   U2450 : MUX2_X1 port map( A => REGISTERS_14_17_port, B => n3104, S => n118, 
                           Z => n2120);
   U2451 : MUX2_X1 port map( A => REGISTERS_14_16_port, B => n3105, S => n118, 
                           Z => n2119);
   U2452 : MUX2_X1 port map( A => REGISTERS_14_15_port, B => n3106, S => n118, 
                           Z => n2118);
   U2453 : MUX2_X1 port map( A => REGISTERS_14_14_port, B => n3107, S => n118, 
                           Z => n2117);
   U2454 : MUX2_X1 port map( A => REGISTERS_14_13_port, B => n3108, S => n118, 
                           Z => n2116);
   U2455 : MUX2_X1 port map( A => REGISTERS_14_12_port, B => n3109, S => n118, 
                           Z => n2115);
   U2456 : MUX2_X1 port map( A => REGISTERS_14_11_port, B => n3110, S => n118, 
                           Z => n2114);
   U2457 : MUX2_X1 port map( A => REGISTERS_14_10_port, B => n3111, S => n118, 
                           Z => n2113);
   U2458 : MUX2_X1 port map( A => REGISTERS_14_9_port, B => n3112, S => n118, Z
                           => n2112);
   U2459 : MUX2_X1 port map( A => REGISTERS_14_8_port, B => n3113, S => n118, Z
                           => n2111);
   U2460 : MUX2_X1 port map( A => REGISTERS_14_7_port, B => n3114, S => n118, Z
                           => n2110);
   U2461 : MUX2_X1 port map( A => REGISTERS_14_6_port, B => n3115, S => n118, Z
                           => n2109);
   U2462 : MUX2_X1 port map( A => REGISTERS_14_5_port, B => n3116, S => n118, Z
                           => n2108);
   U2463 : MUX2_X1 port map( A => REGISTERS_14_4_port, B => n3117, S => n118, Z
                           => n2107);
   U2464 : MUX2_X1 port map( A => REGISTERS_14_3_port, B => n3118, S => n118, Z
                           => n2106);
   U2465 : MUX2_X1 port map( A => REGISTERS_14_2_port, B => n3119, S => n118, Z
                           => n2105);
   U2466 : MUX2_X1 port map( A => REGISTERS_14_1_port, B => n3120, S => n118, Z
                           => n2104);
   U2467 : MUX2_X1 port map( A => REGISTERS_14_0_port, B => n3121, S => n118, Z
                           => n2103);
   U2468 : OAI21_X1 port map( B1 => n3136, B2 => n3143, A => n3124, ZN => n3149
                           );
   U2469 : MUX2_X1 port map( A => REGISTERS_15_31_port, B => n3089, S => n112, 
                           Z => n2102);
   U2470 : MUX2_X1 port map( A => REGISTERS_15_30_port, B => n3091, S => n112, 
                           Z => n2101);
   U2471 : MUX2_X1 port map( A => REGISTERS_15_29_port, B => n3092, S => n112, 
                           Z => n2100);
   U2472 : MUX2_X1 port map( A => REGISTERS_15_28_port, B => n3093, S => n112, 
                           Z => n2099);
   U2473 : MUX2_X1 port map( A => REGISTERS_15_27_port, B => n3094, S => n112, 
                           Z => n2098);
   U2474 : MUX2_X1 port map( A => REGISTERS_15_26_port, B => n3095, S => n112, 
                           Z => n2097);
   U2475 : MUX2_X1 port map( A => REGISTERS_15_25_port, B => n3096, S => n112, 
                           Z => n2096);
   U2476 : MUX2_X1 port map( A => REGISTERS_15_24_port, B => n3097, S => n112, 
                           Z => n2095);
   U2477 : MUX2_X1 port map( A => REGISTERS_15_23_port, B => n3098, S => n112, 
                           Z => n2094);
   U2478 : MUX2_X1 port map( A => REGISTERS_15_22_port, B => n3099, S => n112, 
                           Z => n2093);
   U2479 : MUX2_X1 port map( A => REGISTERS_15_21_port, B => n3100, S => n112, 
                           Z => n2092);
   U2480 : MUX2_X1 port map( A => REGISTERS_15_20_port, B => n3101, S => n112, 
                           Z => n2091);
   U2481 : MUX2_X1 port map( A => REGISTERS_15_19_port, B => n3102, S => n112, 
                           Z => n2090);
   U2482 : MUX2_X1 port map( A => REGISTERS_15_18_port, B => n3103, S => n112, 
                           Z => n2089);
   U2483 : MUX2_X1 port map( A => REGISTERS_15_17_port, B => n3104, S => n112, 
                           Z => n2088);
   U2484 : MUX2_X1 port map( A => REGISTERS_15_16_port, B => n3105, S => n112, 
                           Z => n2087);
   U2485 : MUX2_X1 port map( A => REGISTERS_15_15_port, B => n3106, S => n112, 
                           Z => n2086);
   U2486 : MUX2_X1 port map( A => REGISTERS_15_14_port, B => n3107, S => n112, 
                           Z => n2085);
   U2487 : MUX2_X1 port map( A => REGISTERS_15_13_port, B => n3108, S => n112, 
                           Z => n2084);
   U2488 : MUX2_X1 port map( A => REGISTERS_15_12_port, B => n3109, S => n112, 
                           Z => n2083);
   U2489 : MUX2_X1 port map( A => REGISTERS_15_11_port, B => n3110, S => n112, 
                           Z => n2082);
   U2490 : MUX2_X1 port map( A => REGISTERS_15_10_port, B => n3111, S => n112, 
                           Z => n2081);
   U2491 : MUX2_X1 port map( A => REGISTERS_15_9_port, B => n3112, S => n112, Z
                           => n2080);
   U2492 : MUX2_X1 port map( A => REGISTERS_15_8_port, B => n3113, S => n112, Z
                           => n2079);
   U2493 : MUX2_X1 port map( A => REGISTERS_15_7_port, B => n3114, S => n112, Z
                           => n2078);
   U2494 : MUX2_X1 port map( A => REGISTERS_15_6_port, B => n3115, S => n112, Z
                           => n2077);
   U2495 : MUX2_X1 port map( A => REGISTERS_15_5_port, B => n3116, S => n112, Z
                           => n2076);
   U2496 : MUX2_X1 port map( A => REGISTERS_15_4_port, B => n3117, S => n112, Z
                           => n2075);
   U2497 : MUX2_X1 port map( A => REGISTERS_15_3_port, B => n3118, S => n112, Z
                           => n2074);
   U2498 : MUX2_X1 port map( A => REGISTERS_15_2_port, B => n3119, S => n112, Z
                           => n2073);
   U2499 : MUX2_X1 port map( A => REGISTERS_15_1_port, B => n3120, S => n112, Z
                           => n2072);
   U2500 : MUX2_X1 port map( A => REGISTERS_15_0_port, B => n3121, S => n112, Z
                           => n2071);
   U2501 : OAI21_X1 port map( B1 => n3138, B2 => n3143, A => n3124, ZN => n3150
                           );
   U2502 : NAND3_X1 port map( A1 => n3141, A2 => n3140, A3 => ADD_WR(3), ZN => 
                           n3143);
   U2503 : INV_X1 port map( A => ADD_WR(4), ZN => n3140);
   U2504 : MUX2_X1 port map( A => REGISTERS_16_31_port, B => n3089, S => n114, 
                           Z => n2070);
   U2505 : MUX2_X1 port map( A => REGISTERS_16_30_port, B => n3091, S => n114, 
                           Z => n2069);
   U2506 : MUX2_X1 port map( A => REGISTERS_16_29_port, B => n3092, S => n114, 
                           Z => n2068);
   U2507 : MUX2_X1 port map( A => REGISTERS_16_28_port, B => n3093, S => n114, 
                           Z => n2067);
   U2508 : MUX2_X1 port map( A => REGISTERS_16_27_port, B => n3094, S => n114, 
                           Z => n2066);
   U2509 : MUX2_X1 port map( A => REGISTERS_16_26_port, B => n3095, S => n114, 
                           Z => n2065);
   U2510 : MUX2_X1 port map( A => REGISTERS_16_25_port, B => n3096, S => n114, 
                           Z => n2064);
   U2511 : MUX2_X1 port map( A => REGISTERS_16_24_port, B => n3097, S => n114, 
                           Z => n2063);
   U2512 : MUX2_X1 port map( A => REGISTERS_16_23_port, B => n3098, S => n114, 
                           Z => n2062);
   U2513 : MUX2_X1 port map( A => REGISTERS_16_22_port, B => n3099, S => n114, 
                           Z => n2061);
   U2514 : MUX2_X1 port map( A => REGISTERS_16_21_port, B => n3100, S => n114, 
                           Z => n2060);
   U2515 : MUX2_X1 port map( A => REGISTERS_16_20_port, B => n3101, S => n114, 
                           Z => n2059);
   U2516 : MUX2_X1 port map( A => REGISTERS_16_19_port, B => n3102, S => n114, 
                           Z => n2058);
   U2517 : MUX2_X1 port map( A => REGISTERS_16_18_port, B => n3103, S => n114, 
                           Z => n2057);
   U2518 : MUX2_X1 port map( A => REGISTERS_16_17_port, B => n3104, S => n114, 
                           Z => n2056);
   U2519 : MUX2_X1 port map( A => REGISTERS_16_16_port, B => n3105, S => n114, 
                           Z => n2055);
   U2520 : MUX2_X1 port map( A => REGISTERS_16_15_port, B => n3106, S => n114, 
                           Z => n2054);
   U2521 : MUX2_X1 port map( A => REGISTERS_16_14_port, B => n3107, S => n114, 
                           Z => n2053);
   U2522 : MUX2_X1 port map( A => REGISTERS_16_13_port, B => n3108, S => n114, 
                           Z => n2052);
   U2523 : MUX2_X1 port map( A => REGISTERS_16_12_port, B => n3109, S => n114, 
                           Z => n2051);
   U2524 : MUX2_X1 port map( A => REGISTERS_16_11_port, B => n3110, S => n114, 
                           Z => n2050);
   U2525 : MUX2_X1 port map( A => REGISTERS_16_10_port, B => n3111, S => n114, 
                           Z => n2049);
   U2526 : MUX2_X1 port map( A => REGISTERS_16_9_port, B => n3112, S => n114, Z
                           => n2048);
   U2527 : MUX2_X1 port map( A => REGISTERS_16_8_port, B => n3113, S => n114, Z
                           => n2047);
   U2528 : MUX2_X1 port map( A => REGISTERS_16_7_port, B => n3114, S => n114, Z
                           => n2046);
   U2529 : MUX2_X1 port map( A => REGISTERS_16_6_port, B => n3115, S => n114, Z
                           => n2045);
   U2530 : MUX2_X1 port map( A => REGISTERS_16_5_port, B => n3116, S => n114, Z
                           => n2044);
   U2531 : MUX2_X1 port map( A => REGISTERS_16_4_port, B => n3117, S => n114, Z
                           => n2043);
   U2532 : MUX2_X1 port map( A => REGISTERS_16_3_port, B => n3118, S => n114, Z
                           => n2042);
   U2533 : MUX2_X1 port map( A => REGISTERS_16_2_port, B => n3119, S => n114, Z
                           => n2041);
   U2534 : MUX2_X1 port map( A => REGISTERS_16_1_port, B => n3120, S => n114, Z
                           => n2040);
   U2535 : MUX2_X1 port map( A => REGISTERS_16_0_port, B => n3121, S => n114, Z
                           => n2039);
   U2536 : OAI21_X1 port map( B1 => n3123, B2 => n3152, A => n3124, ZN => n3151
                           );
   U2537 : MUX2_X1 port map( A => REGISTERS_17_31_port, B => n3089, S => n108, 
                           Z => n2038);
   U2538 : MUX2_X1 port map( A => REGISTERS_17_30_port, B => n3091, S => n108, 
                           Z => n2037);
   U2539 : MUX2_X1 port map( A => REGISTERS_17_29_port, B => n3092, S => n108, 
                           Z => n2036);
   U2540 : MUX2_X1 port map( A => REGISTERS_17_28_port, B => n3093, S => n108, 
                           Z => n2035);
   U2541 : MUX2_X1 port map( A => REGISTERS_17_27_port, B => n3094, S => n108, 
                           Z => n2034);
   U2542 : MUX2_X1 port map( A => REGISTERS_17_26_port, B => n3095, S => n108, 
                           Z => n2033);
   U2543 : MUX2_X1 port map( A => REGISTERS_17_25_port, B => n3096, S => n108, 
                           Z => n2032);
   U2544 : MUX2_X1 port map( A => REGISTERS_17_24_port, B => n3097, S => n108, 
                           Z => n2031);
   U2545 : MUX2_X1 port map( A => REGISTERS_17_23_port, B => n3098, S => n108, 
                           Z => n2030);
   U2546 : MUX2_X1 port map( A => REGISTERS_17_22_port, B => n3099, S => n108, 
                           Z => n2029);
   U2547 : MUX2_X1 port map( A => REGISTERS_17_21_port, B => n3100, S => n108, 
                           Z => n2028);
   U2548 : MUX2_X1 port map( A => REGISTERS_17_20_port, B => n3101, S => n108, 
                           Z => n2027);
   U2549 : MUX2_X1 port map( A => REGISTERS_17_19_port, B => n3102, S => n108, 
                           Z => n2026);
   U2550 : MUX2_X1 port map( A => REGISTERS_17_18_port, B => n3103, S => n108, 
                           Z => n2025);
   U2551 : MUX2_X1 port map( A => REGISTERS_17_17_port, B => n3104, S => n108, 
                           Z => n2024);
   U2552 : MUX2_X1 port map( A => REGISTERS_17_16_port, B => n3105, S => n108, 
                           Z => n2023);
   U2553 : MUX2_X1 port map( A => REGISTERS_17_15_port, B => n3106, S => n108, 
                           Z => n2022);
   U2554 : MUX2_X1 port map( A => REGISTERS_17_14_port, B => n3107, S => n108, 
                           Z => n2021);
   U2555 : MUX2_X1 port map( A => REGISTERS_17_13_port, B => n3108, S => n108, 
                           Z => n2020);
   U2556 : MUX2_X1 port map( A => REGISTERS_17_12_port, B => n3109, S => n108, 
                           Z => n2019);
   U2557 : MUX2_X1 port map( A => REGISTERS_17_11_port, B => n3110, S => n108, 
                           Z => n2018);
   U2558 : MUX2_X1 port map( A => REGISTERS_17_10_port, B => n3111, S => n108, 
                           Z => n2017);
   U2559 : MUX2_X1 port map( A => REGISTERS_17_9_port, B => n3112, S => n108, Z
                           => n2016);
   U2560 : MUX2_X1 port map( A => REGISTERS_17_8_port, B => n3113, S => n108, Z
                           => n2015);
   U2561 : MUX2_X1 port map( A => REGISTERS_17_7_port, B => n3114, S => n108, Z
                           => n2014);
   U2562 : MUX2_X1 port map( A => REGISTERS_17_6_port, B => n3115, S => n108, Z
                           => n2013);
   U2563 : MUX2_X1 port map( A => REGISTERS_17_5_port, B => n3116, S => n108, Z
                           => n2012);
   U2564 : MUX2_X1 port map( A => REGISTERS_17_4_port, B => n3117, S => n108, Z
                           => n2011);
   U2565 : MUX2_X1 port map( A => REGISTERS_17_3_port, B => n3118, S => n108, Z
                           => n2010);
   U2566 : MUX2_X1 port map( A => REGISTERS_17_2_port, B => n3119, S => n108, Z
                           => n2009);
   U2567 : MUX2_X1 port map( A => REGISTERS_17_1_port, B => n3120, S => n108, Z
                           => n2008);
   U2568 : MUX2_X1 port map( A => REGISTERS_17_0_port, B => n3121, S => n108, Z
                           => n2007);
   U2569 : OAI21_X1 port map( B1 => n3126, B2 => n3152, A => n3124, ZN => n3153
                           );
   U2570 : MUX2_X1 port map( A => REGISTERS_18_31_port, B => n3089, S => n110, 
                           Z => n2006);
   U2571 : MUX2_X1 port map( A => REGISTERS_18_30_port, B => n3091, S => n110, 
                           Z => n2005);
   U2572 : MUX2_X1 port map( A => REGISTERS_18_29_port, B => n3092, S => n110, 
                           Z => n2004);
   U2573 : MUX2_X1 port map( A => REGISTERS_18_28_port, B => n3093, S => n110, 
                           Z => n2003);
   U2574 : MUX2_X1 port map( A => REGISTERS_18_27_port, B => n3094, S => n110, 
                           Z => n2002);
   U2575 : MUX2_X1 port map( A => REGISTERS_18_26_port, B => n3095, S => n110, 
                           Z => n2001);
   U2576 : MUX2_X1 port map( A => REGISTERS_18_25_port, B => n3096, S => n110, 
                           Z => n2000);
   U2577 : MUX2_X1 port map( A => REGISTERS_18_24_port, B => n3097, S => n110, 
                           Z => n1999);
   U2578 : MUX2_X1 port map( A => REGISTERS_18_23_port, B => n3098, S => n110, 
                           Z => n1998);
   U2579 : MUX2_X1 port map( A => REGISTERS_18_22_port, B => n3099, S => n110, 
                           Z => n1997);
   U2580 : MUX2_X1 port map( A => REGISTERS_18_21_port, B => n3100, S => n110, 
                           Z => n1996);
   U2581 : MUX2_X1 port map( A => REGISTERS_18_20_port, B => n3101, S => n110, 
                           Z => n1995);
   U2582 : MUX2_X1 port map( A => REGISTERS_18_19_port, B => n3102, S => n110, 
                           Z => n1994);
   U2583 : MUX2_X1 port map( A => REGISTERS_18_18_port, B => n3103, S => n110, 
                           Z => n1993);
   U2584 : MUX2_X1 port map( A => REGISTERS_18_17_port, B => n3104, S => n110, 
                           Z => n1992);
   U2585 : MUX2_X1 port map( A => REGISTERS_18_16_port, B => n3105, S => n110, 
                           Z => n1991);
   U2586 : MUX2_X1 port map( A => REGISTERS_18_15_port, B => n3106, S => n110, 
                           Z => n1990);
   U2587 : MUX2_X1 port map( A => REGISTERS_18_14_port, B => n3107, S => n110, 
                           Z => n1989);
   U2588 : MUX2_X1 port map( A => REGISTERS_18_13_port, B => n3108, S => n110, 
                           Z => n1988);
   U2589 : MUX2_X1 port map( A => REGISTERS_18_12_port, B => n3109, S => n110, 
                           Z => n1987);
   U2590 : MUX2_X1 port map( A => REGISTERS_18_11_port, B => n3110, S => n110, 
                           Z => n1986);
   U2591 : MUX2_X1 port map( A => REGISTERS_18_10_port, B => n3111, S => n110, 
                           Z => n1985);
   U2592 : MUX2_X1 port map( A => REGISTERS_18_9_port, B => n3112, S => n110, Z
                           => n1984);
   U2593 : MUX2_X1 port map( A => REGISTERS_18_8_port, B => n3113, S => n110, Z
                           => n1983);
   U2594 : MUX2_X1 port map( A => REGISTERS_18_7_port, B => n3114, S => n110, Z
                           => n1982);
   U2595 : MUX2_X1 port map( A => REGISTERS_18_6_port, B => n3115, S => n110, Z
                           => n1981);
   U2596 : MUX2_X1 port map( A => REGISTERS_18_5_port, B => n3116, S => n110, Z
                           => n1980);
   U2597 : MUX2_X1 port map( A => REGISTERS_18_4_port, B => n3117, S => n110, Z
                           => n1979);
   U2598 : MUX2_X1 port map( A => REGISTERS_18_3_port, B => n3118, S => n110, Z
                           => n1978);
   U2599 : MUX2_X1 port map( A => REGISTERS_18_2_port, B => n3119, S => n110, Z
                           => n1977);
   U2600 : MUX2_X1 port map( A => REGISTERS_18_1_port, B => n3120, S => n110, Z
                           => n1976);
   U2601 : MUX2_X1 port map( A => REGISTERS_18_0_port, B => n3121, S => n110, Z
                           => n1975);
   U2602 : OAI21_X1 port map( B1 => n3128, B2 => n3152, A => n3124, ZN => n3154
                           );
   U2603 : MUX2_X1 port map( A => REGISTERS_19_31_port, B => n3089, S => n104, 
                           Z => n1974);
   U2604 : MUX2_X1 port map( A => REGISTERS_19_30_port, B => n3091, S => n104, 
                           Z => n1973);
   U2605 : MUX2_X1 port map( A => REGISTERS_19_29_port, B => n3092, S => n104, 
                           Z => n1972);
   U2606 : MUX2_X1 port map( A => REGISTERS_19_28_port, B => n3093, S => n104, 
                           Z => n1971);
   U2607 : MUX2_X1 port map( A => REGISTERS_19_27_port, B => n3094, S => n104, 
                           Z => n1970);
   U2608 : MUX2_X1 port map( A => REGISTERS_19_26_port, B => n3095, S => n104, 
                           Z => n1969);
   U2609 : MUX2_X1 port map( A => REGISTERS_19_25_port, B => n3096, S => n104, 
                           Z => n1968);
   U2610 : MUX2_X1 port map( A => REGISTERS_19_24_port, B => n3097, S => n104, 
                           Z => n1967);
   U2611 : MUX2_X1 port map( A => REGISTERS_19_23_port, B => n3098, S => n104, 
                           Z => n1966);
   U2612 : MUX2_X1 port map( A => REGISTERS_19_22_port, B => n3099, S => n104, 
                           Z => n1965);
   U2613 : MUX2_X1 port map( A => REGISTERS_19_21_port, B => n3100, S => n104, 
                           Z => n1964);
   U2614 : MUX2_X1 port map( A => REGISTERS_19_20_port, B => n3101, S => n104, 
                           Z => n1963);
   U2615 : MUX2_X1 port map( A => REGISTERS_19_19_port, B => n3102, S => n104, 
                           Z => n1962);
   U2616 : MUX2_X1 port map( A => REGISTERS_19_18_port, B => n3103, S => n104, 
                           Z => n1961);
   U2617 : MUX2_X1 port map( A => REGISTERS_19_17_port, B => n3104, S => n104, 
                           Z => n1960);
   U2618 : MUX2_X1 port map( A => REGISTERS_19_16_port, B => n3105, S => n104, 
                           Z => n1959);
   U2619 : MUX2_X1 port map( A => REGISTERS_19_15_port, B => n3106, S => n104, 
                           Z => n1958);
   U2620 : MUX2_X1 port map( A => REGISTERS_19_14_port, B => n3107, S => n104, 
                           Z => n1957);
   U2621 : MUX2_X1 port map( A => REGISTERS_19_13_port, B => n3108, S => n104, 
                           Z => n1956);
   U2622 : MUX2_X1 port map( A => REGISTERS_19_12_port, B => n3109, S => n104, 
                           Z => n1955);
   U2623 : MUX2_X1 port map( A => REGISTERS_19_11_port, B => n3110, S => n104, 
                           Z => n1954);
   U2624 : MUX2_X1 port map( A => REGISTERS_19_10_port, B => n3111, S => n104, 
                           Z => n1953);
   U2625 : MUX2_X1 port map( A => REGISTERS_19_9_port, B => n3112, S => n104, Z
                           => n1952);
   U2626 : MUX2_X1 port map( A => REGISTERS_19_8_port, B => n3113, S => n104, Z
                           => n1951);
   U2627 : MUX2_X1 port map( A => REGISTERS_19_7_port, B => n3114, S => n104, Z
                           => n1950);
   U2628 : MUX2_X1 port map( A => REGISTERS_19_6_port, B => n3115, S => n104, Z
                           => n1949);
   U2629 : MUX2_X1 port map( A => REGISTERS_19_5_port, B => n3116, S => n104, Z
                           => n1948);
   U2630 : MUX2_X1 port map( A => REGISTERS_19_4_port, B => n3117, S => n104, Z
                           => n1947);
   U2631 : MUX2_X1 port map( A => REGISTERS_19_3_port, B => n3118, S => n104, Z
                           => n1946);
   U2632 : MUX2_X1 port map( A => REGISTERS_19_2_port, B => n3119, S => n104, Z
                           => n1945);
   U2633 : MUX2_X1 port map( A => REGISTERS_19_1_port, B => n3120, S => n104, Z
                           => n1944);
   U2634 : MUX2_X1 port map( A => REGISTERS_19_0_port, B => n3121, S => n104, Z
                           => n1943);
   U2635 : OAI21_X1 port map( B1 => n3130, B2 => n3152, A => n3124, ZN => n3155
                           );
   U2636 : MUX2_X1 port map( A => REGISTERS_20_31_port, B => n3089, S => n106, 
                           Z => n1942);
   U2637 : MUX2_X1 port map( A => REGISTERS_20_30_port, B => n3091, S => n106, 
                           Z => n1941);
   U2638 : MUX2_X1 port map( A => REGISTERS_20_29_port, B => n3092, S => n106, 
                           Z => n1940);
   U2639 : MUX2_X1 port map( A => REGISTERS_20_28_port, B => n3093, S => n106, 
                           Z => n1939);
   U2640 : MUX2_X1 port map( A => REGISTERS_20_27_port, B => n3094, S => n106, 
                           Z => n1938);
   U2641 : MUX2_X1 port map( A => REGISTERS_20_26_port, B => n3095, S => n106, 
                           Z => n1937);
   U2642 : MUX2_X1 port map( A => REGISTERS_20_25_port, B => n3096, S => n106, 
                           Z => n1936);
   U2643 : MUX2_X1 port map( A => REGISTERS_20_24_port, B => n3097, S => n106, 
                           Z => n1935);
   U2644 : MUX2_X1 port map( A => REGISTERS_20_23_port, B => n3098, S => n106, 
                           Z => n1934);
   U2645 : MUX2_X1 port map( A => REGISTERS_20_22_port, B => n3099, S => n106, 
                           Z => n1933);
   U2646 : MUX2_X1 port map( A => REGISTERS_20_21_port, B => n3100, S => n106, 
                           Z => n1932);
   U2647 : MUX2_X1 port map( A => REGISTERS_20_20_port, B => n3101, S => n106, 
                           Z => n1931);
   U2648 : MUX2_X1 port map( A => REGISTERS_20_19_port, B => n3102, S => n106, 
                           Z => n1930);
   U2649 : MUX2_X1 port map( A => REGISTERS_20_18_port, B => n3103, S => n106, 
                           Z => n1929);
   U2650 : MUX2_X1 port map( A => REGISTERS_20_17_port, B => n3104, S => n106, 
                           Z => n1928);
   U2651 : MUX2_X1 port map( A => REGISTERS_20_16_port, B => n3105, S => n106, 
                           Z => n1927);
   U2652 : MUX2_X1 port map( A => REGISTERS_20_15_port, B => n3106, S => n106, 
                           Z => n1926);
   U2653 : MUX2_X1 port map( A => REGISTERS_20_14_port, B => n3107, S => n106, 
                           Z => n1925);
   U2654 : MUX2_X1 port map( A => REGISTERS_20_13_port, B => n3108, S => n106, 
                           Z => n1924);
   U2655 : MUX2_X1 port map( A => REGISTERS_20_12_port, B => n3109, S => n106, 
                           Z => n1923);
   U2656 : MUX2_X1 port map( A => REGISTERS_20_11_port, B => n3110, S => n106, 
                           Z => n1922);
   U2657 : MUX2_X1 port map( A => REGISTERS_20_10_port, B => n3111, S => n106, 
                           Z => n1921);
   U2658 : MUX2_X1 port map( A => REGISTERS_20_9_port, B => n3112, S => n106, Z
                           => n1920);
   U2659 : MUX2_X1 port map( A => REGISTERS_20_8_port, B => n3113, S => n106, Z
                           => n1919);
   U2660 : MUX2_X1 port map( A => REGISTERS_20_7_port, B => n3114, S => n106, Z
                           => n1918);
   U2661 : MUX2_X1 port map( A => REGISTERS_20_6_port, B => n3115, S => n106, Z
                           => n1917);
   U2662 : MUX2_X1 port map( A => REGISTERS_20_5_port, B => n3116, S => n106, Z
                           => n1916);
   U2663 : MUX2_X1 port map( A => REGISTERS_20_4_port, B => n3117, S => n106, Z
                           => n1915);
   U2664 : MUX2_X1 port map( A => REGISTERS_20_3_port, B => n3118, S => n106, Z
                           => n1914);
   U2665 : MUX2_X1 port map( A => REGISTERS_20_2_port, B => n3119, S => n106, Z
                           => n1913);
   U2666 : MUX2_X1 port map( A => REGISTERS_20_1_port, B => n3120, S => n106, Z
                           => n1912);
   U2667 : MUX2_X1 port map( A => REGISTERS_20_0_port, B => n3121, S => n106, Z
                           => n1911);
   U2668 : OAI21_X1 port map( B1 => n3132, B2 => n3152, A => n3124, ZN => n3156
                           );
   U2669 : MUX2_X1 port map( A => REGISTERS_21_31_port, B => n3089, S => n100, 
                           Z => n1910);
   U2670 : MUX2_X1 port map( A => REGISTERS_21_30_port, B => n3091, S => n100, 
                           Z => n1909);
   U2671 : MUX2_X1 port map( A => REGISTERS_21_29_port, B => n3092, S => n100, 
                           Z => n1908);
   U2672 : MUX2_X1 port map( A => REGISTERS_21_28_port, B => n3093, S => n100, 
                           Z => n1907);
   U2673 : MUX2_X1 port map( A => REGISTERS_21_27_port, B => n3094, S => n100, 
                           Z => n1906);
   U2674 : MUX2_X1 port map( A => REGISTERS_21_26_port, B => n3095, S => n100, 
                           Z => n1905);
   U2675 : MUX2_X1 port map( A => REGISTERS_21_25_port, B => n3096, S => n100, 
                           Z => n1904);
   U2676 : MUX2_X1 port map( A => REGISTERS_21_24_port, B => n3097, S => n100, 
                           Z => n1903);
   U2677 : MUX2_X1 port map( A => REGISTERS_21_23_port, B => n3098, S => n100, 
                           Z => n1902);
   U2678 : MUX2_X1 port map( A => REGISTERS_21_22_port, B => n3099, S => n100, 
                           Z => n1901);
   U2679 : MUX2_X1 port map( A => REGISTERS_21_21_port, B => n3100, S => n100, 
                           Z => n1900);
   U2680 : MUX2_X1 port map( A => REGISTERS_21_20_port, B => n3101, S => n100, 
                           Z => n1899);
   U2681 : MUX2_X1 port map( A => REGISTERS_21_19_port, B => n3102, S => n100, 
                           Z => n1898);
   U2682 : MUX2_X1 port map( A => REGISTERS_21_18_port, B => n3103, S => n100, 
                           Z => n1897);
   U2683 : MUX2_X1 port map( A => REGISTERS_21_17_port, B => n3104, S => n100, 
                           Z => n1896);
   U2684 : MUX2_X1 port map( A => REGISTERS_21_16_port, B => n3105, S => n100, 
                           Z => n1895);
   U2685 : MUX2_X1 port map( A => REGISTERS_21_15_port, B => n3106, S => n100, 
                           Z => n1894);
   U2686 : MUX2_X1 port map( A => REGISTERS_21_14_port, B => n3107, S => n100, 
                           Z => n1893);
   U2687 : MUX2_X1 port map( A => REGISTERS_21_13_port, B => n3108, S => n100, 
                           Z => n1892);
   U2688 : MUX2_X1 port map( A => REGISTERS_21_12_port, B => n3109, S => n100, 
                           Z => n1891);
   U2689 : MUX2_X1 port map( A => REGISTERS_21_11_port, B => n3110, S => n100, 
                           Z => n1890);
   U2690 : MUX2_X1 port map( A => REGISTERS_21_10_port, B => n3111, S => n100, 
                           Z => n1889);
   U2691 : MUX2_X1 port map( A => REGISTERS_21_9_port, B => n3112, S => n100, Z
                           => n1888);
   U2692 : MUX2_X1 port map( A => REGISTERS_21_8_port, B => n3113, S => n100, Z
                           => n1887);
   U2693 : MUX2_X1 port map( A => REGISTERS_21_7_port, B => n3114, S => n100, Z
                           => n1886);
   U2694 : MUX2_X1 port map( A => REGISTERS_21_6_port, B => n3115, S => n100, Z
                           => n1885);
   U2695 : MUX2_X1 port map( A => REGISTERS_21_5_port, B => n3116, S => n100, Z
                           => n1884);
   U2696 : MUX2_X1 port map( A => REGISTERS_21_4_port, B => n3117, S => n100, Z
                           => n1883);
   U2697 : MUX2_X1 port map( A => REGISTERS_21_3_port, B => n3118, S => n100, Z
                           => n1882);
   U2698 : MUX2_X1 port map( A => REGISTERS_21_2_port, B => n3119, S => n100, Z
                           => n1881);
   U2699 : MUX2_X1 port map( A => REGISTERS_21_1_port, B => n3120, S => n100, Z
                           => n1880);
   U2700 : MUX2_X1 port map( A => REGISTERS_21_0_port, B => n3121, S => n100, Z
                           => n1879);
   U2701 : OAI21_X1 port map( B1 => n3134, B2 => n3152, A => n3124, ZN => n3157
                           );
   U2702 : MUX2_X1 port map( A => REGISTERS_22_31_port, B => n3089, S => n102, 
                           Z => n1878);
   U2703 : MUX2_X1 port map( A => REGISTERS_22_30_port, B => n3091, S => n102, 
                           Z => n1877);
   U2704 : MUX2_X1 port map( A => REGISTERS_22_29_port, B => n3092, S => n102, 
                           Z => n1876);
   U2705 : MUX2_X1 port map( A => REGISTERS_22_28_port, B => n3093, S => n102, 
                           Z => n1875);
   U2706 : MUX2_X1 port map( A => REGISTERS_22_27_port, B => n3094, S => n102, 
                           Z => n1874);
   U2707 : MUX2_X1 port map( A => REGISTERS_22_26_port, B => n3095, S => n102, 
                           Z => n1873);
   U2708 : MUX2_X1 port map( A => REGISTERS_22_25_port, B => n3096, S => n102, 
                           Z => n1872);
   U2709 : MUX2_X1 port map( A => REGISTERS_22_24_port, B => n3097, S => n102, 
                           Z => n1871);
   U2710 : MUX2_X1 port map( A => REGISTERS_22_23_port, B => n3098, S => n102, 
                           Z => n1870);
   U2711 : MUX2_X1 port map( A => REGISTERS_22_22_port, B => n3099, S => n102, 
                           Z => n1869);
   U2712 : MUX2_X1 port map( A => REGISTERS_22_21_port, B => n3100, S => n102, 
                           Z => n1868);
   U2713 : MUX2_X1 port map( A => REGISTERS_22_20_port, B => n3101, S => n102, 
                           Z => n1867);
   U2714 : MUX2_X1 port map( A => REGISTERS_22_19_port, B => n3102, S => n102, 
                           Z => n1866);
   U2715 : MUX2_X1 port map( A => REGISTERS_22_18_port, B => n3103, S => n102, 
                           Z => n1865);
   U2716 : MUX2_X1 port map( A => REGISTERS_22_17_port, B => n3104, S => n102, 
                           Z => n1864);
   U2717 : MUX2_X1 port map( A => REGISTERS_22_16_port, B => n3105, S => n102, 
                           Z => n1863);
   U2718 : MUX2_X1 port map( A => REGISTERS_22_15_port, B => n3106, S => n102, 
                           Z => n1862);
   U2719 : MUX2_X1 port map( A => REGISTERS_22_14_port, B => n3107, S => n102, 
                           Z => n1861);
   U2720 : MUX2_X1 port map( A => REGISTERS_22_13_port, B => n3108, S => n102, 
                           Z => n1860);
   U2721 : MUX2_X1 port map( A => REGISTERS_22_12_port, B => n3109, S => n102, 
                           Z => n1859);
   U2722 : MUX2_X1 port map( A => REGISTERS_22_11_port, B => n3110, S => n102, 
                           Z => n1858);
   U2723 : MUX2_X1 port map( A => REGISTERS_22_10_port, B => n3111, S => n102, 
                           Z => n1857);
   U2724 : MUX2_X1 port map( A => REGISTERS_22_9_port, B => n3112, S => n102, Z
                           => n1856);
   U2725 : MUX2_X1 port map( A => REGISTERS_22_8_port, B => n3113, S => n102, Z
                           => n1855);
   U2726 : MUX2_X1 port map( A => REGISTERS_22_7_port, B => n3114, S => n102, Z
                           => n1854);
   U2727 : MUX2_X1 port map( A => REGISTERS_22_6_port, B => n3115, S => n102, Z
                           => n1853);
   U2728 : MUX2_X1 port map( A => REGISTERS_22_5_port, B => n3116, S => n102, Z
                           => n1852);
   U2729 : MUX2_X1 port map( A => REGISTERS_22_4_port, B => n3117, S => n102, Z
                           => n1851);
   U2730 : MUX2_X1 port map( A => REGISTERS_22_3_port, B => n3118, S => n102, Z
                           => n1850);
   U2731 : MUX2_X1 port map( A => REGISTERS_22_2_port, B => n3119, S => n102, Z
                           => n1849);
   U2732 : MUX2_X1 port map( A => REGISTERS_22_1_port, B => n3120, S => n102, Z
                           => n1848);
   U2733 : MUX2_X1 port map( A => REGISTERS_22_0_port, B => n3121, S => n102, Z
                           => n1847);
   U2734 : OAI21_X1 port map( B1 => n3136, B2 => n3152, A => n3124, ZN => n3158
                           );
   U2735 : MUX2_X1 port map( A => REGISTERS_23_31_port, B => n3089, S => n82, Z
                           => n1846);
   U2736 : MUX2_X1 port map( A => REGISTERS_23_30_port, B => n3091, S => n82, Z
                           => n1845);
   U2737 : MUX2_X1 port map( A => REGISTERS_23_29_port, B => n3092, S => n82, Z
                           => n1844);
   U2738 : MUX2_X1 port map( A => REGISTERS_23_28_port, B => n3093, S => n82, Z
                           => n1843);
   U2739 : MUX2_X1 port map( A => REGISTERS_23_27_port, B => n3094, S => n82, Z
                           => n1842);
   U2740 : MUX2_X1 port map( A => REGISTERS_23_26_port, B => n3095, S => n82, Z
                           => n1841);
   U2741 : MUX2_X1 port map( A => REGISTERS_23_25_port, B => n3096, S => n82, Z
                           => n1840);
   U2742 : MUX2_X1 port map( A => REGISTERS_23_24_port, B => n3097, S => n82, Z
                           => n1839);
   U2743 : MUX2_X1 port map( A => REGISTERS_23_23_port, B => n3098, S => n82, Z
                           => n1838);
   U2744 : MUX2_X1 port map( A => REGISTERS_23_22_port, B => n3099, S => n82, Z
                           => n1837);
   U2745 : MUX2_X1 port map( A => REGISTERS_23_21_port, B => n3100, S => n82, Z
                           => n1836);
   U2746 : MUX2_X1 port map( A => REGISTERS_23_20_port, B => n3101, S => n82, Z
                           => n1835);
   U2747 : MUX2_X1 port map( A => REGISTERS_23_19_port, B => n3102, S => n82, Z
                           => n1834);
   U2748 : MUX2_X1 port map( A => REGISTERS_23_18_port, B => n3103, S => n82, Z
                           => n1833);
   U2749 : MUX2_X1 port map( A => REGISTERS_23_17_port, B => n3104, S => n82, Z
                           => n1832);
   U2750 : MUX2_X1 port map( A => REGISTERS_23_16_port, B => n3105, S => n82, Z
                           => n1831);
   U2751 : MUX2_X1 port map( A => REGISTERS_23_15_port, B => n3106, S => n82, Z
                           => n1830);
   U2752 : MUX2_X1 port map( A => REGISTERS_23_14_port, B => n3107, S => n82, Z
                           => n1829);
   U2753 : MUX2_X1 port map( A => REGISTERS_23_13_port, B => n3108, S => n82, Z
                           => n1828);
   U2754 : MUX2_X1 port map( A => REGISTERS_23_12_port, B => n3109, S => n82, Z
                           => n1827);
   U2755 : MUX2_X1 port map( A => REGISTERS_23_11_port, B => n3110, S => n82, Z
                           => n1826);
   U2756 : MUX2_X1 port map( A => REGISTERS_23_10_port, B => n3111, S => n82, Z
                           => n1825);
   U2757 : MUX2_X1 port map( A => REGISTERS_23_9_port, B => n3112, S => n82, Z 
                           => n1824);
   U2758 : MUX2_X1 port map( A => REGISTERS_23_8_port, B => n3113, S => n82, Z 
                           => n1823);
   U2759 : MUX2_X1 port map( A => REGISTERS_23_7_port, B => n3114, S => n82, Z 
                           => n1822);
   U2760 : MUX2_X1 port map( A => REGISTERS_23_6_port, B => n3115, S => n82, Z 
                           => n1821);
   U2761 : MUX2_X1 port map( A => REGISTERS_23_5_port, B => n3116, S => n82, Z 
                           => n1820);
   U2762 : MUX2_X1 port map( A => REGISTERS_23_4_port, B => n3117, S => n82, Z 
                           => n1819);
   U2763 : MUX2_X1 port map( A => REGISTERS_23_3_port, B => n3118, S => n82, Z 
                           => n1818);
   U2764 : MUX2_X1 port map( A => REGISTERS_23_2_port, B => n3119, S => n82, Z 
                           => n1817);
   U2765 : MUX2_X1 port map( A => REGISTERS_23_1_port, B => n3120, S => n82, Z 
                           => n1816);
   U2766 : MUX2_X1 port map( A => REGISTERS_23_0_port, B => n3121, S => n82, Z 
                           => n1815);
   U2767 : OAI21_X1 port map( B1 => n3138, B2 => n3152, A => n3124, ZN => n3159
                           );
   U2768 : NAND3_X1 port map( A1 => n3141, A2 => n3139, A3 => ADD_WR(4), ZN => 
                           n3152);
   U2769 : INV_X1 port map( A => ADD_WR(3), ZN => n3139);
   U2770 : MUX2_X1 port map( A => REGISTERS_24_31_port, B => n3089, S => n84, Z
                           => n1814);
   U2771 : MUX2_X1 port map( A => REGISTERS_24_30_port, B => n3091, S => n84, Z
                           => n1813);
   U2772 : MUX2_X1 port map( A => REGISTERS_24_29_port, B => n3092, S => n84, Z
                           => n1812);
   U2773 : MUX2_X1 port map( A => REGISTERS_24_28_port, B => n3093, S => n84, Z
                           => n1811);
   U2774 : MUX2_X1 port map( A => REGISTERS_24_27_port, B => n3094, S => n84, Z
                           => n1810);
   U2775 : MUX2_X1 port map( A => REGISTERS_24_26_port, B => n3095, S => n84, Z
                           => n1809);
   U2776 : MUX2_X1 port map( A => REGISTERS_24_25_port, B => n3096, S => n84, Z
                           => n1808);
   U2777 : MUX2_X1 port map( A => REGISTERS_24_24_port, B => n3097, S => n84, Z
                           => n1807);
   U2778 : MUX2_X1 port map( A => REGISTERS_24_23_port, B => n3098, S => n84, Z
                           => n1806);
   U2779 : MUX2_X1 port map( A => REGISTERS_24_22_port, B => n3099, S => n84, Z
                           => n1805);
   U2780 : MUX2_X1 port map( A => REGISTERS_24_21_port, B => n3100, S => n84, Z
                           => n1804);
   U2781 : MUX2_X1 port map( A => REGISTERS_24_20_port, B => n3101, S => n84, Z
                           => n1803);
   U2782 : MUX2_X1 port map( A => REGISTERS_24_19_port, B => n3102, S => n84, Z
                           => n1802);
   U2783 : MUX2_X1 port map( A => REGISTERS_24_18_port, B => n3103, S => n84, Z
                           => n1801);
   U2784 : MUX2_X1 port map( A => REGISTERS_24_17_port, B => n3104, S => n84, Z
                           => n1800);
   U2785 : MUX2_X1 port map( A => REGISTERS_24_16_port, B => n3105, S => n84, Z
                           => n1799);
   U2786 : MUX2_X1 port map( A => REGISTERS_24_15_port, B => n3106, S => n84, Z
                           => n1798);
   U2787 : MUX2_X1 port map( A => REGISTERS_24_14_port, B => n3107, S => n84, Z
                           => n1797);
   U2788 : MUX2_X1 port map( A => REGISTERS_24_13_port, B => n3108, S => n84, Z
                           => n1796);
   U2789 : MUX2_X1 port map( A => REGISTERS_24_12_port, B => n3109, S => n84, Z
                           => n1795);
   U2790 : MUX2_X1 port map( A => REGISTERS_24_11_port, B => n3110, S => n84, Z
                           => n1794);
   U2791 : MUX2_X1 port map( A => REGISTERS_24_10_port, B => n3111, S => n84, Z
                           => n1793);
   U2792 : MUX2_X1 port map( A => REGISTERS_24_9_port, B => n3112, S => n84, Z 
                           => n1792);
   U2793 : MUX2_X1 port map( A => REGISTERS_24_8_port, B => n3113, S => n84, Z 
                           => n1791);
   U2794 : MUX2_X1 port map( A => REGISTERS_24_7_port, B => n3114, S => n84, Z 
                           => n1790);
   U2795 : MUX2_X1 port map( A => REGISTERS_24_6_port, B => n3115, S => n84, Z 
                           => n1789);
   U2796 : MUX2_X1 port map( A => REGISTERS_24_5_port, B => n3116, S => n84, Z 
                           => n1788);
   U2797 : MUX2_X1 port map( A => REGISTERS_24_4_port, B => n3117, S => n84, Z 
                           => n1787);
   U2798 : MUX2_X1 port map( A => REGISTERS_24_3_port, B => n3118, S => n84, Z 
                           => n1786);
   U2799 : MUX2_X1 port map( A => REGISTERS_24_2_port, B => n3119, S => n84, Z 
                           => n1785);
   U2800 : MUX2_X1 port map( A => REGISTERS_24_1_port, B => n3120, S => n84, Z 
                           => n1784);
   U2801 : MUX2_X1 port map( A => REGISTERS_24_0_port, B => n3121, S => n84, Z 
                           => n1783);
   U2802 : OAI21_X1 port map( B1 => n3123, B2 => n3161, A => n3124, ZN => n3160
                           );
   U2803 : NAND3_X1 port map( A1 => n3162, A2 => n3163, A3 => n3164, ZN => 
                           n3123);
   U2804 : MUX2_X1 port map( A => REGISTERS_25_31_port, B => n3089, S => n86, Z
                           => n1782);
   U2805 : MUX2_X1 port map( A => REGISTERS_25_30_port, B => n3091, S => n86, Z
                           => n1781);
   U2806 : MUX2_X1 port map( A => REGISTERS_25_29_port, B => n3092, S => n86, Z
                           => n1780);
   U2807 : MUX2_X1 port map( A => REGISTERS_25_28_port, B => n3093, S => n86, Z
                           => n1779);
   U2808 : MUX2_X1 port map( A => REGISTERS_25_27_port, B => n3094, S => n86, Z
                           => n1778);
   U2809 : MUX2_X1 port map( A => REGISTERS_25_26_port, B => n3095, S => n86, Z
                           => n1777);
   U2810 : MUX2_X1 port map( A => REGISTERS_25_25_port, B => n3096, S => n86, Z
                           => n1776);
   U2811 : MUX2_X1 port map( A => REGISTERS_25_24_port, B => n3097, S => n86, Z
                           => n1775);
   U2812 : MUX2_X1 port map( A => REGISTERS_25_23_port, B => n3098, S => n86, Z
                           => n1774);
   U2813 : MUX2_X1 port map( A => REGISTERS_25_22_port, B => n3099, S => n86, Z
                           => n1773);
   U2814 : MUX2_X1 port map( A => REGISTERS_25_21_port, B => n3100, S => n86, Z
                           => n1772);
   U2815 : MUX2_X1 port map( A => REGISTERS_25_20_port, B => n3101, S => n86, Z
                           => n1771);
   U2816 : MUX2_X1 port map( A => REGISTERS_25_19_port, B => n3102, S => n86, Z
                           => n1770);
   U2817 : MUX2_X1 port map( A => REGISTERS_25_18_port, B => n3103, S => n86, Z
                           => n1769);
   U2818 : MUX2_X1 port map( A => REGISTERS_25_17_port, B => n3104, S => n86, Z
                           => n1768);
   U2819 : MUX2_X1 port map( A => REGISTERS_25_16_port, B => n3105, S => n86, Z
                           => n1767);
   U2820 : MUX2_X1 port map( A => REGISTERS_25_15_port, B => n3106, S => n86, Z
                           => n1766);
   U2821 : MUX2_X1 port map( A => REGISTERS_25_14_port, B => n3107, S => n86, Z
                           => n1765);
   U2822 : MUX2_X1 port map( A => REGISTERS_25_13_port, B => n3108, S => n86, Z
                           => n1764);
   U2823 : MUX2_X1 port map( A => REGISTERS_25_12_port, B => n3109, S => n86, Z
                           => n1763);
   U2824 : MUX2_X1 port map( A => REGISTERS_25_11_port, B => n3110, S => n86, Z
                           => n1762);
   U2825 : MUX2_X1 port map( A => REGISTERS_25_10_port, B => n3111, S => n86, Z
                           => n1761);
   U2826 : MUX2_X1 port map( A => REGISTERS_25_9_port, B => n3112, S => n86, Z 
                           => n1760);
   U2827 : MUX2_X1 port map( A => REGISTERS_25_8_port, B => n3113, S => n86, Z 
                           => n1759);
   U2828 : MUX2_X1 port map( A => REGISTERS_25_7_port, B => n3114, S => n86, Z 
                           => n1758);
   U2829 : MUX2_X1 port map( A => REGISTERS_25_6_port, B => n3115, S => n86, Z 
                           => n1757);
   U2830 : MUX2_X1 port map( A => REGISTERS_25_5_port, B => n3116, S => n86, Z 
                           => n1756);
   U2831 : MUX2_X1 port map( A => REGISTERS_25_4_port, B => n3117, S => n86, Z 
                           => n1755);
   U2832 : MUX2_X1 port map( A => REGISTERS_25_3_port, B => n3118, S => n86, Z 
                           => n1754);
   U2833 : MUX2_X1 port map( A => REGISTERS_25_2_port, B => n3119, S => n86, Z 
                           => n1753);
   U2834 : MUX2_X1 port map( A => REGISTERS_25_1_port, B => n3120, S => n86, Z 
                           => n1752);
   U2835 : MUX2_X1 port map( A => REGISTERS_25_0_port, B => n3121, S => n86, Z 
                           => n1751);
   U2836 : OAI21_X1 port map( B1 => n3126, B2 => n3161, A => n3124, ZN => n3165
                           );
   U2837 : NAND3_X1 port map( A1 => n3162, A2 => n3163, A3 => ADD_WR(0), ZN => 
                           n3126);
   U2838 : MUX2_X1 port map( A => REGISTERS_26_31_port, B => n3089, S => n88, Z
                           => n1750);
   U2839 : MUX2_X1 port map( A => REGISTERS_26_30_port, B => n3091, S => n88, Z
                           => n1749);
   U2840 : MUX2_X1 port map( A => REGISTERS_26_29_port, B => n3092, S => n88, Z
                           => n1748);
   U2841 : MUX2_X1 port map( A => REGISTERS_26_28_port, B => n3093, S => n88, Z
                           => n1747);
   U2842 : MUX2_X1 port map( A => REGISTERS_26_27_port, B => n3094, S => n88, Z
                           => n1746);
   U2843 : MUX2_X1 port map( A => REGISTERS_26_26_port, B => n3095, S => n88, Z
                           => n1745);
   U2844 : MUX2_X1 port map( A => REGISTERS_26_25_port, B => n3096, S => n88, Z
                           => n1744);
   U2845 : MUX2_X1 port map( A => REGISTERS_26_24_port, B => n3097, S => n88, Z
                           => n1743);
   U2846 : MUX2_X1 port map( A => REGISTERS_26_23_port, B => n3098, S => n88, Z
                           => n1742);
   U2847 : MUX2_X1 port map( A => REGISTERS_26_22_port, B => n3099, S => n88, Z
                           => n1741);
   U2848 : MUX2_X1 port map( A => REGISTERS_26_21_port, B => n3100, S => n88, Z
                           => n1740);
   U2849 : MUX2_X1 port map( A => REGISTERS_26_20_port, B => n3101, S => n88, Z
                           => n1739);
   U2850 : MUX2_X1 port map( A => REGISTERS_26_19_port, B => n3102, S => n88, Z
                           => n1738);
   U2851 : MUX2_X1 port map( A => REGISTERS_26_18_port, B => n3103, S => n88, Z
                           => n1737);
   U2852 : MUX2_X1 port map( A => REGISTERS_26_17_port, B => n3104, S => n88, Z
                           => n1736);
   U2853 : MUX2_X1 port map( A => REGISTERS_26_16_port, B => n3105, S => n88, Z
                           => n1735);
   U2854 : MUX2_X1 port map( A => REGISTERS_26_15_port, B => n3106, S => n88, Z
                           => n1734);
   U2855 : MUX2_X1 port map( A => REGISTERS_26_14_port, B => n3107, S => n88, Z
                           => n1733);
   U2856 : MUX2_X1 port map( A => REGISTERS_26_13_port, B => n3108, S => n88, Z
                           => n1732);
   U2857 : MUX2_X1 port map( A => REGISTERS_26_12_port, B => n3109, S => n88, Z
                           => n1731);
   U2858 : MUX2_X1 port map( A => REGISTERS_26_11_port, B => n3110, S => n88, Z
                           => n1730);
   U2859 : MUX2_X1 port map( A => REGISTERS_26_10_port, B => n3111, S => n88, Z
                           => n1729);
   U2860 : MUX2_X1 port map( A => REGISTERS_26_9_port, B => n3112, S => n88, Z 
                           => n1728);
   U2861 : MUX2_X1 port map( A => REGISTERS_26_8_port, B => n3113, S => n88, Z 
                           => n1727);
   U2862 : MUX2_X1 port map( A => REGISTERS_26_7_port, B => n3114, S => n88, Z 
                           => n1726);
   U2863 : MUX2_X1 port map( A => REGISTERS_26_6_port, B => n3115, S => n88, Z 
                           => n1725);
   U2864 : MUX2_X1 port map( A => REGISTERS_26_5_port, B => n3116, S => n88, Z 
                           => n1724);
   U2865 : MUX2_X1 port map( A => REGISTERS_26_4_port, B => n3117, S => n88, Z 
                           => n1723);
   U2866 : MUX2_X1 port map( A => REGISTERS_26_3_port, B => n3118, S => n88, Z 
                           => n1722);
   U2867 : MUX2_X1 port map( A => REGISTERS_26_2_port, B => n3119, S => n88, Z 
                           => n1721);
   U2868 : MUX2_X1 port map( A => REGISTERS_26_1_port, B => n3120, S => n88, Z 
                           => n1720);
   U2869 : MUX2_X1 port map( A => REGISTERS_26_0_port, B => n3121, S => n88, Z 
                           => n1719);
   U2870 : OAI21_X1 port map( B1 => n3128, B2 => n3161, A => n3124, ZN => n3166
                           );
   U2871 : NAND3_X1 port map( A1 => n3164, A2 => n3163, A3 => ADD_WR(1), ZN => 
                           n3128);
   U2872 : MUX2_X1 port map( A => REGISTERS_27_31_port, B => n3089, S => n90, Z
                           => n1718);
   U2873 : MUX2_X1 port map( A => REGISTERS_27_30_port, B => n3091, S => n90, Z
                           => n1717);
   U2874 : MUX2_X1 port map( A => REGISTERS_27_29_port, B => n3092, S => n90, Z
                           => n1716);
   U2875 : MUX2_X1 port map( A => REGISTERS_27_28_port, B => n3093, S => n90, Z
                           => n1715);
   U2876 : MUX2_X1 port map( A => REGISTERS_27_27_port, B => n3094, S => n90, Z
                           => n1714);
   U2877 : MUX2_X1 port map( A => REGISTERS_27_26_port, B => n3095, S => n90, Z
                           => n1713);
   U2878 : MUX2_X1 port map( A => REGISTERS_27_25_port, B => n3096, S => n90, Z
                           => n1712);
   U2879 : MUX2_X1 port map( A => REGISTERS_27_24_port, B => n3097, S => n90, Z
                           => n1711);
   U2880 : MUX2_X1 port map( A => REGISTERS_27_23_port, B => n3098, S => n90, Z
                           => n1710);
   U2881 : MUX2_X1 port map( A => REGISTERS_27_22_port, B => n3099, S => n90, Z
                           => n1709);
   U2882 : MUX2_X1 port map( A => REGISTERS_27_21_port, B => n3100, S => n90, Z
                           => n1708);
   U2883 : MUX2_X1 port map( A => REGISTERS_27_20_port, B => n3101, S => n90, Z
                           => n1707);
   U2884 : MUX2_X1 port map( A => REGISTERS_27_19_port, B => n3102, S => n90, Z
                           => n1706);
   U2885 : MUX2_X1 port map( A => REGISTERS_27_18_port, B => n3103, S => n90, Z
                           => n1705);
   U2886 : MUX2_X1 port map( A => REGISTERS_27_17_port, B => n3104, S => n90, Z
                           => n1704);
   U2887 : MUX2_X1 port map( A => REGISTERS_27_16_port, B => n3105, S => n90, Z
                           => n1703);
   U2888 : MUX2_X1 port map( A => REGISTERS_27_15_port, B => n3106, S => n90, Z
                           => n1702);
   U2889 : MUX2_X1 port map( A => REGISTERS_27_14_port, B => n3107, S => n90, Z
                           => n1701);
   U2890 : MUX2_X1 port map( A => REGISTERS_27_13_port, B => n3108, S => n90, Z
                           => n1700);
   U2891 : MUX2_X1 port map( A => REGISTERS_27_12_port, B => n3109, S => n90, Z
                           => n1699);
   U2892 : MUX2_X1 port map( A => REGISTERS_27_11_port, B => n3110, S => n90, Z
                           => n1698);
   U2893 : MUX2_X1 port map( A => REGISTERS_27_10_port, B => n3111, S => n90, Z
                           => n1697);
   U2894 : MUX2_X1 port map( A => REGISTERS_27_9_port, B => n3112, S => n90, Z 
                           => n1696);
   U2895 : MUX2_X1 port map( A => REGISTERS_27_8_port, B => n3113, S => n90, Z 
                           => n1695);
   U2896 : MUX2_X1 port map( A => REGISTERS_27_7_port, B => n3114, S => n90, Z 
                           => n1694);
   U2897 : MUX2_X1 port map( A => REGISTERS_27_6_port, B => n3115, S => n90, Z 
                           => n1693);
   U2898 : MUX2_X1 port map( A => REGISTERS_27_5_port, B => n3116, S => n90, Z 
                           => n1692);
   U2899 : MUX2_X1 port map( A => REGISTERS_27_4_port, B => n3117, S => n90, Z 
                           => n1691);
   U2900 : MUX2_X1 port map( A => REGISTERS_27_3_port, B => n3118, S => n90, Z 
                           => n1690);
   U2901 : MUX2_X1 port map( A => REGISTERS_27_2_port, B => n3119, S => n90, Z 
                           => n1689);
   U2902 : MUX2_X1 port map( A => REGISTERS_27_1_port, B => n3120, S => n90, Z 
                           => n1688);
   U2903 : MUX2_X1 port map( A => REGISTERS_27_0_port, B => n3121, S => n90, Z 
                           => n1687);
   U2904 : OAI21_X1 port map( B1 => n3130, B2 => n3161, A => n3124, ZN => n3167
                           );
   U2905 : NAND3_X1 port map( A1 => ADD_WR(0), A2 => n3163, A3 => ADD_WR(1), ZN
                           => n3130);
   U2906 : INV_X1 port map( A => ADD_WR(2), ZN => n3163);
   U2907 : MUX2_X1 port map( A => REGISTERS_28_31_port, B => n3089, S => n92, Z
                           => n1686);
   U2908 : MUX2_X1 port map( A => REGISTERS_28_30_port, B => n3091, S => n92, Z
                           => n1685);
   U2909 : MUX2_X1 port map( A => REGISTERS_28_29_port, B => n3092, S => n92, Z
                           => n1684);
   U2910 : MUX2_X1 port map( A => REGISTERS_28_28_port, B => n3093, S => n92, Z
                           => n1683);
   U2911 : MUX2_X1 port map( A => REGISTERS_28_27_port, B => n3094, S => n92, Z
                           => n1682);
   U2912 : MUX2_X1 port map( A => REGISTERS_28_26_port, B => n3095, S => n92, Z
                           => n1681);
   U2913 : MUX2_X1 port map( A => REGISTERS_28_25_port, B => n3096, S => n92, Z
                           => n1680);
   U2914 : MUX2_X1 port map( A => REGISTERS_28_24_port, B => n3097, S => n92, Z
                           => n1679);
   U2915 : MUX2_X1 port map( A => REGISTERS_28_23_port, B => n3098, S => n92, Z
                           => n1678);
   U2916 : MUX2_X1 port map( A => REGISTERS_28_22_port, B => n3099, S => n92, Z
                           => n1677);
   U2917 : MUX2_X1 port map( A => REGISTERS_28_21_port, B => n3100, S => n92, Z
                           => n1676);
   U2918 : MUX2_X1 port map( A => REGISTERS_28_20_port, B => n3101, S => n92, Z
                           => n1675);
   U2919 : MUX2_X1 port map( A => REGISTERS_28_19_port, B => n3102, S => n92, Z
                           => n1674);
   U2920 : MUX2_X1 port map( A => REGISTERS_28_18_port, B => n3103, S => n92, Z
                           => n1673);
   U2921 : MUX2_X1 port map( A => REGISTERS_28_17_port, B => n3104, S => n92, Z
                           => n1672);
   U2922 : MUX2_X1 port map( A => REGISTERS_28_16_port, B => n3105, S => n92, Z
                           => n1671);
   U2923 : MUX2_X1 port map( A => REGISTERS_28_15_port, B => n3106, S => n92, Z
                           => n1670);
   U2924 : MUX2_X1 port map( A => REGISTERS_28_14_port, B => n3107, S => n92, Z
                           => n1669);
   U2925 : MUX2_X1 port map( A => REGISTERS_28_13_port, B => n3108, S => n92, Z
                           => n1668);
   U2926 : MUX2_X1 port map( A => REGISTERS_28_12_port, B => n3109, S => n92, Z
                           => n1667);
   U2927 : MUX2_X1 port map( A => REGISTERS_28_11_port, B => n3110, S => n92, Z
                           => n1666);
   U2928 : MUX2_X1 port map( A => REGISTERS_28_10_port, B => n3111, S => n92, Z
                           => n1665);
   U2929 : MUX2_X1 port map( A => REGISTERS_28_9_port, B => n3112, S => n92, Z 
                           => n1664);
   U2930 : MUX2_X1 port map( A => REGISTERS_28_8_port, B => n3113, S => n92, Z 
                           => n1663);
   U2931 : MUX2_X1 port map( A => REGISTERS_28_7_port, B => n3114, S => n92, Z 
                           => n1662);
   U2932 : MUX2_X1 port map( A => REGISTERS_28_6_port, B => n3115, S => n92, Z 
                           => n1661);
   U2933 : MUX2_X1 port map( A => REGISTERS_28_5_port, B => n3116, S => n92, Z 
                           => n1660);
   U2934 : MUX2_X1 port map( A => REGISTERS_28_4_port, B => n3117, S => n92, Z 
                           => n1659);
   U2935 : MUX2_X1 port map( A => REGISTERS_28_3_port, B => n3118, S => n92, Z 
                           => n1658);
   U2936 : MUX2_X1 port map( A => REGISTERS_28_2_port, B => n3119, S => n92, Z 
                           => n1657);
   U2937 : MUX2_X1 port map( A => REGISTERS_28_1_port, B => n3120, S => n92, Z 
                           => n1656);
   U2938 : MUX2_X1 port map( A => REGISTERS_28_0_port, B => n3121, S => n92, Z 
                           => n1655);
   U2939 : OAI21_X1 port map( B1 => n3132, B2 => n3161, A => n3124, ZN => n3168
                           );
   U2940 : NAND3_X1 port map( A1 => n3164, A2 => n3162, A3 => ADD_WR(2), ZN => 
                           n3132);
   U2941 : MUX2_X1 port map( A => REGISTERS_29_31_port, B => n3089, S => n94, Z
                           => n1654);
   U2942 : MUX2_X1 port map( A => REGISTERS_29_30_port, B => n3091, S => n94, Z
                           => n1653);
   U2943 : MUX2_X1 port map( A => REGISTERS_29_29_port, B => n3092, S => n94, Z
                           => n1652);
   U2944 : MUX2_X1 port map( A => REGISTERS_29_28_port, B => n3093, S => n94, Z
                           => n1651);
   U2945 : MUX2_X1 port map( A => REGISTERS_29_27_port, B => n3094, S => n94, Z
                           => n1650);
   U2946 : MUX2_X1 port map( A => REGISTERS_29_26_port, B => n3095, S => n94, Z
                           => n1649);
   U2947 : MUX2_X1 port map( A => REGISTERS_29_25_port, B => n3096, S => n94, Z
                           => n1648);
   U2948 : MUX2_X1 port map( A => REGISTERS_29_24_port, B => n3097, S => n94, Z
                           => n1647);
   U2949 : MUX2_X1 port map( A => REGISTERS_29_23_port, B => n3098, S => n94, Z
                           => n1646);
   U2950 : MUX2_X1 port map( A => REGISTERS_29_22_port, B => n3099, S => n94, Z
                           => n1645);
   U2951 : MUX2_X1 port map( A => REGISTERS_29_21_port, B => n3100, S => n94, Z
                           => n1644);
   U2952 : MUX2_X1 port map( A => REGISTERS_29_20_port, B => n3101, S => n94, Z
                           => n1643);
   U2953 : MUX2_X1 port map( A => REGISTERS_29_19_port, B => n3102, S => n94, Z
                           => n1642);
   U2954 : MUX2_X1 port map( A => REGISTERS_29_18_port, B => n3103, S => n94, Z
                           => n1641);
   U2955 : MUX2_X1 port map( A => REGISTERS_29_17_port, B => n3104, S => n94, Z
                           => n1640);
   U2956 : MUX2_X1 port map( A => REGISTERS_29_16_port, B => n3105, S => n94, Z
                           => n1639);
   U2957 : MUX2_X1 port map( A => REGISTERS_29_15_port, B => n3106, S => n94, Z
                           => n1638);
   U2958 : MUX2_X1 port map( A => REGISTERS_29_14_port, B => n3107, S => n94, Z
                           => n1637);
   U2959 : MUX2_X1 port map( A => REGISTERS_29_13_port, B => n3108, S => n94, Z
                           => n1636);
   U2960 : MUX2_X1 port map( A => REGISTERS_29_12_port, B => n3109, S => n94, Z
                           => n1635);
   U2961 : MUX2_X1 port map( A => REGISTERS_29_11_port, B => n3110, S => n94, Z
                           => n1634);
   U2962 : MUX2_X1 port map( A => REGISTERS_29_10_port, B => n3111, S => n94, Z
                           => n1633);
   U2963 : MUX2_X1 port map( A => REGISTERS_29_9_port, B => n3112, S => n94, Z 
                           => n1632);
   U2964 : MUX2_X1 port map( A => REGISTERS_29_8_port, B => n3113, S => n94, Z 
                           => n1631);
   U2965 : MUX2_X1 port map( A => REGISTERS_29_7_port, B => n3114, S => n94, Z 
                           => n1630);
   U2966 : MUX2_X1 port map( A => REGISTERS_29_6_port, B => n3115, S => n94, Z 
                           => n1629);
   U2967 : MUX2_X1 port map( A => REGISTERS_29_5_port, B => n3116, S => n94, Z 
                           => n1628);
   U2968 : MUX2_X1 port map( A => REGISTERS_29_4_port, B => n3117, S => n94, Z 
                           => n1627);
   U2969 : MUX2_X1 port map( A => REGISTERS_29_3_port, B => n3118, S => n94, Z 
                           => n1626);
   U2970 : MUX2_X1 port map( A => REGISTERS_29_2_port, B => n3119, S => n94, Z 
                           => n1625);
   U2971 : MUX2_X1 port map( A => REGISTERS_29_1_port, B => n3120, S => n94, Z 
                           => n1624);
   U2972 : MUX2_X1 port map( A => REGISTERS_29_0_port, B => n3121, S => n94, Z 
                           => n1623);
   U2973 : OAI21_X1 port map( B1 => n3134, B2 => n3161, A => n3124, ZN => n3169
                           );
   U2974 : NAND3_X1 port map( A1 => ADD_WR(0), A2 => n3162, A3 => ADD_WR(2), ZN
                           => n3134);
   U2975 : INV_X1 port map( A => ADD_WR(1), ZN => n3162);
   U2976 : MUX2_X1 port map( A => REGISTERS_30_31_port, B => n3089, S => n96, Z
                           => n1622);
   U2977 : MUX2_X1 port map( A => REGISTERS_30_30_port, B => n3091, S => n96, Z
                           => n1621);
   U2978 : MUX2_X1 port map( A => REGISTERS_30_29_port, B => n3092, S => n96, Z
                           => n1620);
   U2979 : MUX2_X1 port map( A => REGISTERS_30_28_port, B => n3093, S => n96, Z
                           => n1619);
   U2980 : MUX2_X1 port map( A => REGISTERS_30_27_port, B => n3094, S => n96, Z
                           => n1618);
   U2981 : MUX2_X1 port map( A => REGISTERS_30_26_port, B => n3095, S => n96, Z
                           => n1617);
   U2982 : MUX2_X1 port map( A => REGISTERS_30_25_port, B => n3096, S => n96, Z
                           => n1616);
   U2983 : MUX2_X1 port map( A => REGISTERS_30_24_port, B => n3097, S => n96, Z
                           => n1615);
   U2984 : MUX2_X1 port map( A => REGISTERS_30_23_port, B => n3098, S => n96, Z
                           => n1614);
   U2985 : MUX2_X1 port map( A => REGISTERS_30_22_port, B => n3099, S => n96, Z
                           => n1613);
   U2986 : MUX2_X1 port map( A => REGISTERS_30_21_port, B => n3100, S => n96, Z
                           => n1612);
   U2987 : MUX2_X1 port map( A => REGISTERS_30_20_port, B => n3101, S => n96, Z
                           => n1611);
   U2988 : MUX2_X1 port map( A => REGISTERS_30_19_port, B => n3102, S => n96, Z
                           => n1610);
   U2989 : MUX2_X1 port map( A => REGISTERS_30_18_port, B => n3103, S => n96, Z
                           => n1609);
   U2990 : MUX2_X1 port map( A => REGISTERS_30_17_port, B => n3104, S => n96, Z
                           => n1608);
   U2991 : MUX2_X1 port map( A => REGISTERS_30_16_port, B => n3105, S => n96, Z
                           => n1607);
   U2992 : MUX2_X1 port map( A => REGISTERS_30_15_port, B => n3106, S => n96, Z
                           => n1606);
   U2993 : MUX2_X1 port map( A => REGISTERS_30_14_port, B => n3107, S => n96, Z
                           => n1605);
   U2994 : MUX2_X1 port map( A => REGISTERS_30_13_port, B => n3108, S => n96, Z
                           => n1604);
   U2995 : MUX2_X1 port map( A => REGISTERS_30_12_port, B => n3109, S => n96, Z
                           => n1603);
   U2996 : MUX2_X1 port map( A => REGISTERS_30_11_port, B => n3110, S => n96, Z
                           => n1602);
   U2997 : MUX2_X1 port map( A => REGISTERS_30_10_port, B => n3111, S => n96, Z
                           => n1601);
   U2998 : MUX2_X1 port map( A => REGISTERS_30_9_port, B => n3112, S => n96, Z 
                           => n1600);
   U2999 : MUX2_X1 port map( A => REGISTERS_30_8_port, B => n3113, S => n96, Z 
                           => n1599);
   U3000 : MUX2_X1 port map( A => REGISTERS_30_7_port, B => n3114, S => n96, Z 
                           => n1598);
   U3001 : MUX2_X1 port map( A => REGISTERS_30_6_port, B => n3115, S => n96, Z 
                           => n1597);
   U3002 : MUX2_X1 port map( A => REGISTERS_30_5_port, B => n3116, S => n96, Z 
                           => n1596);
   U3003 : MUX2_X1 port map( A => REGISTERS_30_4_port, B => n3117, S => n96, Z 
                           => n1595);
   U3004 : MUX2_X1 port map( A => REGISTERS_30_3_port, B => n3118, S => n96, Z 
                           => n1594);
   U3005 : MUX2_X1 port map( A => REGISTERS_30_2_port, B => n3119, S => n96, Z 
                           => n1593);
   U3006 : MUX2_X1 port map( A => REGISTERS_30_1_port, B => n3120, S => n96, Z 
                           => n1592);
   U3007 : MUX2_X1 port map( A => REGISTERS_30_0_port, B => n3121, S => n96, Z 
                           => n1591);
   U3008 : OAI21_X1 port map( B1 => n3136, B2 => n3161, A => n3124, ZN => n3170
                           );
   U3009 : NAND3_X1 port map( A1 => ADD_WR(1), A2 => n3164, A3 => ADD_WR(2), ZN
                           => n3136);
   U3010 : INV_X1 port map( A => ADD_WR(0), ZN => n3164);
   U3011 : MUX2_X1 port map( A => REGISTERS_31_31_port, B => n3089, S => n98, Z
                           => n1590);
   U3012 : AND2_X1 port map( A1 => DATAIN(31), A2 => n3124, ZN => n3089);
   U3013 : MUX2_X1 port map( A => REGISTERS_31_30_port, B => n3091, S => n98, Z
                           => n1589);
   U3014 : AND2_X1 port map( A1 => DATAIN(30), A2 => n3124, ZN => n3091);
   U3015 : MUX2_X1 port map( A => REGISTERS_31_29_port, B => n3092, S => n98, Z
                           => n1588);
   U3016 : AND2_X1 port map( A1 => DATAIN(29), A2 => n3124, ZN => n3092);
   U3017 : MUX2_X1 port map( A => REGISTERS_31_28_port, B => n3093, S => n98, Z
                           => n1587);
   U3018 : AND2_X1 port map( A1 => DATAIN(28), A2 => n3124, ZN => n3093);
   U3019 : MUX2_X1 port map( A => REGISTERS_31_27_port, B => n3094, S => n98, Z
                           => n1586);
   U3020 : AND2_X1 port map( A1 => DATAIN(27), A2 => n3124, ZN => n3094);
   U3021 : MUX2_X1 port map( A => REGISTERS_31_26_port, B => n3095, S => n98, Z
                           => n1585);
   U3022 : AND2_X1 port map( A1 => DATAIN(26), A2 => n3124, ZN => n3095);
   U3023 : MUX2_X1 port map( A => REGISTERS_31_25_port, B => n3096, S => n98, Z
                           => n1584);
   U3024 : AND2_X1 port map( A1 => DATAIN(25), A2 => n3124, ZN => n3096);
   U3025 : MUX2_X1 port map( A => REGISTERS_31_24_port, B => n3097, S => n98, Z
                           => n1583);
   U3026 : AND2_X1 port map( A1 => DATAIN(24), A2 => n3124, ZN => n3097);
   U3027 : MUX2_X1 port map( A => REGISTERS_31_23_port, B => n3098, S => n98, Z
                           => n1582);
   U3028 : AND2_X1 port map( A1 => DATAIN(23), A2 => n3124, ZN => n3098);
   U3029 : MUX2_X1 port map( A => REGISTERS_31_22_port, B => n3099, S => n98, Z
                           => n1581);
   U3030 : AND2_X1 port map( A1 => DATAIN(22), A2 => n3124, ZN => n3099);
   U3031 : MUX2_X1 port map( A => REGISTERS_31_21_port, B => n3100, S => n98, Z
                           => n1580);
   U3032 : AND2_X1 port map( A1 => DATAIN(21), A2 => n3124, ZN => n3100);
   U3033 : MUX2_X1 port map( A => REGISTERS_31_20_port, B => n3101, S => n98, Z
                           => n1579);
   U3034 : AND2_X1 port map( A1 => DATAIN(20), A2 => n3124, ZN => n3101);
   U3035 : MUX2_X1 port map( A => REGISTERS_31_19_port, B => n3102, S => n98, Z
                           => n1578);
   U3036 : AND2_X1 port map( A1 => DATAIN(19), A2 => n3124, ZN => n3102);
   U3037 : MUX2_X1 port map( A => REGISTERS_31_18_port, B => n3103, S => n98, Z
                           => n1577);
   U3038 : AND2_X1 port map( A1 => DATAIN(18), A2 => n3124, ZN => n3103);
   U3039 : MUX2_X1 port map( A => REGISTERS_31_17_port, B => n3104, S => n98, Z
                           => n1576);
   U3040 : AND2_X1 port map( A1 => DATAIN(17), A2 => n3124, ZN => n3104);
   U3041 : MUX2_X1 port map( A => REGISTERS_31_16_port, B => n3105, S => n98, Z
                           => n1575);
   U3042 : AND2_X1 port map( A1 => DATAIN(16), A2 => n3124, ZN => n3105);
   U3043 : MUX2_X1 port map( A => REGISTERS_31_15_port, B => n3106, S => n98, Z
                           => n1574);
   U3044 : AND2_X1 port map( A1 => DATAIN(15), A2 => n3124, ZN => n3106);
   U3045 : MUX2_X1 port map( A => REGISTERS_31_14_port, B => n3107, S => n98, Z
                           => n1573);
   U3046 : AND2_X1 port map( A1 => DATAIN(14), A2 => n3124, ZN => n3107);
   U3047 : MUX2_X1 port map( A => REGISTERS_31_13_port, B => n3108, S => n98, Z
                           => n1572);
   U3048 : AND2_X1 port map( A1 => DATAIN(13), A2 => n3124, ZN => n3108);
   U3049 : MUX2_X1 port map( A => REGISTERS_31_12_port, B => n3109, S => n98, Z
                           => n1571);
   U3050 : AND2_X1 port map( A1 => DATAIN(12), A2 => n3124, ZN => n3109);
   U3051 : MUX2_X1 port map( A => REGISTERS_31_11_port, B => n3110, S => n98, Z
                           => n1570);
   U3052 : AND2_X1 port map( A1 => DATAIN(11), A2 => n3124, ZN => n3110);
   U3053 : MUX2_X1 port map( A => REGISTERS_31_10_port, B => n3111, S => n98, Z
                           => n1569);
   U3054 : AND2_X1 port map( A1 => DATAIN(10), A2 => n3124, ZN => n3111);
   U3055 : MUX2_X1 port map( A => REGISTERS_31_9_port, B => n3112, S => n98, Z 
                           => n1568);
   U3056 : AND2_X1 port map( A1 => DATAIN(9), A2 => n3124, ZN => n3112);
   U3057 : MUX2_X1 port map( A => REGISTERS_31_8_port, B => n3113, S => n98, Z 
                           => n1567);
   U3058 : AND2_X1 port map( A1 => DATAIN(8), A2 => n3124, ZN => n3113);
   U3059 : MUX2_X1 port map( A => REGISTERS_31_7_port, B => n3114, S => n98, Z 
                           => n1566);
   U3060 : AND2_X1 port map( A1 => DATAIN(7), A2 => n3124, ZN => n3114);
   U3061 : MUX2_X1 port map( A => REGISTERS_31_6_port, B => n3115, S => n98, Z 
                           => n1565);
   U3062 : AND2_X1 port map( A1 => DATAIN(6), A2 => n3124, ZN => n3115);
   U3063 : MUX2_X1 port map( A => REGISTERS_31_5_port, B => n3116, S => n98, Z 
                           => n1564);
   U3064 : AND2_X1 port map( A1 => DATAIN(5), A2 => n3124, ZN => n3116);
   U3065 : MUX2_X1 port map( A => REGISTERS_31_4_port, B => n3117, S => n98, Z 
                           => n1563);
   U3066 : AND2_X1 port map( A1 => DATAIN(4), A2 => n3124, ZN => n3117);
   U3067 : MUX2_X1 port map( A => REGISTERS_31_3_port, B => n3118, S => n98, Z 
                           => n1562);
   U3068 : AND2_X1 port map( A1 => DATAIN(3), A2 => n3124, ZN => n3118);
   U3069 : MUX2_X1 port map( A => REGISTERS_31_2_port, B => n3119, S => n98, Z 
                           => n1561);
   U3070 : AND2_X1 port map( A1 => DATAIN(2), A2 => n3124, ZN => n3119);
   U3071 : MUX2_X1 port map( A => REGISTERS_31_1_port, B => n3120, S => n98, Z 
                           => n1560);
   U3072 : AND2_X1 port map( A1 => DATAIN(1), A2 => n3124, ZN => n3120);
   U3073 : MUX2_X1 port map( A => REGISTERS_31_0_port, B => n3121, S => n98, Z 
                           => n1559);
   U3074 : OAI21_X1 port map( B1 => n3138, B2 => n3161, A => n3124, ZN => n3171
                           );
   U3075 : NAND3_X1 port map( A1 => ADD_WR(3), A2 => n3141, A3 => ADD_WR(4), ZN
                           => n3161);
   U3076 : AND2_X1 port map( A1 => WR, A2 => ENABLE, ZN => n3141);
   U3077 : NAND3_X1 port map( A1 => ADD_WR(1), A2 => ADD_WR(0), A3 => ADD_WR(2)
                           , ZN => n3138);
   U3078 : AND2_X1 port map( A1 => DATAIN(0), A2 => n3124, ZN => n3121);
   U3079 : OAI21_X1 port map( B1 => n3086, B2 => n49, A => n3172, ZN => n1558);
   U3080 : OAI21_X1 port map( B1 => n3086, B2 => n50, A => n3172, ZN => n1557);
   U3081 : OAI21_X1 port map( B1 => n3086, B2 => n51, A => n3172, ZN => n1556);
   U3082 : OAI21_X1 port map( B1 => n3086, B2 => n52, A => n3172, ZN => n1555);
   U3083 : OAI21_X1 port map( B1 => n3086, B2 => n53, A => n3172, ZN => n1554);
   U3084 : OAI21_X1 port map( B1 => n3086, B2 => n54, A => n3172, ZN => n1553);
   U3085 : OAI21_X1 port map( B1 => n3086, B2 => n55, A => n3172, ZN => n1552);
   U3086 : OAI21_X1 port map( B1 => n3086, B2 => n56, A => n3172, ZN => n1551);
   U3087 : OAI21_X1 port map( B1 => n3086, B2 => n57, A => n3172, ZN => n1550);
   U3088 : OAI21_X1 port map( B1 => n3086, B2 => n58, A => n3172, ZN => n1549);
   U3089 : OAI21_X1 port map( B1 => n3086, B2 => n59, A => n3172, ZN => n1548);
   U3090 : OAI21_X1 port map( B1 => n3086, B2 => n60, A => n3172, ZN => n1547);
   U3091 : OAI21_X1 port map( B1 => n3086, B2 => n61, A => n3172, ZN => n1546);
   U3092 : OAI21_X1 port map( B1 => n3086, B2 => n62, A => n3172, ZN => n1545);
   U3093 : OAI21_X1 port map( B1 => n3086, B2 => n63, A => n3172, ZN => n1544);
   U3094 : OAI21_X1 port map( B1 => n3086, B2 => n64, A => n3172, ZN => n1543);
   U3095 : OAI21_X1 port map( B1 => n3086, B2 => n65, A => n3172, ZN => n1542);
   U3096 : OAI21_X1 port map( B1 => n3086, B2 => n66, A => n3172, ZN => n1541);
   U3097 : OAI21_X1 port map( B1 => n3086, B2 => n67, A => n3172, ZN => n1540);
   U3098 : OAI21_X1 port map( B1 => n3086, B2 => n68, A => n3172, ZN => n1539);
   U3099 : OAI21_X1 port map( B1 => n3086, B2 => n69, A => n3172, ZN => n1538);
   U3100 : OAI21_X1 port map( B1 => n3086, B2 => n70, A => n3172, ZN => n1537);
   U3101 : OAI21_X1 port map( B1 => n3086, B2 => n71, A => n3172, ZN => n1536);
   U3102 : OAI21_X1 port map( B1 => n3086, B2 => n72, A => n3172, ZN => n1535);
   U3103 : OAI21_X1 port map( B1 => n3086, B2 => n73, A => n3172, ZN => n1534);
   U3104 : OAI21_X1 port map( B1 => n3086, B2 => n74, A => n3172, ZN => n1533);
   U3105 : OAI21_X1 port map( B1 => n3086, B2 => n75, A => n3172, ZN => n1532);
   U3106 : OAI21_X1 port map( B1 => n3086, B2 => n76, A => n3172, ZN => n1531);
   U3107 : OAI21_X1 port map( B1 => n3086, B2 => n77, A => n3172, ZN => n1530);
   U3108 : OAI21_X1 port map( B1 => n3086, B2 => n78, A => n3172, ZN => n1529);
   U3109 : OAI21_X1 port map( B1 => n3086, B2 => n79, A => n3172, ZN => n1528);
   U3110 : OAI21_X1 port map( B1 => n3086, B2 => n80, A => n3172, ZN => n1527);
   U3111 : MUX2_X1 port map( A => N220, B => n3299, S => n3088, Z => n1494);
   U3112 : MUX2_X1 port map( A => N219, B => n3297, S => n3088, Z => n1493);
   U3113 : MUX2_X1 port map( A => N218, B => n3295, S => n3088, Z => n1492);
   U3114 : MUX2_X1 port map( A => N217, B => n3293, S => n3088, Z => n1491);
   U3115 : MUX2_X1 port map( A => N216, B => n3291, S => n3088, Z => n1490);
   U3116 : MUX2_X1 port map( A => N215, B => n3289, S => n3088, Z => n1489);
   U3117 : MUX2_X1 port map( A => N214, B => n3287, S => n3088, Z => n1488);
   U3118 : MUX2_X1 port map( A => N213, B => n3285, S => n3088, Z => n1487);
   U3119 : MUX2_X1 port map( A => N212, B => n3283, S => n3088, Z => n1486);
   U3120 : MUX2_X1 port map( A => N211, B => n3281, S => n3088, Z => n1485);
   U3121 : MUX2_X1 port map( A => N210, B => n3279, S => n3088, Z => n1484);
   U3122 : MUX2_X1 port map( A => N209, B => n3277, S => n3088, Z => n1483);
   U3123 : MUX2_X1 port map( A => N208, B => n3275, S => n3088, Z => n1482);
   U3124 : MUX2_X1 port map( A => N207, B => n3273, S => n3088, Z => n1481);
   U3125 : MUX2_X1 port map( A => N206, B => n3271, S => n3088, Z => n1480);
   U3126 : MUX2_X1 port map( A => N205, B => n3269, S => n3088, Z => n1479);
   U3127 : MUX2_X1 port map( A => N204, B => n3267, S => n3088, Z => n1478);
   U3128 : MUX2_X1 port map( A => N203, B => n3265, S => n3088, Z => n1477);
   U3129 : MUX2_X1 port map( A => N202, B => n3263, S => n3088, Z => n1476);
   U3130 : MUX2_X1 port map( A => N201, B => n3261, S => n3088, Z => n1475);
   U3131 : MUX2_X1 port map( A => N200, B => n3259, S => n3088, Z => n1474);
   U3132 : MUX2_X1 port map( A => N199, B => n3257, S => n3088, Z => n1473);
   U3133 : MUX2_X1 port map( A => N198, B => n3255, S => n3088, Z => n1472);
   U3134 : MUX2_X1 port map( A => N197, B => n3253, S => n3088, Z => n1471);
   U3135 : MUX2_X1 port map( A => N196, B => n3251, S => n3088, Z => n1470);
   U3136 : MUX2_X1 port map( A => N195, B => n3249, S => n3088, Z => n1469);
   U3137 : MUX2_X1 port map( A => N194, B => n3247, S => n3088, Z => n1468);
   U3138 : MUX2_X1 port map( A => N193, B => n3245, S => n3088, Z => n1467);
   U3139 : MUX2_X1 port map( A => N192, B => n3243, S => n3088, Z => n1466);
   U3140 : MUX2_X1 port map( A => N191, B => n3241, S => n3088, Z => n1465);
   U3141 : MUX2_X1 port map( A => N190, B => n3239, S => n3088, Z => n1464);
   U3142 : MUX2_X1 port map( A => N189, B => n3237, S => n3088, Z => n1463);
   U3143 : MUX2_X1 port map( A => N187, B => n3235, S => n3088, Z => n1461);
   U3144 : MUX2_X1 port map( A => N186, B => n3233, S => n3088, Z => n1459);
   U3145 : MUX2_X1 port map( A => N185, B => n3231, S => n3088, Z => n1457);
   U3146 : MUX2_X1 port map( A => N184, B => n3229, S => n3088, Z => n1455);
   U3147 : MUX2_X1 port map( A => N183, B => n3227, S => n3088, Z => n1453);
   U3148 : MUX2_X1 port map( A => N182, B => n3225, S => n3088, Z => n1451);
   U3149 : MUX2_X1 port map( A => N181, B => n3223, S => n3088, Z => n1449);
   U3150 : MUX2_X1 port map( A => N180, B => n3221, S => n3088, Z => n1447);
   U3151 : MUX2_X1 port map( A => N179, B => n3219, S => n3088, Z => n1445);
   U3152 : MUX2_X1 port map( A => N178, B => n3217, S => n3088, Z => n1443);
   U3153 : MUX2_X1 port map( A => N177, B => n3215, S => n3088, Z => n1441);
   U3154 : MUX2_X1 port map( A => N176, B => n3213, S => n3088, Z => n1439);
   U3155 : MUX2_X1 port map( A => N175, B => n3211, S => n3088, Z => n1437);
   U3156 : MUX2_X1 port map( A => N174, B => n3209, S => n3088, Z => n1435);
   U3157 : MUX2_X1 port map( A => N173, B => n3207, S => n3088, Z => n1433);
   U3158 : MUX2_X1 port map( A => N172, B => n3205, S => n3088, Z => n1431);
   U3159 : MUX2_X1 port map( A => N171, B => n3203, S => n3088, Z => n1429);
   U3160 : MUX2_X1 port map( A => N170, B => n3201, S => n3088, Z => n1427);
   U3161 : MUX2_X1 port map( A => N169, B => n3199, S => n3088, Z => n1425);
   U3162 : MUX2_X1 port map( A => N168, B => n3197, S => n3088, Z => n1423);
   U3163 : MUX2_X1 port map( A => N167, B => n3195, S => n3088, Z => n1421);
   U3164 : MUX2_X1 port map( A => N166, B => n3193, S => n3088, Z => n1419);
   U3165 : MUX2_X1 port map( A => N165, B => n3191, S => n3088, Z => n1417);
   U3166 : MUX2_X1 port map( A => N164, B => n3189, S => n3088, Z => n1415);
   U3167 : MUX2_X1 port map( A => N163, B => n3187, S => n3088, Z => n1413);
   U3168 : MUX2_X1 port map( A => N162, B => n3185, S => n3088, Z => n1411);
   U3169 : MUX2_X1 port map( A => N161, B => n3183, S => n3088, Z => n1409);
   U3170 : MUX2_X1 port map( A => N160, B => n3181, S => n3088, Z => n1407);
   U3171 : MUX2_X1 port map( A => N159, B => n3179, S => n3088, Z => n1405);
   U3172 : MUX2_X1 port map( A => N158, B => n3177, S => n3088, Z => n1403);
   U3173 : MUX2_X1 port map( A => N157, B => n3175, S => n3088, Z => n1401);
   U3174 : MUX2_X1 port map( A => N156, B => n3173, S => n3088, Z => n1399);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_entity.all;

entity Addr_Transformer_Addr_bits5_M4_in_loc_out12 is

   port( ENABLE, RD1, RD2, WR : in std_logic;  ADDR_WR_IN, ADDR_RD1_IN, 
         ADDR_RD2_IN : in std_logic_vector (3 downto 0);  CWP : in 
         std_logic_vector (4 downto 0);  ADDR_WR_OUT, ADDR_RD1_OUT, 
         ADDR_RD2_OUT : out std_logic_vector (4 downto 0));

end Addr_Transformer_Addr_bits5_M4_in_loc_out12;

architecture SYN_Behavioral of Addr_Transformer_Addr_bits5_M4_in_loc_out12 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N29, N52, N75, N76, N77, N78, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10
      , n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, 
      n25, n26, n27, n28, n29_port, n30, n31, n32, n33, n34, n35, n36, n37, n38
      , n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, 
      n52_port, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65
      , n66, n67, n68, n69, n70, n71, n72, n73, n74, n75_port, n76_port, 
      n77_port, n78_port, n79, n80, n81, n82, n83 : std_logic;

begin
   
   ADDR_WR_OUT_reg_4_inst : DLH_X1 port map( G => N78, D => N75, Q => 
                           ADDR_WR_OUT(4));
   ADDR_WR_OUT_reg_3_inst : DLH_X1 port map( G => N78, D => n80, Q => 
                           ADDR_WR_OUT(3));
   ADDR_WR_OUT_reg_2_inst : DLH_X1 port map( G => N78, D => n81, Q => 
                           ADDR_WR_OUT(2));
   ADDR_WR_OUT_reg_1_inst : DLH_X1 port map( G => N78, D => n82, Q => 
                           ADDR_WR_OUT(1));
   ADDR_WR_OUT_reg_0_inst : DLH_X1 port map( G => N78, D => n83, Q => 
                           ADDR_WR_OUT(0));
   ADDR_RD1_OUT_reg_4_inst : DLH_X1 port map( G => N76, D => N29, Q => 
                           ADDR_RD1_OUT(4));
   ADDR_RD1_OUT_reg_3_inst : DLH_X1 port map( G => N76, D => n72, Q => 
                           ADDR_RD1_OUT(3));
   ADDR_RD1_OUT_reg_2_inst : DLH_X1 port map( G => N76, D => n73, Q => 
                           ADDR_RD1_OUT(2));
   ADDR_RD1_OUT_reg_1_inst : DLH_X1 port map( G => N76, D => n74, Q => 
                           ADDR_RD1_OUT(1));
   ADDR_RD1_OUT_reg_0_inst : DLH_X1 port map( G => N76, D => n75_port, Q => 
                           ADDR_RD1_OUT(0));
   ADDR_RD2_OUT_reg_4_inst : DLH_X1 port map( G => N77, D => N52, Q => 
                           ADDR_RD2_OUT(4));
   ADDR_RD2_OUT_reg_3_inst : DLH_X1 port map( G => N77, D => n76_port, Q => 
                           ADDR_RD2_OUT(3));
   ADDR_RD2_OUT_reg_2_inst : DLH_X1 port map( G => N77, D => n77_port, Q => 
                           ADDR_RD2_OUT(2));
   ADDR_RD2_OUT_reg_1_inst : DLH_X1 port map( G => N77, D => n78_port, Q => 
                           ADDR_RD2_OUT(1));
   ADDR_RD2_OUT_reg_0_inst : DLH_X1 port map( G => N77, D => n79, Q => 
                           ADDR_RD2_OUT(0));
   U3 : XOR2_X1 port map( A => ADDR_RD1_IN(3), B => n1, Z => n72);
   U4 : NOR2_X1 port map( A1 => n2, A2 => n3, ZN => n1);
   U5 : XOR2_X1 port map( A => CWP(3), B => n4, Z => n3);
   U6 : XOR2_X1 port map( A => n5, B => n6, Z => n73);
   U7 : NAND2_X1 port map( A1 => n7, A2 => n8, ZN => n6);
   U8 : XOR2_X1 port map( A => n9, B => n10, Z => n7);
   U9 : XNOR2_X1 port map( A => ADDR_RD1_IN(1), B => n11, ZN => n74);
   U10 : NAND2_X1 port map( A1 => n12, A2 => n8, ZN => n11);
   U11 : XOR2_X1 port map( A => n13, B => n14, Z => n12);
   U12 : XOR2_X1 port map( A => ADDR_RD1_IN(0), B => n15, Z => n75_port);
   U13 : NOR2_X1 port map( A1 => n2, A2 => n16, ZN => n15);
   U14 : XOR2_X1 port map( A => ADDR_RD2_IN(3), B => n17, Z => n76_port);
   U15 : NOR2_X1 port map( A1 => n18, A2 => n19, ZN => n17);
   U16 : XOR2_X1 port map( A => CWP(3), B => n20, Z => n19);
   U17 : XOR2_X1 port map( A => n21, B => n22, Z => n77_port);
   U18 : NAND2_X1 port map( A1 => n23, A2 => n24, ZN => n22);
   U19 : XOR2_X1 port map( A => n9, B => n25, Z => n23);
   U20 : XOR2_X1 port map( A => n26, B => n27, Z => n78_port);
   U21 : NAND2_X1 port map( A1 => n28, A2 => n24, ZN => n27);
   U22 : XOR2_X1 port map( A => n13, B => n29_port, Z => n28);
   U23 : XOR2_X1 port map( A => ADDR_RD2_IN(0), B => n30, Z => n79);
   U24 : NOR2_X1 port map( A1 => n18, A2 => n16, ZN => n30);
   U25 : XOR2_X1 port map( A => ADDR_WR_IN(3), B => n31, Z => n80);
   U26 : NOR2_X1 port map( A1 => n32, A2 => n33, ZN => n31);
   U27 : XOR2_X1 port map( A => CWP(3), B => n34, Z => n33);
   U28 : XOR2_X1 port map( A => n35, B => n36, Z => n81);
   U29 : NAND2_X1 port map( A1 => n37, A2 => n38, ZN => n36);
   U30 : XOR2_X1 port map( A => n9, B => n39, Z => n37);
   U31 : XOR2_X1 port map( A => n40, B => n41, Z => n82);
   U32 : NAND2_X1 port map( A1 => n42, A2 => n38, ZN => n41);
   U33 : XOR2_X1 port map( A => n13, B => n43, Z => n42);
   U34 : INV_X1 port map( A => CWP(1), ZN => n13);
   U35 : XOR2_X1 port map( A => ADDR_WR_IN(0), B => n44, Z => n83);
   U36 : NOR2_X1 port map( A1 => n32, A2 => n16, ZN => n44);
   U37 : INV_X1 port map( A => CWP(0), ZN => n16);
   U38 : AND2_X1 port map( A1 => WR, A2 => ENABLE, ZN => N78);
   U39 : AND2_X1 port map( A1 => RD2, A2 => ENABLE, ZN => N77);
   U40 : AND2_X1 port map( A1 => RD1, A2 => ENABLE, ZN => N76);
   U41 : NOR2_X1 port map( A1 => n32, A2 => n45, ZN => N75);
   U42 : XOR2_X1 port map( A => n46, B => CWP(4), Z => n45);
   U43 : OAI22_X1 port map( A1 => n34, A2 => n47, B1 => n48, B2 => n49, ZN => 
                           n46);
   U44 : AND2_X1 port map( A1 => n47, A2 => n34, ZN => n48);
   U45 : AOI21_X1 port map( B1 => n50, B2 => ADDR_WR_IN(2), A => n51, ZN => n34
                           );
   U46 : AOI21_X1 port map( B1 => n35, B2 => n39, A => n9, ZN => n51);
   U47 : INV_X1 port map( A => n50, ZN => n39);
   U48 : OAI21_X1 port map( B1 => n43, B2 => n40, A => n52_port, ZN => n50);
   U49 : OAI21_X1 port map( B1 => n53, B2 => ADDR_WR_IN(1), A => CWP(1), ZN => 
                           n52_port);
   U50 : INV_X1 port map( A => n43, ZN => n53);
   U51 : INV_X1 port map( A => ADDR_WR_IN(1), ZN => n40);
   U52 : NAND2_X1 port map( A1 => ADDR_WR_IN(0), A2 => CWP(0), ZN => n43);
   U53 : INV_X1 port map( A => n38, ZN => n32);
   U54 : NAND2_X1 port map( A1 => n35, A2 => n47, ZN => n38);
   U55 : INV_X1 port map( A => ADDR_WR_IN(3), ZN => n47);
   U56 : INV_X1 port map( A => ADDR_WR_IN(2), ZN => n35);
   U57 : NOR2_X1 port map( A1 => n18, A2 => n54, ZN => N52);
   U58 : XOR2_X1 port map( A => n55, B => CWP(4), Z => n54);
   U59 : OAI22_X1 port map( A1 => n20, A2 => n56, B1 => n57, B2 => n49, ZN => 
                           n55);
   U60 : INV_X1 port map( A => CWP(3), ZN => n49);
   U61 : AND2_X1 port map( A1 => n56, A2 => n20, ZN => n57);
   U62 : AOI21_X1 port map( B1 => n58, B2 => ADDR_RD2_IN(2), A => n59, ZN => 
                           n20);
   U63 : AOI21_X1 port map( B1 => n21, B2 => n25, A => n9, ZN => n59);
   U64 : INV_X1 port map( A => CWP(2), ZN => n9);
   U65 : INV_X1 port map( A => n58, ZN => n25);
   U66 : OAI21_X1 port map( B1 => n29_port, B2 => n26, A => n60, ZN => n58);
   U67 : OAI21_X1 port map( B1 => n61, B2 => ADDR_RD2_IN(1), A => CWP(1), ZN =>
                           n60);
   U68 : INV_X1 port map( A => n29_port, ZN => n61);
   U69 : INV_X1 port map( A => ADDR_RD2_IN(1), ZN => n26);
   U70 : NAND2_X1 port map( A1 => ADDR_RD2_IN(0), A2 => CWP(0), ZN => n29_port)
                           ;
   U71 : INV_X1 port map( A => n24, ZN => n18);
   U72 : NAND2_X1 port map( A1 => n21, A2 => n56, ZN => n24);
   U73 : INV_X1 port map( A => ADDR_RD2_IN(3), ZN => n56);
   U74 : INV_X1 port map( A => ADDR_RD2_IN(2), ZN => n21);
   U75 : NOR2_X1 port map( A1 => n2, A2 => n62, ZN => N29);
   U76 : XNOR2_X1 port map( A => CWP(4), B => n63, ZN => n62);
   U77 : AOI22_X1 port map( A1 => CWP(3), A2 => n64, B1 => ADDR_RD1_IN(3), B2 
                           => n65, ZN => n63);
   U78 : NAND2_X1 port map( A1 => n4, A2 => n66, ZN => n64);
   U79 : INV_X1 port map( A => n65, ZN => n4);
   U80 : OAI21_X1 port map( B1 => n10, B2 => n5, A => n67, ZN => n65);
   U81 : OAI21_X1 port map( B1 => ADDR_RD1_IN(2), B2 => n68, A => CWP(2), ZN =>
                           n67);
   U82 : INV_X1 port map( A => n10, ZN => n68);
   U83 : AOI21_X1 port map( B1 => n69, B2 => ADDR_RD1_IN(1), A => n70, ZN => 
                           n10);
   U84 : INV_X1 port map( A => n71, ZN => n70);
   U85 : OAI21_X1 port map( B1 => n69, B2 => ADDR_RD1_IN(1), A => CWP(1), ZN =>
                           n71);
   U86 : INV_X1 port map( A => n14, ZN => n69);
   U87 : NAND2_X1 port map( A1 => CWP(0), A2 => ADDR_RD1_IN(0), ZN => n14);
   U88 : INV_X1 port map( A => n8, ZN => n2);
   U89 : NAND2_X1 port map( A1 => n5, A2 => n66, ZN => n8);
   U90 : INV_X1 port map( A => ADDR_RD1_IN(3), ZN => n66);
   U91 : INV_X1 port map( A => ADDR_RD1_IN(2), ZN => n5);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_entity.all;

entity window_reg_fsm_Nbit32_M4_N4_F3_bit_F2_IN_LOC8_bit_inloc3 is

   port( Clk, Rst, CALL, RET, ACK_FILL, ACK_SPILL : in std_logic;  FILL, SPILL 
         : out std_logic;  CWP, SWP : out std_logic_vector (4 downto 0));

end window_reg_fsm_Nbit32_M4_N4_F3_bit_F2_IN_LOC8_bit_inloc3;

architecture SYN_Behavioral of 
   window_reg_fsm_Nbit32_M4_N4_F3_bit_F2_IN_LOC8_bit_inloc3 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal FILL_port, SPILL_port, N160, N161, n56, n57, n58, n59, n60, n61, n62,
      n63, n64, n65, n66, n69, n73, n74, n75, n132, n133, n134, n135, n136, 
      n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, 
      n149, n150, n151, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
      n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28
      , n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, 
      n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n67, n68
      , n70, n71, n72, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, 
      n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, 
      n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, 
      n113, n114, n115, n116, n117, n118, n119, n_2088, n_2089, n_2090, n_2091,
      n_2092, n_2093, n_2094 : std_logic;

begin
   FILL <= FILL_port;
   SPILL <= SPILL_port;
   
   TransferRegsCounter_reg_0_inst : DFF_X1 port map( D => n151, CK => n9, Q => 
                           n_2088, QN => n75);
   TransferRegsCounter_reg_2_inst : DFF_X1 port map( D => n150, CK => n9, Q => 
                           n_2089, QN => n73);
   CurrState_reg_1_inst : DFFR_X1 port map( D => N161, CK => n9, RN => n119, Q 
                           => n8, QN => n56);
   CurrState_reg_0_inst : DFFR_X1 port map( D => N160, CK => n9, RN => n119, Q 
                           => n_2090, QN => n114);
   TransferRegsCounter_reg_1_inst : DFF_X1 port map( D => n141, CK => n9, Q => 
                           n7, QN => n74);
   cwp_s_reg_4_inst : DFF_X1 port map( D => n149, CK => n11, Q => CWP(4), QN =>
                           n62);
   swp_s_reg_0_inst : DFF_X1 port map( D => n140, CK => n10, Q => SWP(0), QN =>
                           n61);
   swp_s_reg_1_inst : DFF_X1 port map( D => n139, CK => n10, Q => SWP(1), QN =>
                           n60);
   swp_s_reg_2_inst : DFF_X1 port map( D => n138, CK => n10, Q => SWP(2), QN =>
                           n59);
   cwp_s_reg_3_inst : DFF_X1 port map( D => n133, CK => n9, Q => CWP(3), QN => 
                           n63);
   cwp_s_reg_0_inst : DFF_X1 port map( D => n136, CK => n9, Q => CWP(0), QN => 
                           n66);
   cwp_s_reg_1_inst : DFF_X1 port map( D => n135, CK => n9, Q => CWP(1), QN => 
                           n65);
   CANRESTORE_reg_2_inst : DFF_X1 port map( D => n147, CK => n10, Q => n116, QN
                           => n3);
   CANSAVE_reg_0_inst : DFF_X1 port map( D => n143, CK => n10, Q => n6, QN => 
                           n69);
   CANSAVE_reg_1_inst : DFF_X1 port map( D => n144, CK => n10, Q => n_2091, QN 
                           => n2);
   CANSAVE_reg_2_inst : DFF_X1 port map( D => n142, CK => n10, Q => n_2092, QN 
                           => n4);
   CANRESTORE_reg_0_inst : DFF_X1 port map( D => n145, CK => n10, Q => n115, QN
                           => n1);
   CANRESTORE_reg_1_inst : DFF_X1 port map( D => n146, CK => n9, Q => n117, QN 
                           => n5);
   cwp_s_reg_2_inst : DFF_X1 port map( D => n134, CK => n10, Q => CWP(2), QN =>
                           n64);
   swp_s_reg_3_inst : DFF_X1 port map( D => n137, CK => n9, Q => SWP(3), QN => 
                           n58);
   swp_s_reg_4_inst : DFF_X1 port map( D => n148, CK => n10, Q => SWP(4), QN =>
                           n57);
   FILL_reg : DFF_X1 port map( D => n118, CK => n10, Q => FILL_port, QN => 
                           n_2093);
   SPILL_reg : DFF_X1 port map( D => n132, CK => n9, Q => SPILL_port, QN => 
                           n_2094);
   U3 : BUF_X1 port map( A => Clk, Z => n11);
   U4 : BUF_X1 port map( A => n11, Z => n9);
   U5 : BUF_X1 port map( A => n11, Z => n10);
   U6 : MUX2_X1 port map( A => FILL_port, B => n12, S => n13, Z => n118);
   U7 : NOR2_X1 port map( A1 => n14, A2 => Rst, ZN => n13);
   U8 : AOI21_X1 port map( B1 => n15, B2 => n16, A => n17, ZN => n14);
   U9 : MUX2_X1 port map( A => n18, B => n19, S => n75, Z => n151);
   U10 : NOR2_X1 port map( A1 => n18, A2 => n20, ZN => n19);
   U11 : INV_X1 port map( A => n21, ZN => n150);
   U12 : AOI21_X1 port map( B1 => n7, B2 => n22, A => n23, ZN => n21);
   U13 : AOI21_X1 port map( B1 => n20, B2 => n24, A => n73, ZN => n23);
   U14 : INV_X1 port map( A => n18, ZN => n24);
   U15 : OAI221_X1 port map( B1 => n25, B2 => n26, C1 => n62, C2 => n27, A => 
                           n28, ZN => n149);
   U16 : INV_X1 port map( A => n29, ZN => n28);
   U17 : OAI21_X1 port map( B1 => n30, B2 => n31, A => n32, ZN => n29);
   U18 : XOR2_X1 port map( A => n62, B => n63, Z => n31);
   U19 : NAND2_X1 port map( A1 => n33, A2 => n34, ZN => n148);
   U20 : MUX2_X1 port map( A => n25, B => n57, S => n35, Z => n33);
   U21 : XNOR2_X1 port map( A => n36, B => n37, ZN => n25);
   U22 : XOR2_X1 port map( A => n38, B => n39, Z => n37);
   U23 : OAI21_X1 port map( B1 => n40, B2 => n41, A => n42, ZN => n39);
   U24 : OAI22_X1 port map( A1 => n57, A2 => n43, B1 => n62, B2 => n44, ZN => 
                           n36);
   U25 : OAI22_X1 port map( A1 => n45, A2 => n3, B1 => n46, B2 => n47, ZN => 
                           n147);
   U26 : XOR2_X1 port map( A => n48, B => n49, Z => n47);
   U27 : XNOR2_X1 port map( A => n50, B => n3, ZN => n49);
   U28 : OAI22_X1 port map( A1 => n5, A2 => n1, B1 => n51, B2 => n50, ZN => n48
                           );
   U29 : NOR2_X1 port map( A1 => n115, A2 => n117, ZN => n51);
   U30 : OAI22_X1 port map( A1 => n45, A2 => n5, B1 => n46, B2 => n52, ZN => 
                           n146);
   U31 : XOR2_X1 port map( A => n50, B => n53, Z => n52);
   U32 : XNOR2_X1 port map( A => n1, B => n117, ZN => n53);
   U33 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n115, B2 => n46, ZN => 
                           n145);
   U34 : OAI21_X1 port map( B1 => n54, B2 => n46, A => n55, ZN => n144);
   U35 : MUX2_X1 port map( A => n67, B => n2, S => n68, Z => n55);
   U36 : AOI21_X1 port map( B1 => n70, B2 => n40, A => n71, ZN => n54);
   U37 : OAI21_X1 port map( B1 => n6, B2 => n46, A => n72, ZN => n143);
   U38 : MUX2_X1 port map( A => n67, B => n69, S => n68, Z => n72);
   U39 : MUX2_X1 port map( A => n76, B => n77, S => n4, Z => n142);
   U40 : NOR4_X1 port map( A1 => n69, A2 => n78, A3 => n46, A4 => n2, ZN => n77
                           );
   U41 : NAND2_X1 port map( A1 => n45, A2 => n12, ZN => n46);
   U42 : OAI21_X1 port map( B1 => n41, B2 => n79, A => n45, ZN => n76);
   U43 : INV_X1 port map( A => n68, ZN => n45);
   U44 : OAI21_X1 port map( B1 => n80, B2 => n81, A => n119, ZN => n68);
   U45 : MUX2_X1 port map( A => n71, B => n40, S => n82, Z => n79);
   U46 : NOR2_X1 port map( A1 => n69, A2 => n2, ZN => n82);
   U47 : NOR2_X1 port map( A1 => n40, A2 => n70, ZN => n71);
   U48 : XNOR2_X1 port map( A => n6, B => n2, ZN => n70);
   U49 : MUX2_X1 port map( A => n22, B => n83, S => n7, Z => n141);
   U50 : INV_X1 port map( A => n84, ZN => n83);
   U51 : AOI21_X1 port map( B1 => n85, B2 => n75, A => n18, ZN => n84);
   U52 : NOR3_X1 port map( A1 => n18, A2 => n75, A3 => n20, ZN => n22);
   U53 : NAND2_X1 port map( A1 => n119, A2 => n86, ZN => n18);
   U54 : NAND3_X1 port map( A1 => n20, A2 => n67, A3 => n87, ZN => n86);
   U55 : NAND2_X1 port map( A1 => n61, A2 => n34, ZN => n140);
   U56 : NAND2_X1 port map( A1 => n60, A2 => n34, ZN => n139);
   U57 : NAND2_X1 port map( A1 => n59, A2 => n34, ZN => n138);
   U58 : NAND2_X1 port map( A1 => n88, A2 => n80, ZN => n34);
   U59 : INV_X1 port map( A => n89, ZN => n137);
   U60 : MUX2_X1 port map( A => n38, B => n58, S => n35, Z => n89);
   U61 : NAND2_X1 port map( A1 => n66, A2 => n32, ZN => n136);
   U62 : NAND2_X1 port map( A1 => n65, A2 => n32, ZN => n135);
   U63 : NAND2_X1 port map( A1 => n64, A2 => n32, ZN => n134);
   U64 : OAI211_X1 port map( C1 => n38, C2 => n26, A => n32, B => n90, ZN => 
                           n133);
   U65 : MUX2_X1 port map( A => n27, B => n30, S => n63, Z => n90);
   U66 : NAND2_X1 port map( A1 => n27, A2 => n91, ZN => n30);
   U67 : NAND2_X1 port map( A1 => n80, A2 => n27, ZN => n32);
   U68 : INV_X1 port map( A => n67, ZN => n80);
   U69 : NAND2_X1 port map( A1 => n12, A2 => n27, ZN => n26);
   U70 : NAND2_X1 port map( A1 => n35, A2 => n92, ZN => n27);
   U71 : OR3_X1 port map( A1 => n93, A2 => Rst, A3 => n41, ZN => n92);
   U72 : AOI21_X1 port map( B1 => n94, B2 => RET, A => n78, ZN => n93);
   U73 : INV_X1 port map( A => n40, ZN => n78);
   U74 : INV_X1 port map( A => n88, ZN => n35);
   U75 : AOI21_X1 port map( B1 => n43, B2 => n67, A => Rst, ZN => n88);
   U76 : OAI22_X1 port map( A1 => n58, A2 => n43, B1 => n63, B2 => n44, ZN => 
                           n38);
   U77 : NOR2_X1 port map( A1 => n81, A2 => n16, ZN => n44);
   U78 : OAI21_X1 port map( B1 => n41, B2 => n40, A => n50, ZN => n81);
   U79 : NAND4_X1 port map( A1 => RET, A2 => n12, A3 => n95, A4 => n94, ZN => 
                           n50);
   U80 : NAND3_X1 port map( A1 => n3, A2 => n1, A3 => n5, ZN => n95);
   U81 : NAND2_X1 port map( A1 => CALL, A2 => n96, ZN => n40);
   U82 : NAND3_X1 port map( A1 => n2, A2 => n4, A3 => n69, ZN => n96);
   U83 : OR2_X1 port map( A1 => n97, A2 => n87, ZN => n43);
   U84 : AOI22_X1 port map( A1 => n98, A2 => ACK_SPILL, B1 => n17, B2 => 
                           ACK_FILL, ZN => n87);
   U85 : MUX2_X1 port map( A => n12, B => SPILL_port, S => n99, Z => n132);
   U86 : OAI21_X1 port map( B1 => n100, B2 => n98, A => n119, ZN => n99);
   U87 : INV_X1 port map( A => Rst, ZN => n119);
   U88 : OAI221_X1 port map( B1 => ACK_FILL, B2 => n101, C1 => ACK_SPILL, C2 =>
                           n102, A => n103, ZN => N161);
   U89 : AOI211_X1 port map( C1 => n15, C2 => n16, A => n100, B => n85, ZN => 
                           n103);
   U90 : INV_X1 port map( A => n20, ZN => n85);
   U91 : NAND2_X1 port map( A1 => n91, A2 => n97, ZN => n20);
   U92 : INV_X1 port map( A => n104, ZN => n97);
   U93 : NAND2_X1 port map( A1 => n102, A2 => n101, ZN => n91);
   U94 : NOR2_X1 port map( A1 => n105, A2 => n41, ZN => n100);
   U95 : INV_X1 port map( A => n12, ZN => n41);
   U96 : AND4_X1 port map( A1 => n12, A2 => n94, A3 => RET, A4 => n106, ZN => 
                           n16);
   U97 : NOR3_X1 port map( A1 => n117, A2 => n115, A3 => n116, ZN => n106);
   U98 : INV_X1 port map( A => CALL, ZN => n94);
   U99 : AND4_X1 port map( A1 => n107, A2 => n108, A3 => n109, A4 => n110, ZN 
                           => n15);
   U100 : NOR2_X1 port map( A1 => n111, A2 => n112, ZN => n110);
   U101 : XOR2_X1 port map( A => n62, B => n57, Z => n112);
   U102 : XOR2_X1 port map( A => n66, B => n61, Z => n111);
   U103 : XNOR2_X1 port map( A => n59, B => n64, ZN => n109);
   U104 : XNOR2_X1 port map( A => n60, B => n65, ZN => n108);
   U105 : XNOR2_X1 port map( A => n58, B => n63, ZN => n107);
   U106 : NAND4_X1 port map( A1 => n113, A2 => n101, A3 => n42, A4 => n67, ZN 
                           => N160);
   U107 : NAND2_X1 port map( A1 => n114, A2 => n56, ZN => n67);
   U108 : NAND3_X1 port map( A1 => ACK_SPILL, A2 => n98, A3 => n104, ZN => n42)
                           ;
   U109 : NOR3_X1 port map( A1 => n74, A2 => n75, A3 => n73, ZN => n104);
   U110 : INV_X1 port map( A => n102, ZN => n98);
   U111 : NAND2_X1 port map( A1 => n114, A2 => n8, ZN => n102);
   U112 : INV_X1 port map( A => n17, ZN => n101);
   U113 : NOR2_X1 port map( A1 => n114, A2 => n56, ZN => n17);
   U114 : NAND2_X1 port map( A1 => n12, A2 => n105, ZN => n113);
   U115 : NAND4_X1 port map( A1 => CALL, A2 => n69, A3 => n2, A4 => n4, ZN => 
                           n105);
   U116 : NOR2_X1 port map( A1 => n8, A2 => n114, ZN => n12);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_entity.all;

entity top_entity is

   port( Clk, Rst, CALL, RET, ACK_FILL, ACK_SPILL : in std_logic;  FILL, SPILL 
         : out std_logic;  CWP, SWP : out std_logic_vector (4 downto 0);  
         ENABLE, RD1, RD2, WR : in std_logic;  ADDR_WR_IN, ADDR_RD1_IN, 
         ADDR_RD2_IN : in std_logic_vector (3 downto 0);  DATAIN : in 
         std_logic_vector (31 downto 0);  OUT1, OUT2 : out std_logic_vector (31
         downto 0));

end top_entity;

architecture SYN_structural of top_entity is

   component register_file_nbit32_addr_bits5
      port( CLK, RESET, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
            ADD_RD2 : in std_logic_vector (4 downto 0);  DATAIN : in 
            std_logic_vector (31 downto 0);  OUT1, OUT2 : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component Addr_Transformer_Addr_bits5_M4_in_loc_out12
      port( ENABLE, RD1, RD2, WR : in std_logic;  ADDR_WR_IN, ADDR_RD1_IN, 
            ADDR_RD2_IN : in std_logic_vector (3 downto 0);  CWP : in 
            std_logic_vector (4 downto 0);  ADDR_WR_OUT, ADDR_RD1_OUT, 
            ADDR_RD2_OUT : out std_logic_vector (4 downto 0));
   end component;
   
   component window_reg_fsm_Nbit32_M4_N4_F3_bit_F2_IN_LOC8_bit_inloc3
      port( Clk, Rst, CALL, RET, ACK_FILL, ACK_SPILL : in std_logic;  FILL, 
            SPILL : out std_logic;  CWP, SWP : out std_logic_vector (4 downto 
            0));
   end component;
   
   signal cwp_s_4_port, cwp_s_3_port, cwp_s_2_port, cwp_s_1_port, cwp_s_0_port,
      ADDR_WR_4_port, ADDR_WR_3_port, ADDR_WR_2_port, ADDR_WR_1_port, 
      ADDR_WR_0_port, ADDR_RD1_4_port, ADDR_RD1_3_port, ADDR_RD1_2_port, 
      ADDR_RD1_1_port, ADDR_RD1_0_port, ADDR_RD2_4_port, ADDR_RD2_3_port, 
      ADDR_RD2_2_port, ADDR_RD2_1_port, ADDR_RD2_0_port, n_2107, n_2108, n_2109
      , n_2110, n_2111, n_2112, n_2113 : std_logic;

begin
   
   fsm : window_reg_fsm_Nbit32_M4_N4_F3_bit_F2_IN_LOC8_bit_inloc3 port map( Clk
                           => Clk, Rst => Rst, CALL => CALL, RET => RET, 
                           ACK_FILL => ACK_FILL, ACK_SPILL => ACK_SPILL, FILL 
                           => n_2107, SPILL => n_2108, CWP(4) => cwp_s_4_port, 
                           CWP(3) => cwp_s_3_port, CWP(2) => cwp_s_2_port, 
                           CWP(1) => cwp_s_1_port, CWP(0) => cwp_s_0_port, 
                           SWP(4) => n_2109, SWP(3) => n_2110, SWP(2) => n_2111
                           , SWP(1) => n_2112, SWP(0) => n_2113);
   addr_trsf : Addr_Transformer_Addr_bits5_M4_in_loc_out12 port map( ENABLE => 
                           ENABLE, RD1 => RD1, RD2 => RD2, WR => WR, 
                           ADDR_WR_IN(3) => ADDR_WR_IN(3), ADDR_WR_IN(2) => 
                           ADDR_WR_IN(2), ADDR_WR_IN(1) => ADDR_WR_IN(1), 
                           ADDR_WR_IN(0) => ADDR_WR_IN(0), ADDR_RD1_IN(3) => 
                           ADDR_RD1_IN(3), ADDR_RD1_IN(2) => ADDR_RD1_IN(2), 
                           ADDR_RD1_IN(1) => ADDR_RD1_IN(1), ADDR_RD1_IN(0) => 
                           ADDR_RD1_IN(0), ADDR_RD2_IN(3) => ADDR_RD2_IN(3), 
                           ADDR_RD2_IN(2) => ADDR_RD2_IN(2), ADDR_RD2_IN(1) => 
                           ADDR_RD2_IN(1), ADDR_RD2_IN(0) => ADDR_RD2_IN(0), 
                           CWP(4) => cwp_s_4_port, CWP(3) => cwp_s_3_port, 
                           CWP(2) => cwp_s_2_port, CWP(1) => cwp_s_1_port, 
                           CWP(0) => cwp_s_0_port, ADDR_WR_OUT(4) => 
                           ADDR_WR_4_port, ADDR_WR_OUT(3) => ADDR_WR_3_port, 
                           ADDR_WR_OUT(2) => ADDR_WR_2_port, ADDR_WR_OUT(1) => 
                           ADDR_WR_1_port, ADDR_WR_OUT(0) => ADDR_WR_0_port, 
                           ADDR_RD1_OUT(4) => ADDR_RD1_4_port, ADDR_RD1_OUT(3) 
                           => ADDR_RD1_3_port, ADDR_RD1_OUT(2) => 
                           ADDR_RD1_2_port, ADDR_RD1_OUT(1) => ADDR_RD1_1_port,
                           ADDR_RD1_OUT(0) => ADDR_RD1_0_port, ADDR_RD2_OUT(4) 
                           => ADDR_RD2_4_port, ADDR_RD2_OUT(3) => 
                           ADDR_RD2_3_port, ADDR_RD2_OUT(2) => ADDR_RD2_2_port,
                           ADDR_RD2_OUT(1) => ADDR_RD2_1_port, ADDR_RD2_OUT(0) 
                           => ADDR_RD2_0_port);
   regfile : register_file_nbit32_addr_bits5 port map( CLK => Clk, RESET => Rst
                           , ENABLE => ENABLE, RD1 => RD1, RD2 => RD2, WR => WR
                           , ADD_WR(4) => ADDR_WR_4_port, ADD_WR(3) => 
                           ADDR_WR_3_port, ADD_WR(2) => ADDR_WR_2_port, 
                           ADD_WR(1) => ADDR_WR_1_port, ADD_WR(0) => 
                           ADDR_WR_0_port, ADD_RD1(4) => ADDR_RD1_4_port, 
                           ADD_RD1(3) => ADDR_RD1_3_port, ADD_RD1(2) => 
                           ADDR_RD1_2_port, ADD_RD1(1) => ADDR_RD1_1_port, 
                           ADD_RD1(0) => ADDR_RD1_0_port, ADD_RD2(4) => 
                           ADDR_RD2_4_port, ADD_RD2(3) => ADDR_RD2_3_port, 
                           ADD_RD2(2) => ADDR_RD2_2_port, ADD_RD2(1) => 
                           ADDR_RD2_1_port, ADD_RD2(0) => ADDR_RD2_0_port, 
                           DATAIN(31) => DATAIN(31), DATAIN(30) => DATAIN(30), 
                           DATAIN(29) => DATAIN(29), DATAIN(28) => DATAIN(28), 
                           DATAIN(27) => DATAIN(27), DATAIN(26) => DATAIN(26), 
                           DATAIN(25) => DATAIN(25), DATAIN(24) => DATAIN(24), 
                           DATAIN(23) => DATAIN(23), DATAIN(22) => DATAIN(22), 
                           DATAIN(21) => DATAIN(21), DATAIN(20) => DATAIN(20), 
                           DATAIN(19) => DATAIN(19), DATAIN(18) => DATAIN(18), 
                           DATAIN(17) => DATAIN(17), DATAIN(16) => DATAIN(16), 
                           DATAIN(15) => DATAIN(15), DATAIN(14) => DATAIN(14), 
                           DATAIN(13) => DATAIN(13), DATAIN(12) => DATAIN(12), 
                           DATAIN(11) => DATAIN(11), DATAIN(10) => DATAIN(10), 
                           DATAIN(9) => DATAIN(9), DATAIN(8) => DATAIN(8), 
                           DATAIN(7) => DATAIN(7), DATAIN(6) => DATAIN(6), 
                           DATAIN(5) => DATAIN(5), DATAIN(4) => DATAIN(4), 
                           DATAIN(3) => DATAIN(3), DATAIN(2) => DATAIN(2), 
                           DATAIN(1) => DATAIN(1), DATAIN(0) => DATAIN(0), 
                           OUT1(31) => OUT1(31), OUT1(30) => OUT1(30), OUT1(29)
                           => OUT1(29), OUT1(28) => OUT1(28), OUT1(27) => 
                           OUT1(27), OUT1(26) => OUT1(26), OUT1(25) => OUT1(25)
                           , OUT1(24) => OUT1(24), OUT1(23) => OUT1(23), 
                           OUT1(22) => OUT1(22), OUT1(21) => OUT1(21), OUT1(20)
                           => OUT1(20), OUT1(19) => OUT1(19), OUT1(18) => 
                           OUT1(18), OUT1(17) => OUT1(17), OUT1(16) => OUT1(16)
                           , OUT1(15) => OUT1(15), OUT1(14) => OUT1(14), 
                           OUT1(13) => OUT1(13), OUT1(12) => OUT1(12), OUT1(11)
                           => OUT1(11), OUT1(10) => OUT1(10), OUT1(9) => 
                           OUT1(9), OUT1(8) => OUT1(8), OUT1(7) => OUT1(7), 
                           OUT1(6) => OUT1(6), OUT1(5) => OUT1(5), OUT1(4) => 
                           OUT1(4), OUT1(3) => OUT1(3), OUT1(2) => OUT1(2), 
                           OUT1(1) => OUT1(1), OUT1(0) => OUT1(0), OUT2(31) => 
                           OUT2(31), OUT2(30) => OUT2(30), OUT2(29) => OUT2(29)
                           , OUT2(28) => OUT2(28), OUT2(27) => OUT2(27), 
                           OUT2(26) => OUT2(26), OUT2(25) => OUT2(25), OUT2(24)
                           => OUT2(24), OUT2(23) => OUT2(23), OUT2(22) => 
                           OUT2(22), OUT2(21) => OUT2(21), OUT2(20) => OUT2(20)
                           , OUT2(19) => OUT2(19), OUT2(18) => OUT2(18), 
                           OUT2(17) => OUT2(17), OUT2(16) => OUT2(16), OUT2(15)
                           => OUT2(15), OUT2(14) => OUT2(14), OUT2(13) => 
                           OUT2(13), OUT2(12) => OUT2(12), OUT2(11) => OUT2(11)
                           , OUT2(10) => OUT2(10), OUT2(9) => OUT2(9), OUT2(8) 
                           => OUT2(8), OUT2(7) => OUT2(7), OUT2(6) => OUT2(6), 
                           OUT2(5) => OUT2(5), OUT2(4) => OUT2(4), OUT2(3) => 
                           OUT2(3), OUT2(2) => OUT2(2), OUT2(1) => OUT2(1), 
                           OUT2(0) => OUT2(0));

end SYN_structural;
