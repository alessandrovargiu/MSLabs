
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_BOOTHMUL is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_BOOTHMUL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_1022 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1022;

architecture SYN_BEHAVIORAL of FA_1022 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n6, n7, n8, n9, n10 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => n9);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => n6);
   U3 : BUF_X1 port map( A => Ci, Z => n10);
   U4 : AOI21_X1 port map( B1 => Ci, B2 => n8, A => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : INV_X1 port map( A => n9, ZN => n8);
   U7 : XNOR2_X1 port map( A => n10, B => n9, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_1021 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1021;

architecture SYN_BEHAVIORAL of FA_1021 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U2 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_1020 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1020;

architecture SYN_BEHAVIORAL of FA_1020 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n6, n7, n9, n10, n11, n12, n14 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n14);
   U2 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => Ci, A2 => n14, ZN => n7);
   U4 : NAND2_X1 port map( A1 => n6, A2 => n7, ZN => Co);
   U5 : OR2_X1 port map( A1 => Ci, A2 => n9, ZN => n12);
   U6 : INV_X1 port map( A => n14, ZN => n9);
   U7 : NAND2_X1 port map( A1 => n12, A2 => n11, ZN => S);
   U8 : NAND2_X1 port map( A1 => Ci, A2 => n10, ZN => n11);
   U9 : INV_X1 port map( A => n14, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_1019 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1019;

architecture SYN_BEHAVIORAL of FA_1019 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n6, n7, n8, n9, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : OAI22_X1 port map( A1 => n6, A2 => n7, B1 => n8, B2 => n9, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n6);
   U5 : INV_X1 port map( A => A, ZN => n7);
   U6 : INV_X1 port map( A => Ci, ZN => n8);
   U7 : INV_X1 port map( A => n11, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_1018 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1018;

architecture SYN_BEHAVIORAL of FA_1018 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n6, n7, n8, n9, n11 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : OAI22_X1 port map( A1 => n6, A2 => n7, B1 => n8, B2 => n9, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n6);
   U5 : INV_X1 port map( A => A, ZN => n7);
   U6 : INV_X1 port map( A => Ci, ZN => n8);
   U7 : INV_X1 port map( A => n11, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_1017 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1017;

architecture SYN_BEHAVIORAL of FA_1017 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n6, n7, n8 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => n8);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => n6);
   U3 : AOI21_X1 port map( B1 => Ci, B2 => n7, A => n6, ZN => n2);
   U4 : INV_X1 port map( A => n8, ZN => n7);
   U5 : XNOR2_X1 port map( A => Ci, B => n8, ZN => S);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_1016 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1016;

architecture SYN_BEHAVIORAL of FA_1016 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n6, n8, n9 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n8);
   U1 : INV_X1 port map( A => n8, ZN => n6);
   U2 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n8, ZN => n9);
   U5 : INV_X1 port map( A => n9, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_1015 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1015;

architecture SYN_BEHAVIORAL of FA_1015 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);
   U1 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : INV_X1 port map( A => n8, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_1014 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1014;

architecture SYN_BEHAVIORAL of FA_1014 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n6, n7, n9 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => n9, ZN => n7);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n9, ZN => n6);
   U3 : INV_X1 port map( A => n6, ZN => Co);
   U5 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_1013 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1013;

architecture SYN_BEHAVIORAL of FA_1013 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n6, n8, n9 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n8);
   U1 : INV_X1 port map( A => n8, ZN => n6);
   U2 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n8, ZN => n9);
   U5 : INV_X1 port map( A => n9, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_1012 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1012;

architecture SYN_BEHAVIORAL of FA_1012 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);
   U1 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : INV_X1 port map( A => n8, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_1011 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1011;

architecture SYN_BEHAVIORAL of FA_1011 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);
   U1 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U3 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_1010 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1010;

architecture SYN_BEHAVIORAL of FA_1010 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n6, n8, n9 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n8);
   U1 : INV_X1 port map( A => n8, ZN => n6);
   U2 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);
   U3 : INV_X1 port map( A => n9, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n8, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_1009 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1009;

architecture SYN_BEHAVIORAL of FA_1009 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);
   U1 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U3 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_1008 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1008;

architecture SYN_BEHAVIORAL of FA_1008 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);
   U1 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U3 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_1007 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1007;

architecture SYN_BEHAVIORAL of FA_1007 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);
   U1 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : INV_X1 port map( A => n8, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n7, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_1006 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1006;

architecture SYN_BEHAVIORAL of FA_1006 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n6, n8, n9 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);
   U2 : XOR2_X1 port map( A => A, B => B, Z => n8);
   U3 : INV_X1 port map( A => n8, ZN => n6);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n8, ZN => n9);
   U5 : INV_X1 port map( A => n9, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_1005 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1005;

architecture SYN_BEHAVIORAL of FA_1005 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);
   U1 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : INV_X1 port map( A => n8, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_1004 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1004;

architecture SYN_BEHAVIORAL of FA_1004 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);
   U1 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n7, B2 => Ci, ZN => n8);
   U3 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_1003 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1003;

architecture SYN_BEHAVIORAL of FA_1003 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X2
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n6, n8, n9 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n8);
   U1 : INV_X1 port map( A => n8, ZN => n6);
   U2 : XNOR2_X2 port map( A => Ci, B => n6, ZN => S);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n8, B2 => Ci, ZN => n9);
   U5 : INV_X1 port map( A => n9, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_1002 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1002;

architecture SYN_BEHAVIORAL of FA_1002 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);
   U1 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : INV_X1 port map( A => n8, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n7, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_1001 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1001;

architecture SYN_BEHAVIORAL of FA_1001 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);
   U1 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n7, B2 => Ci, ZN => n8);
   U3 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_1000 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1000;

architecture SYN_BEHAVIORAL of FA_1000 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);
   U1 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : INV_X1 port map( A => n8, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n7, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_999 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_999;

architecture SYN_BEHAVIORAL of FA_999 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);
   U1 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n7, B2 => Ci, ZN => n8);
   U3 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_998 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_998;

architecture SYN_BEHAVIORAL of FA_998 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);
   U1 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U3 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_997 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_997;

architecture SYN_BEHAVIORAL of FA_997 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);
   U1 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : INV_X1 port map( A => n8, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n7, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_996 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_996;

architecture SYN_BEHAVIORAL of FA_996 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);
   U1 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n7, B2 => Ci, ZN => n8);
   U3 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_995 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_995;

architecture SYN_BEHAVIORAL of FA_995 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);
   U1 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : INV_X1 port map( A => n8, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n7, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_994 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_994;

architecture SYN_BEHAVIORAL of FA_994 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);
   U1 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n7, B2 => Ci, ZN => n8);
   U3 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_993 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_993;

architecture SYN_BEHAVIORAL of FA_993 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);
   U1 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n7, B2 => Ci, ZN => n8);
   U3 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_992 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_992;

architecture SYN_BEHAVIORAL of FA_992 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);
   U1 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : INV_X1 port map( A => n8, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_991 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_991;

architecture SYN_BEHAVIORAL of FA_991 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);
   U1 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n7, B2 => Ci, ZN => n8);
   U3 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_990 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_990;

architecture SYN_BEHAVIORAL of FA_990 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);
   U1 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : INV_X1 port map( A => n8, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n7, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_989 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_989;

architecture SYN_BEHAVIORAL of FA_989 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);
   U1 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n7, B2 => Ci, ZN => n8);
   U3 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_988 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_988;

architecture SYN_BEHAVIORAL of FA_988 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);
   U1 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n7, B2 => Ci, ZN => n8);
   U3 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_987 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_987;

architecture SYN_BEHAVIORAL of FA_987 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);
   U1 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : INV_X1 port map( A => n8, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n7, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_986 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_986;

architecture SYN_BEHAVIORAL of FA_986 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);
   U1 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : INV_X1 port map( A => n8, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n7, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_984 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_984;

architecture SYN_BEHAVIORAL of FA_984 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);
   U1 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : INV_X1 port map( A => n8, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n7, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_983 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_983;

architecture SYN_BEHAVIORAL of FA_983 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n7, n8, n9 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n8);
   U1 : INV_X2 port map( A => n7, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => n8, ZN => n7);
   U3 : INV_X1 port map( A => n9, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n8, B2 => Ci, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_982 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_982;

architecture SYN_BEHAVIORAL of FA_982 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n7, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_980 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_980;

architecture SYN_BEHAVIORAL of FA_980 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n9 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n8);
   U1 : NAND2_X1 port map( A1 => Ci, A2 => n7, ZN => n5);
   U2 : NAND2_X1 port map( A1 => n4, A2 => n8, ZN => n6);
   U3 : NAND2_X4 port map( A1 => n5, A2 => n6, ZN => S);
   U5 : INV_X1 port map( A => Ci, ZN => n4);
   U6 : INV_X1 port map( A => n8, ZN => n7);
   U7 : INV_X1 port map( A => n9, ZN => Co);
   U8 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n8, B2 => Ci, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_979 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_979;

architecture SYN_BEHAVIORAL of FA_979 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);
   U3 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_978 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_978;

architecture SYN_BEHAVIORAL of FA_978 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);
   U3 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_977 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_977;

architecture SYN_BEHAVIORAL of FA_977 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U2 : INV_X1 port map( A => n5, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_976 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_976;

architecture SYN_BEHAVIORAL of FA_976 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n5, n6 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : BUF_X2 port map( A => n8, Z => S);
   U2 : XOR2_X1 port map( A => Ci, B => n5, Z => n8);
   U3 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_975 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_975;

architecture SYN_BEHAVIORAL of FA_975 is

   component XOR2_X2
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);
   U3 : XOR2_X2 port map( A => Ci, B => n4, Z => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_974 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_974;

architecture SYN_BEHAVIORAL of FA_974 is

   component XOR2_X2
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);
   U3 : XOR2_X2 port map( A => Ci, B => n4, Z => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_973 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_973;

architecture SYN_BEHAVIORAL of FA_973 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X2
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : XOR2_X2 port map( A => Ci, B => n4, Z => S);
   U2 : INV_X1 port map( A => n5, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_972 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_972;

architecture SYN_BEHAVIORAL of FA_972 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X2
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : XOR2_X2 port map( A => Ci, B => n4, Z => S);
   U2 : INV_X1 port map( A => n5, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_970 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_970;

architecture SYN_BEHAVIORAL of FA_970 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X2
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : XOR2_X2 port map( A => Ci, B => n4, Z => S);
   U2 : INV_X1 port map( A => n5, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_969 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_969;

architecture SYN_BEHAVIORAL of FA_969 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_968 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_968;

architecture SYN_BEHAVIORAL of FA_968 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_967 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_967;

architecture SYN_BEHAVIORAL of FA_967 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_966 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_966;

architecture SYN_BEHAVIORAL of FA_966 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_965 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_965;

architecture SYN_BEHAVIORAL of FA_965 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_964 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_964;

architecture SYN_BEHAVIORAL of FA_964 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_963 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_963;

architecture SYN_BEHAVIORAL of FA_963 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_962 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_962;

architecture SYN_BEHAVIORAL of FA_962 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_961 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_961;

architecture SYN_BEHAVIORAL of FA_961 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_960 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_960;

architecture SYN_BEHAVIORAL of FA_960 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_959 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_959;

architecture SYN_BEHAVIORAL of FA_959 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_958 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_958;

architecture SYN_BEHAVIORAL of FA_958 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_957 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_957;

architecture SYN_BEHAVIORAL of FA_957 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal net156153, n2, n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => net156153, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => n5, B1 => n4, B2 => Ci, ZN => n2);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U5 : CLKBUF_X1 port map( A => A, Z => n5);
   U6 : CLKBUF_X1 port map( A => n4, Z => net156153);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_956 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_956;

architecture SYN_BEHAVIORAL of FA_956 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal net154989, net156164, n2, n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => net154989, B => net156164, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => n5, B1 => Ci, B2 => n4, ZN => n2);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U5 : CLKBUF_X1 port map( A => A, Z => n5);
   U6 : CLKBUF_X1 port map( A => Ci, Z => net156164);
   U7 : CLKBUF_X1 port map( A => n4, Z => net154989);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_955 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_955;

architecture SYN_BEHAVIORAL of FA_955 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U2 : INV_X1 port map( A => n4, ZN => n8);
   U5 : OAI22_X1 port map( A1 => n5, A2 => n6, B1 => n7, B2 => n8, ZN => Co);
   U6 : INV_X1 port map( A => B, ZN => n5);
   U7 : INV_X1 port map( A => A, ZN => n6);
   U8 : INV_X1 port map( A => Ci, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_954 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_954;

architecture SYN_BEHAVIORAL of FA_954 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net166205, n4, n5 : std_logic;

begin
   
   U1 : OAI21_X1 port map( B1 => n4, B2 => n5, A => net166205, ZN => Co);
   U2 : INV_X1 port map( A => Ci, ZN => n4);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => net166205);
   U4 : XNOR2_X1 port map( A => Ci, B => n5, ZN => S);
   U5 : XNOR2_X1 port map( A => A, B => B, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_953 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_953;

architecture SYN_BEHAVIORAL of FA_953 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => n4);
   U2 : AOI21_X1 port map( B1 => Ci, B2 => n6, A => n4, ZN => n2);
   U3 : INV_X1 port map( A => n2, ZN => Co);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n6);
   U5 : XNOR2_X1 port map( A => Ci, B => n5, ZN => S);
   U6 : XNOR2_X1 port map( A => A, B => B, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_952 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_952;

architecture SYN_BEHAVIORAL of FA_952 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : AOI22_X1 port map( A1 => B, A2 => n5, B1 => Ci, B2 => n4, ZN => n2);
   U2 : CLKBUF_X1 port map( A => A, Z => n5);
   U5 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_951 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_951;

architecture SYN_BEHAVIORAL of FA_951 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => n4);
   U2 : AOI21_X1 port map( B1 => n5, B2 => Ci, A => n4, ZN => n2);
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U4 : INV_X1 port map( A => n6, ZN => n5);
   U5 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_950 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_950;

architecture SYN_BEHAVIORAL of FA_950 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : CLKBUF_X1 port map( A => A, Z => n4);
   U2 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => n4, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_949 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_949;

architecture SYN_BEHAVIORAL of FA_949 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n8);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n5, B1 => n6, B2 => n7, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U5 : INV_X1 port map( A => A, ZN => n5);
   U6 : INV_X1 port map( A => Ci, ZN => n6);
   U7 : INV_X1 port map( A => n8, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_948 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_948;

architecture SYN_BEHAVIORAL of FA_948 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => Ci, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_947 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_947;

architecture SYN_BEHAVIORAL of FA_947 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_946 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_946;

architecture SYN_BEHAVIORAL of FA_946 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_945 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_945;

architecture SYN_BEHAVIORAL of FA_945 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : CLKBUF_X1 port map( A => A, Z => n4);
   U2 : AOI22_X1 port map( A1 => B, A2 => n4, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_944 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_944;

architecture SYN_BEHAVIORAL of FA_944 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_943 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_943;

architecture SYN_BEHAVIORAL of FA_943 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_942 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_942;

architecture SYN_BEHAVIORAL of FA_942 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : CLKBUF_X1 port map( A => A, Z => n4);
   U2 : AOI22_X1 port map( A1 => B, A2 => n4, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_941 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_941;

architecture SYN_BEHAVIORAL of FA_941 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_940 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_940;

architecture SYN_BEHAVIORAL of FA_940 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_939 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_939;

architecture SYN_BEHAVIORAL of FA_939 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_938 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_938;

architecture SYN_BEHAVIORAL of FA_938 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n9);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : INV_X1 port map( A => B, ZN => n5);
   U5 : NAND2_X1 port map( A1 => n7, A2 => n8, ZN => Co);
   U6 : OR2_X1 port map( A1 => n4, A2 => n5, ZN => n7);
   U7 : NAND2_X1 port map( A1 => n9, A2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_937 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_937;

architecture SYN_BEHAVIORAL of FA_937 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_936 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_936;

architecture SYN_BEHAVIORAL of FA_936 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n6);
   U1 : CLKBUF_X1 port map( A => Ci, Z => n4);
   U2 : XNOR2_X1 port map( A => n4, B => n5, ZN => S);
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n5);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_935 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_935;

architecture SYN_BEHAVIORAL of FA_935 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_934 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_934;

architecture SYN_BEHAVIORAL of FA_934 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_933 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_933;

architecture SYN_BEHAVIORAL of FA_933 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_932 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_932;

architecture SYN_BEHAVIORAL of FA_932 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_931 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_931;

architecture SYN_BEHAVIORAL of FA_931 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_930 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_930;

architecture SYN_BEHAVIORAL of FA_930 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_929 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_929;

architecture SYN_BEHAVIORAL of FA_929 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_928 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_928;

architecture SYN_BEHAVIORAL of FA_928 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_927 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_927;

architecture SYN_BEHAVIORAL of FA_927 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_926 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_926;

architecture SYN_BEHAVIORAL of FA_926 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_925 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_925;

architecture SYN_BEHAVIORAL of FA_925 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_924 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_924;

architecture SYN_BEHAVIORAL of FA_924 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_923 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_923;

architecture SYN_BEHAVIORAL of FA_923 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_922 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_922;

architecture SYN_BEHAVIORAL of FA_922 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_921 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_921;

architecture SYN_BEHAVIORAL of FA_921 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_920 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_920;

architecture SYN_BEHAVIORAL of FA_920 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_919 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_919;

architecture SYN_BEHAVIORAL of FA_919 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_918 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_918;

architecture SYN_BEHAVIORAL of FA_918 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_917 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_917;

architecture SYN_BEHAVIORAL of FA_917 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_916 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_916;

architecture SYN_BEHAVIORAL of FA_916 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_915 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_915;

architecture SYN_BEHAVIORAL of FA_915 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_914 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_914;

architecture SYN_BEHAVIORAL of FA_914 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_913 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_913;

architecture SYN_BEHAVIORAL of FA_913 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_912 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_912;

architecture SYN_BEHAVIORAL of FA_912 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_911 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_911;

architecture SYN_BEHAVIORAL of FA_911 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_910 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_910;

architecture SYN_BEHAVIORAL of FA_910 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_909 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_909;

architecture SYN_BEHAVIORAL of FA_909 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_908 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_908;

architecture SYN_BEHAVIORAL of FA_908 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_907 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_907;

architecture SYN_BEHAVIORAL of FA_907 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_906 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_906;

architecture SYN_BEHAVIORAL of FA_906 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_905 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_905;

architecture SYN_BEHAVIORAL of FA_905 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_904 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_904;

architecture SYN_BEHAVIORAL of FA_904 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_903 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_903;

architecture SYN_BEHAVIORAL of FA_903 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_902 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_902;

architecture SYN_BEHAVIORAL of FA_902 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_901 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_901;

architecture SYN_BEHAVIORAL of FA_901 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_900 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_900;

architecture SYN_BEHAVIORAL of FA_900 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_899 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_899;

architecture SYN_BEHAVIORAL of FA_899 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_898 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_898;

architecture SYN_BEHAVIORAL of FA_898 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_897 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_897;

architecture SYN_BEHAVIORAL of FA_897 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_896 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_896;

architecture SYN_BEHAVIORAL of FA_896 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_895 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_895;

architecture SYN_BEHAVIORAL of FA_895 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_894 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_894;

architecture SYN_BEHAVIORAL of FA_894 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_893 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_893;

architecture SYN_BEHAVIORAL of FA_893 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_892 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_892;

architecture SYN_BEHAVIORAL of FA_892 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_891 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_891;

architecture SYN_BEHAVIORAL of FA_891 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal net160811, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => net160811, Z => S);
   U1 : OAI21_X1 port map( B1 => n5, B2 => n6, A => n7, ZN => Co);
   U2 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n7);
   U4 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U5 : INV_X1 port map( A => n8, ZN => net160811);
   U6 : CLKBUF_X1 port map( A => n6, Z => n8);
   U7 : INV_X1 port map( A => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_890 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_890;

architecture SYN_BEHAVIORAL of FA_890 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U2 : OR2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : OAI21_X1 port map( B1 => n7, B2 => Ci, A => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);
   U6 : AND2_X1 port map( A1 => A, A2 => B, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_889 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_889;

architecture SYN_BEHAVIORAL of FA_889 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U1 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => n4, B2 => Ci, ZN => n2);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_888 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_888;

architecture SYN_BEHAVIORAL of FA_888 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U1 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_887 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_887;

architecture SYN_BEHAVIORAL of FA_887 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U2 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_886 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_886;

architecture SYN_BEHAVIORAL of FA_886 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_885 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_885;

architecture SYN_BEHAVIORAL of FA_885 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U1 : XNOR2_X1 port map( A => B, B => n5, ZN => n8);
   U2 : OAI22_X1 port map( A1 => n4, A2 => n5, B1 => n6, B2 => n7, ZN => Co);
   U4 : INV_X1 port map( A => B, ZN => n4);
   U5 : INV_X1 port map( A => A, ZN => n5);
   U6 : INV_X1 port map( A => Ci, ZN => n6);
   U7 : INV_X1 port map( A => n8, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_884 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_884;

architecture SYN_BEHAVIORAL of FA_884 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => n6, B => B, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_883 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_883;

architecture SYN_BEHAVIORAL of FA_883 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_882 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_882;

architecture SYN_BEHAVIORAL of FA_882 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => n4);
   U2 : AOI21_X1 port map( B1 => n5, B2 => Ci, A => n4, ZN => n2);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U4 : INV_X1 port map( A => n6, ZN => n5);
   U5 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_881 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_881;

architecture SYN_BEHAVIORAL of FA_881 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => n6, B => B, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_880 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_880;

architecture SYN_BEHAVIORAL of FA_880 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U5 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_879 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_879;

architecture SYN_BEHAVIORAL of FA_879 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_878 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_878;

architecture SYN_BEHAVIORAL of FA_878 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_877 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_877;

architecture SYN_BEHAVIORAL of FA_877 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => n5, B => B, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_876 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_876;

architecture SYN_BEHAVIORAL of FA_876 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_875 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_875;

architecture SYN_BEHAVIORAL of FA_875 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_874 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_874;

architecture SYN_BEHAVIORAL of FA_874 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_873 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_873;

architecture SYN_BEHAVIORAL of FA_873 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_872 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_872;

architecture SYN_BEHAVIORAL of FA_872 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_871 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_871;

architecture SYN_BEHAVIORAL of FA_871 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_870 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_870;

architecture SYN_BEHAVIORAL of FA_870 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_869 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_869;

architecture SYN_BEHAVIORAL of FA_869 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_868 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_868;

architecture SYN_BEHAVIORAL of FA_868 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_867 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_867;

architecture SYN_BEHAVIORAL of FA_867 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_866 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_866;

architecture SYN_BEHAVIORAL of FA_866 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n4);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n8, ZN => n5);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => n7, B => B, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_865 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_865;

architecture SYN_BEHAVIORAL of FA_865 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_864 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_864;

architecture SYN_BEHAVIORAL of FA_864 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_863 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_863;

architecture SYN_BEHAVIORAL of FA_863 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_862 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_862;

architecture SYN_BEHAVIORAL of FA_862 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_861 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_861;

architecture SYN_BEHAVIORAL of FA_861 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_860 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_860;

architecture SYN_BEHAVIORAL of FA_860 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_859 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_859;

architecture SYN_BEHAVIORAL of FA_859 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_858 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_858;

architecture SYN_BEHAVIORAL of FA_858 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_857 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_857;

architecture SYN_BEHAVIORAL of FA_857 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_856 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_856;

architecture SYN_BEHAVIORAL of FA_856 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_855 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_855;

architecture SYN_BEHAVIORAL of FA_855 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => n5, B => B, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_854 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_854;

architecture SYN_BEHAVIORAL of FA_854 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_853 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_853;

architecture SYN_BEHAVIORAL of FA_853 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => n6, B2 => Ci, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_852 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_852;

architecture SYN_BEHAVIORAL of FA_852 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_851 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_851;

architecture SYN_BEHAVIORAL of FA_851 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_850 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_850;

architecture SYN_BEHAVIORAL of FA_850 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_849 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_849;

architecture SYN_BEHAVIORAL of FA_849 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_848 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_848;

architecture SYN_BEHAVIORAL of FA_848 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_847 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_847;

architecture SYN_BEHAVIORAL of FA_847 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_846 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_846;

architecture SYN_BEHAVIORAL of FA_846 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_845 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_845;

architecture SYN_BEHAVIORAL of FA_845 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_844 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_844;

architecture SYN_BEHAVIORAL of FA_844 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_843 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_843;

architecture SYN_BEHAVIORAL of FA_843 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_842 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_842;

architecture SYN_BEHAVIORAL of FA_842 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_841 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_841;

architecture SYN_BEHAVIORAL of FA_841 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_840 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_840;

architecture SYN_BEHAVIORAL of FA_840 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_839 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_839;

architecture SYN_BEHAVIORAL of FA_839 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_838 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_838;

architecture SYN_BEHAVIORAL of FA_838 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_837 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_837;

architecture SYN_BEHAVIORAL of FA_837 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_836 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_836;

architecture SYN_BEHAVIORAL of FA_836 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_835 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_835;

architecture SYN_BEHAVIORAL of FA_835 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X32
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : XNOR2_X1 port map( A => n4, B => B, ZN => n5);
   U2 : INV_X32 port map( A => A, ZN => n4);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_834 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_834;

architecture SYN_BEHAVIORAL of FA_834 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_833 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_833;

architecture SYN_BEHAVIORAL of FA_833 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : INV_X1 port map( A => A, ZN => n4);
   U4 : XNOR2_X1 port map( A => n4, B => B, ZN => n5);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_832 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_832;

architecture SYN_BEHAVIORAL of FA_832 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_831 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_831;

architecture SYN_BEHAVIORAL of FA_831 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_830 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_830;

architecture SYN_BEHAVIORAL of FA_830 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_829 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_829;

architecture SYN_BEHAVIORAL of FA_829 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_828 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_828;

architecture SYN_BEHAVIORAL of FA_828 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_827 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_827;

architecture SYN_BEHAVIORAL of FA_827 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_826 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_826;

architecture SYN_BEHAVIORAL of FA_826 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_825 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_825;

architecture SYN_BEHAVIORAL of FA_825 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => n7, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n8, ZN => Co);
   U7 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => n7, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_824 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_824;

architecture SYN_BEHAVIORAL of FA_824 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : CLKBUF_X1 port map( A => Ci, Z => n4);
   U4 : CLKBUF_X1 port map( A => n8, Z => n5);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n8);
   U6 : CLKBUF_X1 port map( A => B, Z => n7);
   U7 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n8, ZN => n9);
   U8 : INV_X1 port map( A => n9, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_823 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_823;

architecture SYN_BEHAVIORAL of FA_823 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : NAND2_X1 port map( A1 => n8, A2 => A, ZN => n4);
   U2 : NAND2_X1 port map( A1 => Ci, A2 => n7, ZN => n5);
   U4 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U5 : INV_X1 port map( A => A, ZN => n9);
   U6 : XNOR2_X1 port map( A => B, B => n9, ZN => n7);
   U7 : CLKBUF_X1 port map( A => B, Z => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_822 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_822;

architecture SYN_BEHAVIORAL of FA_822 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n5, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_821 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_821;

architecture SYN_BEHAVIORAL of FA_821 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : OAI22_X1 port map( A1 => n5, A2 => n9, B1 => n6, B2 => n7, ZN => Co);
   U4 : INV_X1 port map( A => n4, ZN => n5);
   U5 : INV_X1 port map( A => Ci, ZN => n6);
   U6 : INV_X1 port map( A => n8, ZN => n7);
   U7 : INV_X1 port map( A => A, ZN => n9);
   U8 : XNOR2_X1 port map( A => B, B => n9, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_820 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_820;

architecture SYN_BEHAVIORAL of FA_820 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => A, ZN => n6);
   U4 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n5, ZN => n2);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_819 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_819;

architecture SYN_BEHAVIORAL of FA_819 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n5);
   U5 : INV_X1 port map( A => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_818 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_818;

architecture SYN_BEHAVIORAL of FA_818 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => B, B => A, Z => n7);
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : NAND2_X1 port map( A1 => n8, A2 => A, ZN => n4);
   U2 : NAND2_X1 port map( A1 => Ci, A2 => n7, ZN => n5);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : CLKBUF_X1 port map( A => B, Z => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_817 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_817;

architecture SYN_BEHAVIORAL of FA_817 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_816 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_816;

architecture SYN_BEHAVIORAL of FA_816 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n2);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_815 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_815;

architecture SYN_BEHAVIORAL of FA_815 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_814 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_814;

architecture SYN_BEHAVIORAL of FA_814 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_813 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_813;

architecture SYN_BEHAVIORAL of FA_813 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_812 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_812;

architecture SYN_BEHAVIORAL of FA_812 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_811 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_811;

architecture SYN_BEHAVIORAL of FA_811 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_810 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_810;

architecture SYN_BEHAVIORAL of FA_810 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_809 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_809;

architecture SYN_BEHAVIORAL of FA_809 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_808 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_808;

architecture SYN_BEHAVIORAL of FA_808 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_807 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_807;

architecture SYN_BEHAVIORAL of FA_807 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_806 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_806;

architecture SYN_BEHAVIORAL of FA_806 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_805 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_805;

architecture SYN_BEHAVIORAL of FA_805 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_804 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_804;

architecture SYN_BEHAVIORAL of FA_804 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_803 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_803;

architecture SYN_BEHAVIORAL of FA_803 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_802 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_802;

architecture SYN_BEHAVIORAL of FA_802 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_801 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_801;

architecture SYN_BEHAVIORAL of FA_801 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_800 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_800;

architecture SYN_BEHAVIORAL of FA_800 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_799 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_799;

architecture SYN_BEHAVIORAL of FA_799 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_798 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_798;

architecture SYN_BEHAVIORAL of FA_798 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_797 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_797;

architecture SYN_BEHAVIORAL of FA_797 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n8);
   U1 : NAND2_X1 port map( A1 => n7, A2 => A, ZN => n4);
   U2 : NAND2_X1 port map( A1 => Ci, A2 => n8, ZN => n5);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : CLKBUF_X1 port map( A => B, Z => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_796 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_796;

architecture SYN_BEHAVIORAL of FA_796 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_795 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_795;

architecture SYN_BEHAVIORAL of FA_795 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_794 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_794;

architecture SYN_BEHAVIORAL of FA_794 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_793 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_793;

architecture SYN_BEHAVIORAL of FA_793 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_792 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_792;

architecture SYN_BEHAVIORAL of FA_792 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_791 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_791;

architecture SYN_BEHAVIORAL of FA_791 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_790 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_790;

architecture SYN_BEHAVIORAL of FA_790 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_789 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_789;

architecture SYN_BEHAVIORAL of FA_789 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_788 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_788;

architecture SYN_BEHAVIORAL of FA_788 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_787 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_787;

architecture SYN_BEHAVIORAL of FA_787 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_786 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_786;

architecture SYN_BEHAVIORAL of FA_786 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_785 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_785;

architecture SYN_BEHAVIORAL of FA_785 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_784 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_784;

architecture SYN_BEHAVIORAL of FA_784 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_783 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_783;

architecture SYN_BEHAVIORAL of FA_783 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_782 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_782;

architecture SYN_BEHAVIORAL of FA_782 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_781 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_781;

architecture SYN_BEHAVIORAL of FA_781 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_780 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_780;

architecture SYN_BEHAVIORAL of FA_780 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_779 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_779;

architecture SYN_BEHAVIORAL of FA_779 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_778 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_778;

architecture SYN_BEHAVIORAL of FA_778 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_777 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_777;

architecture SYN_BEHAVIORAL of FA_777 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_776 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_776;

architecture SYN_BEHAVIORAL of FA_776 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_775 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_775;

architecture SYN_BEHAVIORAL of FA_775 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_774 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_774;

architecture SYN_BEHAVIORAL of FA_774 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_773 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_773;

architecture SYN_BEHAVIORAL of FA_773 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_772 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_772;

architecture SYN_BEHAVIORAL of FA_772 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_771 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_771;

architecture SYN_BEHAVIORAL of FA_771 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_770 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_770;

architecture SYN_BEHAVIORAL of FA_770 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_769 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_769;

architecture SYN_BEHAVIORAL of FA_769 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n7);
   U4 : CLKBUF_X1 port map( A => Ci, Z => n5);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : CLKBUF_X1 port map( A => B, Z => n6);
   U7 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => n7, B2 => n5, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_768 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_768;

architecture SYN_BEHAVIORAL of FA_768 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_767 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_767;

architecture SYN_BEHAVIORAL of FA_767 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_766 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_766;

architecture SYN_BEHAVIORAL of FA_766 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_765 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_765;

architecture SYN_BEHAVIORAL of FA_765 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_764 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_764;

architecture SYN_BEHAVIORAL of FA_764 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_763 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_763;

architecture SYN_BEHAVIORAL of FA_763 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_762 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_762;

architecture SYN_BEHAVIORAL of FA_762 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_761 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_761;

architecture SYN_BEHAVIORAL of FA_761 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_760 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_760;

architecture SYN_BEHAVIORAL of FA_760 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_759 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_759;

architecture SYN_BEHAVIORAL of FA_759 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => n7, Z => n4);
   U4 : XNOR2_X1 port map( A => n5, B => B, ZN => n7);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => n7, B2 => Ci, ZN => n8);
   U7 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_758 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_758;

architecture SYN_BEHAVIORAL of FA_758 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n6, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n8);
   U4 : CLKBUF_X1 port map( A => n8, Z => n5);
   U5 : CLKBUF_X1 port map( A => Ci, Z => n6);
   U6 : CLKBUF_X1 port map( A => B, Z => n7);
   U7 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n8, ZN => n9);
   U8 : INV_X1 port map( A => n9, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_757 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_757;

architecture SYN_BEHAVIORAL of FA_757 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n7, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => n8, ZN => n5);
   U5 : INV_X1 port map( A => Ci, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n7);
   U7 : XNOR2_X1 port map( A => B, B => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_756 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_756;

architecture SYN_BEHAVIORAL of FA_756 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n8);
   U2 : NAND2_X1 port map( A1 => n9, A2 => A, ZN => n4);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n7, ZN => n5);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => B, B => n8, ZN => n7);
   U7 : CLKBUF_X1 port map( A => B, Z => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_755 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_755;

architecture SYN_BEHAVIORAL of FA_755 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n5, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => n5, B2 => Ci, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_754 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_754;

architecture SYN_BEHAVIORAL of FA_754 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : INV_X1 port map( A => n2, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_753 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_753;

architecture SYN_BEHAVIORAL of FA_753 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : XNOR2_X1 port map( A => B, B => n6, ZN => n4);
   U5 : CLKBUF_X1 port map( A => B, Z => n5);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_752 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_752;

architecture SYN_BEHAVIORAL of FA_752 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_751 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_751;

architecture SYN_BEHAVIORAL of FA_751 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_750 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_750;

architecture SYN_BEHAVIORAL of FA_750 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => n5, B => B, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_749 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_749;

architecture SYN_BEHAVIORAL of FA_749 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_748 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_748;

architecture SYN_BEHAVIORAL of FA_748 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_747 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_747;

architecture SYN_BEHAVIORAL of FA_747 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_746 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_746;

architecture SYN_BEHAVIORAL of FA_746 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_745 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_745;

architecture SYN_BEHAVIORAL of FA_745 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_744 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_744;

architecture SYN_BEHAVIORAL of FA_744 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_743 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_743;

architecture SYN_BEHAVIORAL of FA_743 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_742 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_742;

architecture SYN_BEHAVIORAL of FA_742 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_741 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_741;

architecture SYN_BEHAVIORAL of FA_741 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_740 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_740;

architecture SYN_BEHAVIORAL of FA_740 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_739 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_739;

architecture SYN_BEHAVIORAL of FA_739 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_738 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_738;

architecture SYN_BEHAVIORAL of FA_738 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_737 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_737;

architecture SYN_BEHAVIORAL of FA_737 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_736 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_736;

architecture SYN_BEHAVIORAL of FA_736 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_735 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_735;

architecture SYN_BEHAVIORAL of FA_735 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_734 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_734;

architecture SYN_BEHAVIORAL of FA_734 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_733 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_733;

architecture SYN_BEHAVIORAL of FA_733 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_732 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_732;

architecture SYN_BEHAVIORAL of FA_732 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_731 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_731;

architecture SYN_BEHAVIORAL of FA_731 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_730 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_730;

architecture SYN_BEHAVIORAL of FA_730 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_729 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_729;

architecture SYN_BEHAVIORAL of FA_729 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_728 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_728;

architecture SYN_BEHAVIORAL of FA_728 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_727 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_727;

architecture SYN_BEHAVIORAL of FA_727 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_726 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_726;

architecture SYN_BEHAVIORAL of FA_726 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_725 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_725;

architecture SYN_BEHAVIORAL of FA_725 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n7, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : INV_X1 port map( A => n8, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n7);
   U7 : XNOR2_X1 port map( A => n7, B => B, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_724 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_724;

architecture SYN_BEHAVIORAL of FA_724 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_723 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_723;

architecture SYN_BEHAVIORAL of FA_723 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_722 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_722;

architecture SYN_BEHAVIORAL of FA_722 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_721 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_721;

architecture SYN_BEHAVIORAL of FA_721 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_720 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_720;

architecture SYN_BEHAVIORAL of FA_720 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_719 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_719;

architecture SYN_BEHAVIORAL of FA_719 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_718 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_718;

architecture SYN_BEHAVIORAL of FA_718 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n5, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_717 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_717;

architecture SYN_BEHAVIORAL of FA_717 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_716 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_716;

architecture SYN_BEHAVIORAL of FA_716 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_715 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_715;

architecture SYN_BEHAVIORAL of FA_715 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_714 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_714;

architecture SYN_BEHAVIORAL of FA_714 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_713 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_713;

architecture SYN_BEHAVIORAL of FA_713 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_712 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_712;

architecture SYN_BEHAVIORAL of FA_712 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_711 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_711;

architecture SYN_BEHAVIORAL of FA_711 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_710 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_710;

architecture SYN_BEHAVIORAL of FA_710 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_709 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_709;

architecture SYN_BEHAVIORAL of FA_709 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_708 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_708;

architecture SYN_BEHAVIORAL of FA_708 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_707 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_707;

architecture SYN_BEHAVIORAL of FA_707 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n7, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => n8, ZN => n5);
   U5 : INV_X1 port map( A => Ci, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n7);
   U7 : XNOR2_X1 port map( A => n7, B => B, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_706 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_706;

architecture SYN_BEHAVIORAL of FA_706 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_705 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_705;

architecture SYN_BEHAVIORAL of FA_705 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_704 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_704;

architecture SYN_BEHAVIORAL of FA_704 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_703 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_703;

architecture SYN_BEHAVIORAL of FA_703 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_702 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_702;

architecture SYN_BEHAVIORAL of FA_702 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_701 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_701;

architecture SYN_BEHAVIORAL of FA_701 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_700 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_700;

architecture SYN_BEHAVIORAL of FA_700 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_699 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_699;

architecture SYN_BEHAVIORAL of FA_699 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_698 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_698;

architecture SYN_BEHAVIORAL of FA_698 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_697 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_697;

architecture SYN_BEHAVIORAL of FA_697 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_696 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_696;

architecture SYN_BEHAVIORAL of FA_696 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_695 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_695;

architecture SYN_BEHAVIORAL of FA_695 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_694 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_694;

architecture SYN_BEHAVIORAL of FA_694 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_693 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_693;

architecture SYN_BEHAVIORAL of FA_693 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n7, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => n9, ZN => n5);
   U5 : INV_X1 port map( A => Ci, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n7);
   U7 : XNOR2_X1 port map( A => B, B => n7, ZN => n9);
   U8 : CLKBUF_X1 port map( A => n9, Z => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_692 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_692;

architecture SYN_BEHAVIORAL of FA_692 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n9, n10 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n9, B => n7, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n8, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => n10, ZN => n5);
   U5 : INV_X1 port map( A => Ci, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n8);
   U7 : CLKBUF_X1 port map( A => n10, Z => n7);
   U8 : XNOR2_X1 port map( A => B, B => n8, ZN => n10);
   U9 : CLKBUF_X1 port map( A => Ci, Z => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_691 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_691;

architecture SYN_BEHAVIORAL of FA_691 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n6, B2 => Ci, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_690 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_690;

architecture SYN_BEHAVIORAL of FA_690 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U4 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_689 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_689;

architecture SYN_BEHAVIORAL of FA_689 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : XNOR2_X1 port map( A => B, B => n6, ZN => n4);
   U5 : CLKBUF_X1 port map( A => B, Z => n5);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_688 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_688;

architecture SYN_BEHAVIORAL of FA_688 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_687 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_687;

architecture SYN_BEHAVIORAL of FA_687 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_686 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_686;

architecture SYN_BEHAVIORAL of FA_686 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_685 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_685;

architecture SYN_BEHAVIORAL of FA_685 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_684 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_684;

architecture SYN_BEHAVIORAL of FA_684 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_683 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_683;

architecture SYN_BEHAVIORAL of FA_683 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_682 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_682;

architecture SYN_BEHAVIORAL of FA_682 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_681 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_681;

architecture SYN_BEHAVIORAL of FA_681 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_680 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_680;

architecture SYN_BEHAVIORAL of FA_680 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_679 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_679;

architecture SYN_BEHAVIORAL of FA_679 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_678 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_678;

architecture SYN_BEHAVIORAL of FA_678 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_677 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_677;

architecture SYN_BEHAVIORAL of FA_677 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_676 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_676;

architecture SYN_BEHAVIORAL of FA_676 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : CLKBUF_X1 port map( A => B, Z => n5);
   U4 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_675 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_675;

architecture SYN_BEHAVIORAL of FA_675 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_674 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_674;

architecture SYN_BEHAVIORAL of FA_674 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_673 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_673;

architecture SYN_BEHAVIORAL of FA_673 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_672 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_672;

architecture SYN_BEHAVIORAL of FA_672 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_671 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_671;

architecture SYN_BEHAVIORAL of FA_671 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_670 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_670;

architecture SYN_BEHAVIORAL of FA_670 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_669 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_669;

architecture SYN_BEHAVIORAL of FA_669 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_668 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_668;

architecture SYN_BEHAVIORAL of FA_668 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_667 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_667;

architecture SYN_BEHAVIORAL of FA_667 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_666 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_666;

architecture SYN_BEHAVIORAL of FA_666 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_665 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_665;

architecture SYN_BEHAVIORAL of FA_665 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_664 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_664;

architecture SYN_BEHAVIORAL of FA_664 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_663 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_663;

architecture SYN_BEHAVIORAL of FA_663 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_662 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_662;

architecture SYN_BEHAVIORAL of FA_662 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_661 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_661;

architecture SYN_BEHAVIORAL of FA_661 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : NAND2_X1 port map( A1 => n8, A2 => A, ZN => n4);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n9, ZN => n5);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n9);
   U7 : CLKBUF_X1 port map( A => B, Z => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_660 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_660;

architecture SYN_BEHAVIORAL of FA_660 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_659 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_659;

architecture SYN_BEHAVIORAL of FA_659 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : NAND2_X1 port map( A1 => n8, A2 => A, ZN => n4);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n9, ZN => n5);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => n7, B => B, ZN => n9);
   U7 : CLKBUF_X1 port map( A => B, Z => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_658 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_658;

architecture SYN_BEHAVIORAL of FA_658 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_657 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_657;

architecture SYN_BEHAVIORAL of FA_657 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n4);
   U2 : INV_X1 port map( A => n4, ZN => Co);
   U4 : INV_X1 port map( A => A, ZN => n5);
   U5 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_656 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_656;

architecture SYN_BEHAVIORAL of FA_656 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_655 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_655;

architecture SYN_BEHAVIORAL of FA_655 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_654 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_654;

architecture SYN_BEHAVIORAL of FA_654 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n6, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_653 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_653;

architecture SYN_BEHAVIORAL of FA_653 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_652 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_652;

architecture SYN_BEHAVIORAL of FA_652 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_651 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_651;

architecture SYN_BEHAVIORAL of FA_651 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_650 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_650;

architecture SYN_BEHAVIORAL of FA_650 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_649 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_649;

architecture SYN_BEHAVIORAL of FA_649 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_648 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_648;

architecture SYN_BEHAVIORAL of FA_648 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_647 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_647;

architecture SYN_BEHAVIORAL of FA_647 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_646 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_646;

architecture SYN_BEHAVIORAL of FA_646 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_645 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_645;

architecture SYN_BEHAVIORAL of FA_645 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_644 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_644;

architecture SYN_BEHAVIORAL of FA_644 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_643 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_643;

architecture SYN_BEHAVIORAL of FA_643 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_642 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_642;

architecture SYN_BEHAVIORAL of FA_642 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_641 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_641;

architecture SYN_BEHAVIORAL of FA_641 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => n7, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => Co);
   U6 : CLKBUF_X1 port map( A => B, Z => n6);
   U7 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => n4, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_640 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_640;

architecture SYN_BEHAVIORAL of FA_640 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_639 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_639;

architecture SYN_BEHAVIORAL of FA_639 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_638 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_638;

architecture SYN_BEHAVIORAL of FA_638 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_637 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_637;

architecture SYN_BEHAVIORAL of FA_637 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_636 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_636;

architecture SYN_BEHAVIORAL of FA_636 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_635 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_635;

architecture SYN_BEHAVIORAL of FA_635 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_634 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_634;

architecture SYN_BEHAVIORAL of FA_634 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_633 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_633;

architecture SYN_BEHAVIORAL of FA_633 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_632 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_632;

architecture SYN_BEHAVIORAL of FA_632 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_631 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_631;

architecture SYN_BEHAVIORAL of FA_631 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_630 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_630;

architecture SYN_BEHAVIORAL of FA_630 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_629 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_629;

architecture SYN_BEHAVIORAL of FA_629 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_628 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_628;

architecture SYN_BEHAVIORAL of FA_628 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_627 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_627;

architecture SYN_BEHAVIORAL of FA_627 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n6, B2 => Ci, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => n6, Z => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_626 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_626;

architecture SYN_BEHAVIORAL of FA_626 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_625 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_625;

architecture SYN_BEHAVIORAL of FA_625 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : XNOR2_X1 port map( A => B, B => n6, ZN => n4);
   U4 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U5 : CLKBUF_X1 port map( A => B, Z => n5);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_624 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_624;

architecture SYN_BEHAVIORAL of FA_624 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : INV_X1 port map( A => n2, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_623 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_623;

architecture SYN_BEHAVIORAL of FA_623 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : XNOR2_X1 port map( A => B, B => n8, ZN => n4);
   U2 : XNOR2_X1 port map( A => n6, B => n8, ZN => n5);
   U4 : OAI22_X1 port map( A1 => n6, A2 => n8, B1 => n7, B2 => n5, ZN => Co);
   U5 : INV_X1 port map( A => B, ZN => n6);
   U6 : INV_X1 port map( A => Ci, ZN => n7);
   U7 : INV_X1 port map( A => A, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_622 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_622;

architecture SYN_BEHAVIORAL of FA_622 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => n4, B2 => Ci, ZN => n2);
   U4 : INV_X1 port map( A => n2, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_621 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_621;

architecture SYN_BEHAVIORAL of FA_621 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_620 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_620;

architecture SYN_BEHAVIORAL of FA_620 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_619 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_619;

architecture SYN_BEHAVIORAL of FA_619 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_618 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_618;

architecture SYN_BEHAVIORAL of FA_618 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_617 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_617;

architecture SYN_BEHAVIORAL of FA_617 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_616 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_616;

architecture SYN_BEHAVIORAL of FA_616 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_615 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_615;

architecture SYN_BEHAVIORAL of FA_615 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_614 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_614;

architecture SYN_BEHAVIORAL of FA_614 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_613 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_613;

architecture SYN_BEHAVIORAL of FA_613 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_612 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_612;

architecture SYN_BEHAVIORAL of FA_612 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_611 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_611;

architecture SYN_BEHAVIORAL of FA_611 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_610 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_610;

architecture SYN_BEHAVIORAL of FA_610 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_609 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_609;

architecture SYN_BEHAVIORAL of FA_609 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_608 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_608;

architecture SYN_BEHAVIORAL of FA_608 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_607 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_607;

architecture SYN_BEHAVIORAL of FA_607 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_606 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_606;

architecture SYN_BEHAVIORAL of FA_606 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_605 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_605;

architecture SYN_BEHAVIORAL of FA_605 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_604 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_604;

architecture SYN_BEHAVIORAL of FA_604 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_603 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_603;

architecture SYN_BEHAVIORAL of FA_603 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_602 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_602;

architecture SYN_BEHAVIORAL of FA_602 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_601 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_601;

architecture SYN_BEHAVIORAL of FA_601 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_600 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_600;

architecture SYN_BEHAVIORAL of FA_600 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_599 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_599;

architecture SYN_BEHAVIORAL of FA_599 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_598 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_598;

architecture SYN_BEHAVIORAL of FA_598 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => n5, B2 => Ci, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_597 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_597;

architecture SYN_BEHAVIORAL of FA_597 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n8);
   U2 : NAND2_X1 port map( A1 => n9, A2 => A, ZN => n4);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n7, ZN => n5);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : CLKBUF_X1 port map( A => B, Z => n9);
   U7 : XNOR2_X1 port map( A => B, B => n8, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_596 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_596;

architecture SYN_BEHAVIORAL of FA_596 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_595 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_595;

architecture SYN_BEHAVIORAL of FA_595 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_594 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_594;

architecture SYN_BEHAVIORAL of FA_594 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n9);
   U2 : NAND2_X1 port map( A1 => n8, A2 => A, ZN => n4);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n7, ZN => n5);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : CLKBUF_X1 port map( A => B, Z => n8);
   U7 : XNOR2_X1 port map( A => B, B => n9, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_593 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_593;

architecture SYN_BEHAVIORAL of FA_593 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => n7, B => B, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_592 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_592;

architecture SYN_BEHAVIORAL of FA_592 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_591 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_591;

architecture SYN_BEHAVIORAL of FA_591 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_590 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_590;

architecture SYN_BEHAVIORAL of FA_590 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_589 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_589;

architecture SYN_BEHAVIORAL of FA_589 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => n7, B => B, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_588 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_588;

architecture SYN_BEHAVIORAL of FA_588 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_587 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_587;

architecture SYN_BEHAVIORAL of FA_587 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_586 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_586;

architecture SYN_BEHAVIORAL of FA_586 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_585 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_585;

architecture SYN_BEHAVIORAL of FA_585 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_584 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_584;

architecture SYN_BEHAVIORAL of FA_584 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => n7, B => B, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_583 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_583;

architecture SYN_BEHAVIORAL of FA_583 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_582 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_582;

architecture SYN_BEHAVIORAL of FA_582 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n8, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : INV_X1 port map( A => n7, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n8);
   U7 : XNOR2_X1 port map( A => B, B => n8, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_581 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_581;

architecture SYN_BEHAVIORAL of FA_581 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_580 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_580;

architecture SYN_BEHAVIORAL of FA_580 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_579 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_579;

architecture SYN_BEHAVIORAL of FA_579 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_578 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_578;

architecture SYN_BEHAVIORAL of FA_578 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => n4, B2 => Ci, ZN => n2);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_577 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_577;

architecture SYN_BEHAVIORAL of FA_577 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => n7, Z => n5);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n8, ZN => Co);
   U7 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => n5, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_576 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_576;

architecture SYN_BEHAVIORAL of FA_576 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_575 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_575;

architecture SYN_BEHAVIORAL of FA_575 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_574 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_574;

architecture SYN_BEHAVIORAL of FA_574 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_573 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_573;

architecture SYN_BEHAVIORAL of FA_573 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_572 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_572;

architecture SYN_BEHAVIORAL of FA_572 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_571 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_571;

architecture SYN_BEHAVIORAL of FA_571 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_570 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_570;

architecture SYN_BEHAVIORAL of FA_570 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_569 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_569;

architecture SYN_BEHAVIORAL of FA_569 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_568 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_568;

architecture SYN_BEHAVIORAL of FA_568 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_567 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_567;

architecture SYN_BEHAVIORAL of FA_567 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_566 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_566;

architecture SYN_BEHAVIORAL of FA_566 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_565 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_565;

architecture SYN_BEHAVIORAL of FA_565 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_564 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_564;

architecture SYN_BEHAVIORAL of FA_564 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_563 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_563;

architecture SYN_BEHAVIORAL of FA_563 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_562 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_562;

architecture SYN_BEHAVIORAL of FA_562 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_561 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_561;

architecture SYN_BEHAVIORAL of FA_561 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n6, B2 => Ci, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_560 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_560;

architecture SYN_BEHAVIORAL of FA_560 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => n6, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_559 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_559;

architecture SYN_BEHAVIORAL of FA_559 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n7, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => n8, ZN => n5);
   U5 : INV_X1 port map( A => Ci, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n7);
   U7 : XNOR2_X1 port map( A => B, B => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_558 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_558;

architecture SYN_BEHAVIORAL of FA_558 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U4 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_557 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_557;

architecture SYN_BEHAVIORAL of FA_557 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : INV_X1 port map( A => n2, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_556 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_556;

architecture SYN_BEHAVIORAL of FA_556 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_555 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_555;

architecture SYN_BEHAVIORAL of FA_555 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : INV_X1 port map( A => n2, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n5);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_554 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_554;

architecture SYN_BEHAVIORAL of FA_554 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_553 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_553;

architecture SYN_BEHAVIORAL of FA_553 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_552 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_552;

architecture SYN_BEHAVIORAL of FA_552 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_551 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_551;

architecture SYN_BEHAVIORAL of FA_551 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_550 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_550;

architecture SYN_BEHAVIORAL of FA_550 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_549 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_549;

architecture SYN_BEHAVIORAL of FA_549 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_548 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_548;

architecture SYN_BEHAVIORAL of FA_548 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_547 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_547;

architecture SYN_BEHAVIORAL of FA_547 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_546 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_546;

architecture SYN_BEHAVIORAL of FA_546 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_545 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_545;

architecture SYN_BEHAVIORAL of FA_545 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_544 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_544;

architecture SYN_BEHAVIORAL of FA_544 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_543 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_543;

architecture SYN_BEHAVIORAL of FA_543 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_542 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_542;

architecture SYN_BEHAVIORAL of FA_542 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_541 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_541;

architecture SYN_BEHAVIORAL of FA_541 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_540 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_540;

architecture SYN_BEHAVIORAL of FA_540 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_539 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_539;

architecture SYN_BEHAVIORAL of FA_539 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_538 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_538;

architecture SYN_BEHAVIORAL of FA_538 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_537 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_537;

architecture SYN_BEHAVIORAL of FA_537 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_536 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_536;

architecture SYN_BEHAVIORAL of FA_536 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_535 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_535;

architecture SYN_BEHAVIORAL of FA_535 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_534 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_534;

architecture SYN_BEHAVIORAL of FA_534 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_533 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_533;

architecture SYN_BEHAVIORAL of FA_533 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_532 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_532;

architecture SYN_BEHAVIORAL of FA_532 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_531 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_531;

architecture SYN_BEHAVIORAL of FA_531 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_530 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_530;

architecture SYN_BEHAVIORAL of FA_530 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_529 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_529;

architecture SYN_BEHAVIORAL of FA_529 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_528 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_528;

architecture SYN_BEHAVIORAL of FA_528 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_527 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_527;

architecture SYN_BEHAVIORAL of FA_527 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_526 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_526;

architecture SYN_BEHAVIORAL of FA_526 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_525 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_525;

architecture SYN_BEHAVIORAL of FA_525 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_524 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_524;

architecture SYN_BEHAVIORAL of FA_524 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_523 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_523;

architecture SYN_BEHAVIORAL of FA_523 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_522 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_522;

architecture SYN_BEHAVIORAL of FA_522 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_521 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_521;

architecture SYN_BEHAVIORAL of FA_521 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_520 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_520;

architecture SYN_BEHAVIORAL of FA_520 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : NAND2_X1 port map( A1 => n8, A2 => A, ZN => n4);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n9, ZN => n5);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n9);
   U7 : CLKBUF_X1 port map( A => B, Z => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_519 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_519;

architecture SYN_BEHAVIORAL of FA_519 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_518 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_518;

architecture SYN_BEHAVIORAL of FA_518 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_517 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_517;

architecture SYN_BEHAVIORAL of FA_517 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => n5, B => B, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_516 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_516;

architecture SYN_BEHAVIORAL of FA_516 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_515 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_515;

architecture SYN_BEHAVIORAL of FA_515 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_514 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_514;

architecture SYN_BEHAVIORAL of FA_514 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => n4, B2 => Ci, ZN => n2);
   U4 : XNOR2_X1 port map( A => B, B => n6, ZN => n4);
   U5 : CLKBUF_X1 port map( A => B, Z => n5);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_513 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_513;

architecture SYN_BEHAVIORAL of FA_513 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : CLKBUF_X1 port map( A => n7, Z => n4);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n7);
   U6 : INV_X1 port map( A => n8, ZN => Co);
   U7 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => n4, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_512 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_512;

architecture SYN_BEHAVIORAL of FA_512 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_511 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_511;

architecture SYN_BEHAVIORAL of FA_511 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_510 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_510;

architecture SYN_BEHAVIORAL of FA_510 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_509 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_509;

architecture SYN_BEHAVIORAL of FA_509 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_508 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_508;

architecture SYN_BEHAVIORAL of FA_508 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_507 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_507;

architecture SYN_BEHAVIORAL of FA_507 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_506 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_506;

architecture SYN_BEHAVIORAL of FA_506 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_505 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_505;

architecture SYN_BEHAVIORAL of FA_505 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_504 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_504;

architecture SYN_BEHAVIORAL of FA_504 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_503 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_503;

architecture SYN_BEHAVIORAL of FA_503 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_502 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_502;

architecture SYN_BEHAVIORAL of FA_502 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_501 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_501;

architecture SYN_BEHAVIORAL of FA_501 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_500 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_500;

architecture SYN_BEHAVIORAL of FA_500 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_499 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_499;

architecture SYN_BEHAVIORAL of FA_499 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_498 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_498;

architecture SYN_BEHAVIORAL of FA_498 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_497 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_497;

architecture SYN_BEHAVIORAL of FA_497 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_496 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_496;

architecture SYN_BEHAVIORAL of FA_496 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_495 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_495;

architecture SYN_BEHAVIORAL of FA_495 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n7, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => n8, ZN => n5);
   U5 : INV_X1 port map( A => Ci, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n7);
   U7 : XNOR2_X1 port map( A => B, B => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_494 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_494;

architecture SYN_BEHAVIORAL of FA_494 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n6, B2 => Ci, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_493 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_493;

architecture SYN_BEHAVIORAL of FA_493 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U4 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_492 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_492;

architecture SYN_BEHAVIORAL of FA_492 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_491 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_491;

architecture SYN_BEHAVIORAL of FA_491 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : INV_X1 port map( A => n2, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n5);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_490 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_490;

architecture SYN_BEHAVIORAL of FA_490 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_489 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_489;

architecture SYN_BEHAVIORAL of FA_489 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_488 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_488;

architecture SYN_BEHAVIORAL of FA_488 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_487 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_487;

architecture SYN_BEHAVIORAL of FA_487 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_486 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_486;

architecture SYN_BEHAVIORAL of FA_486 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_485 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_485;

architecture SYN_BEHAVIORAL of FA_485 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_484 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_484;

architecture SYN_BEHAVIORAL of FA_484 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_483 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_483;

architecture SYN_BEHAVIORAL of FA_483 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_482 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_482;

architecture SYN_BEHAVIORAL of FA_482 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_481 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_481;

architecture SYN_BEHAVIORAL of FA_481 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_480 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_480;

architecture SYN_BEHAVIORAL of FA_480 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_479 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_479;

architecture SYN_BEHAVIORAL of FA_479 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_478 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_478;

architecture SYN_BEHAVIORAL of FA_478 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_477 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_477;

architecture SYN_BEHAVIORAL of FA_477 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_476 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_476;

architecture SYN_BEHAVIORAL of FA_476 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_475 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_475;

architecture SYN_BEHAVIORAL of FA_475 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_474 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_474;

architecture SYN_BEHAVIORAL of FA_474 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_473 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_473;

architecture SYN_BEHAVIORAL of FA_473 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_472 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_472;

architecture SYN_BEHAVIORAL of FA_472 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_471 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_471;

architecture SYN_BEHAVIORAL of FA_471 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n6, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_470 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_470;

architecture SYN_BEHAVIORAL of FA_470 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => n6, B2 => Ci, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_469 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_469;

architecture SYN_BEHAVIORAL of FA_469 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_468 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_468;

architecture SYN_BEHAVIORAL of FA_468 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_467 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_467;

architecture SYN_BEHAVIORAL of FA_467 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_466 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_466;

architecture SYN_BEHAVIORAL of FA_466 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_465 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_465;

architecture SYN_BEHAVIORAL of FA_465 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_464 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_464;

architecture SYN_BEHAVIORAL of FA_464 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_463 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_463;

architecture SYN_BEHAVIORAL of FA_463 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_462 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_462;

architecture SYN_BEHAVIORAL of FA_462 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n7, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : INV_X1 port map( A => n8, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n7);
   U7 : XNOR2_X1 port map( A => B, B => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_461 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_461;

architecture SYN_BEHAVIORAL of FA_461 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_460 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_460;

architecture SYN_BEHAVIORAL of FA_460 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_459 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_459;

architecture SYN_BEHAVIORAL of FA_459 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_458 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_458;

architecture SYN_BEHAVIORAL of FA_458 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_457 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_457;

architecture SYN_BEHAVIORAL of FA_457 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n6, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_456 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_456;

architecture SYN_BEHAVIORAL of FA_456 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n9, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : NAND2_X1 port map( A1 => n8, A2 => A, ZN => n4);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n9, ZN => n5);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n9);
   U7 : CLKBUF_X1 port map( A => B, Z => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_455 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_455;

architecture SYN_BEHAVIORAL of FA_455 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => n5, B => B, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_454 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_454;

architecture SYN_BEHAVIORAL of FA_454 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n4);
   U2 : INV_X1 port map( A => n4, ZN => Co);
   U4 : INV_X1 port map( A => A, ZN => n5);
   U5 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_453 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_453;

architecture SYN_BEHAVIORAL of FA_453 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_452 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_452;

architecture SYN_BEHAVIORAL of FA_452 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n6, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_451 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_451;

architecture SYN_BEHAVIORAL of FA_451 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n6, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_450 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_450;

architecture SYN_BEHAVIORAL of FA_450 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : XNOR2_X1 port map( A => B, B => n6, ZN => n4);
   U5 : CLKBUF_X1 port map( A => B, Z => n5);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_449 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_449;

architecture SYN_BEHAVIORAL of FA_449 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n8, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : CLKBUF_X1 port map( A => n8, Z => n4);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : CLKBUF_X1 port map( A => Ci, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n8);
   U7 : INV_X1 port map( A => n9, ZN => Co);
   U8 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => n4, B2 => n6, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_448 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_448;

architecture SYN_BEHAVIORAL of FA_448 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_447 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_447;

architecture SYN_BEHAVIORAL of FA_447 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_446 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_446;

architecture SYN_BEHAVIORAL of FA_446 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_445 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_445;

architecture SYN_BEHAVIORAL of FA_445 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_444 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_444;

architecture SYN_BEHAVIORAL of FA_444 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_443 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_443;

architecture SYN_BEHAVIORAL of FA_443 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_442 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_442;

architecture SYN_BEHAVIORAL of FA_442 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_441 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_441;

architecture SYN_BEHAVIORAL of FA_441 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_440 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_440;

architecture SYN_BEHAVIORAL of FA_440 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_439 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_439;

architecture SYN_BEHAVIORAL of FA_439 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_438 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_438;

architecture SYN_BEHAVIORAL of FA_438 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_437 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_437;

architecture SYN_BEHAVIORAL of FA_437 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_436 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_436;

architecture SYN_BEHAVIORAL of FA_436 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_435 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_435;

architecture SYN_BEHAVIORAL of FA_435 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_434 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_434;

architecture SYN_BEHAVIORAL of FA_434 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_433 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_433;

architecture SYN_BEHAVIORAL of FA_433 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_432 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_432;

architecture SYN_BEHAVIORAL of FA_432 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_431 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_431;

architecture SYN_BEHAVIORAL of FA_431 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_430 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_430;

architecture SYN_BEHAVIORAL of FA_430 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_429 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_429;

architecture SYN_BEHAVIORAL of FA_429 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : CLKBUF_X1 port map( A => n7, Z => n5);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n7);
   U6 : INV_X1 port map( A => n8, ZN => Co);
   U7 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n7, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_428 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_428;

architecture SYN_BEHAVIORAL of FA_428 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n7, B2 => Ci, ZN => n4);
   U2 : INV_X1 port map( A => n4, ZN => Co);
   U4 : INV_X1 port map( A => A, ZN => n6);
   U5 : CLKBUF_X1 port map( A => n7, Z => n5);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_427 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_427;

architecture SYN_BEHAVIORAL of FA_427 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : XNOR2_X1 port map( A => B, B => n6, ZN => n4);
   U4 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U5 : CLKBUF_X1 port map( A => B, Z => n5);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_426 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_426;

architecture SYN_BEHAVIORAL of FA_426 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n5, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_425 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_425;

architecture SYN_BEHAVIORAL of FA_425 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : XNOR2_X1 port map( A => B, B => n6, ZN => n4);
   U5 : CLKBUF_X1 port map( A => B, Z => n5);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_424 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_424;

architecture SYN_BEHAVIORAL of FA_424 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_423 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_423;

architecture SYN_BEHAVIORAL of FA_423 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_422 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_422;

architecture SYN_BEHAVIORAL of FA_422 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_421 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_421;

architecture SYN_BEHAVIORAL of FA_421 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_420 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_420;

architecture SYN_BEHAVIORAL of FA_420 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : XNOR2_X1 port map( A => B, B => n6, ZN => n4);
   U5 : CLKBUF_X1 port map( A => B, Z => n5);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_419 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_419;

architecture SYN_BEHAVIORAL of FA_419 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_418 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_418;

architecture SYN_BEHAVIORAL of FA_418 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_417 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_417;

architecture SYN_BEHAVIORAL of FA_417 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_416 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_416;

architecture SYN_BEHAVIORAL of FA_416 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_415 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_415;

architecture SYN_BEHAVIORAL of FA_415 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_414 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_414;

architecture SYN_BEHAVIORAL of FA_414 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_413 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_413;

architecture SYN_BEHAVIORAL of FA_413 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_412 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_412;

architecture SYN_BEHAVIORAL of FA_412 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_411 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_411;

architecture SYN_BEHAVIORAL of FA_411 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_410 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_410;

architecture SYN_BEHAVIORAL of FA_410 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_409 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_409;

architecture SYN_BEHAVIORAL of FA_409 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_408 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_408;

architecture SYN_BEHAVIORAL of FA_408 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_407 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_407;

architecture SYN_BEHAVIORAL of FA_407 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n6, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n6, B2 => Ci, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_406 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_406;

architecture SYN_BEHAVIORAL of FA_406 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_405 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_405;

architecture SYN_BEHAVIORAL of FA_405 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n6, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_404 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_404;

architecture SYN_BEHAVIORAL of FA_404 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_403 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_403;

architecture SYN_BEHAVIORAL of FA_403 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_402 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_402;

architecture SYN_BEHAVIORAL of FA_402 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_401 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_401;

architecture SYN_BEHAVIORAL of FA_401 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_400 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_400;

architecture SYN_BEHAVIORAL of FA_400 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_399 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_399;

architecture SYN_BEHAVIORAL of FA_399 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_398 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_398;

architecture SYN_BEHAVIORAL of FA_398 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_397 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_397;

architecture SYN_BEHAVIORAL of FA_397 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n6, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_396 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_396;

architecture SYN_BEHAVIORAL of FA_396 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_395 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_395;

architecture SYN_BEHAVIORAL of FA_395 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_394 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_394;

architecture SYN_BEHAVIORAL of FA_394 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_393 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_393;

architecture SYN_BEHAVIORAL of FA_393 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : OAI22_X1 port map( A1 => n5, A2 => n8, B1 => n6, B2 => n7, ZN => Co);
   U4 : INV_X1 port map( A => n4, ZN => n5);
   U5 : INV_X1 port map( A => Ci, ZN => n6);
   U6 : INV_X1 port map( A => n9, ZN => n7);
   U7 : INV_X1 port map( A => A, ZN => n8);
   U8 : XNOR2_X1 port map( A => B, B => n8, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_392 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_392;

architecture SYN_BEHAVIORAL of FA_392 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n6, B2 => Ci, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_391 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_391;

architecture SYN_BEHAVIORAL of FA_391 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_390 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_390;

architecture SYN_BEHAVIORAL of FA_390 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_389 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_389;

architecture SYN_BEHAVIORAL of FA_389 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n8);
   U2 : NAND2_X1 port map( A1 => n7, A2 => A, ZN => n4);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n9, ZN => n5);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : CLKBUF_X1 port map( A => B, Z => n7);
   U7 : XNOR2_X1 port map( A => B, B => n8, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_388 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_388;

architecture SYN_BEHAVIORAL of FA_388 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n6, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_387 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_387;

architecture SYN_BEHAVIORAL of FA_387 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n6, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_386 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_386;

architecture SYN_BEHAVIORAL of FA_386 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U4 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => n4, B2 => Ci, ZN => n2);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_385 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_385;

architecture SYN_BEHAVIORAL of FA_385 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => n7, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n8, ZN => Co);
   U7 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => n4, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_384 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_384;

architecture SYN_BEHAVIORAL of FA_384 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_383 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_383;

architecture SYN_BEHAVIORAL of FA_383 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_382 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_382;

architecture SYN_BEHAVIORAL of FA_382 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_381 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_381;

architecture SYN_BEHAVIORAL of FA_381 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_380 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_380;

architecture SYN_BEHAVIORAL of FA_380 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_379 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_379;

architecture SYN_BEHAVIORAL of FA_379 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_378 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_378;

architecture SYN_BEHAVIORAL of FA_378 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_377 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_377;

architecture SYN_BEHAVIORAL of FA_377 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_376 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_376;

architecture SYN_BEHAVIORAL of FA_376 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_375 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_375;

architecture SYN_BEHAVIORAL of FA_375 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_374 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_374;

architecture SYN_BEHAVIORAL of FA_374 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_373 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_373;

architecture SYN_BEHAVIORAL of FA_373 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_372 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_372;

architecture SYN_BEHAVIORAL of FA_372 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_371 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_371;

architecture SYN_BEHAVIORAL of FA_371 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_370 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_370;

architecture SYN_BEHAVIORAL of FA_370 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_369 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_369;

architecture SYN_BEHAVIORAL of FA_369 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_368 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_368;

architecture SYN_BEHAVIORAL of FA_368 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_367 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_367;

architecture SYN_BEHAVIORAL of FA_367 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_366 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_366;

architecture SYN_BEHAVIORAL of FA_366 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_365 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_365;

architecture SYN_BEHAVIORAL of FA_365 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_364 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_364;

architecture SYN_BEHAVIORAL of FA_364 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_363 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_363;

architecture SYN_BEHAVIORAL of FA_363 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => n6, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n6, B2 => Ci, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_362 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_362;

architecture SYN_BEHAVIORAL of FA_362 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : CLKBUF_X1 port map( A => Ci, Z => n4);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n7);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => n7, B2 => Ci, ZN => n8);
   U7 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_361 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_361;

architecture SYN_BEHAVIORAL of FA_361 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : XNOR2_X1 port map( A => B, B => n6, ZN => n4);
   U4 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U5 : CLKBUF_X1 port map( A => B, Z => n5);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_360 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_360;

architecture SYN_BEHAVIORAL of FA_360 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_359 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_359;

architecture SYN_BEHAVIORAL of FA_359 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_358 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_358;

architecture SYN_BEHAVIORAL of FA_358 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_357 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_357;

architecture SYN_BEHAVIORAL of FA_357 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_356 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_356;

architecture SYN_BEHAVIORAL of FA_356 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : XNOR2_X1 port map( A => B, B => n6, ZN => n4);
   U5 : CLKBUF_X1 port map( A => B, Z => n5);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_355 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_355;

architecture SYN_BEHAVIORAL of FA_355 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_354 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_354;

architecture SYN_BEHAVIORAL of FA_354 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_353 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_353;

architecture SYN_BEHAVIORAL of FA_353 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => n6, B2 => Ci, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_352 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_352;

architecture SYN_BEHAVIORAL of FA_352 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_351 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_351;

architecture SYN_BEHAVIORAL of FA_351 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_350 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_350;

architecture SYN_BEHAVIORAL of FA_350 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_349 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_349;

architecture SYN_BEHAVIORAL of FA_349 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_348 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_348;

architecture SYN_BEHAVIORAL of FA_348 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_347 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_347;

architecture SYN_BEHAVIORAL of FA_347 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_346 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_346;

architecture SYN_BEHAVIORAL of FA_346 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_345 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_345;

architecture SYN_BEHAVIORAL of FA_345 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_344 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_344;

architecture SYN_BEHAVIORAL of FA_344 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_343 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_343;

architecture SYN_BEHAVIORAL of FA_343 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_342 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_342;

architecture SYN_BEHAVIORAL of FA_342 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_341 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_341;

architecture SYN_BEHAVIORAL of FA_341 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_340 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_340;

architecture SYN_BEHAVIORAL of FA_340 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n6, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_339 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_339;

architecture SYN_BEHAVIORAL of FA_339 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_338 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_338;

architecture SYN_BEHAVIORAL of FA_338 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_337 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_337;

architecture SYN_BEHAVIORAL of FA_337 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_336 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_336;

architecture SYN_BEHAVIORAL of FA_336 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n7, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : INV_X1 port map( A => n8, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n7);
   U7 : XNOR2_X1 port map( A => B, B => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_335 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_335;

architecture SYN_BEHAVIORAL of FA_335 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_334 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_334;

architecture SYN_BEHAVIORAL of FA_334 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_333 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_333;

architecture SYN_BEHAVIORAL of FA_333 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_332 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_332;

architecture SYN_BEHAVIORAL of FA_332 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_331 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_331;

architecture SYN_BEHAVIORAL of FA_331 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_330 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_330;

architecture SYN_BEHAVIORAL of FA_330 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => n5, B => B, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_329 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_329;

architecture SYN_BEHAVIORAL of FA_329 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_328 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_328;

architecture SYN_BEHAVIORAL of FA_328 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_327 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_327;

architecture SYN_BEHAVIORAL of FA_327 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_326 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_326;

architecture SYN_BEHAVIORAL of FA_326 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : NAND2_X1 port map( A1 => n8, A2 => A, ZN => n4);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n9, ZN => n5);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n9);
   U7 : CLKBUF_X1 port map( A => B, Z => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_325 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_325;

architecture SYN_BEHAVIORAL of FA_325 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n6, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => n6, B2 => Ci, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_324 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_324;

architecture SYN_BEHAVIORAL of FA_324 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => n6, B2 => Ci, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_323 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_323;

architecture SYN_BEHAVIORAL of FA_323 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n6, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_322 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_322;

architecture SYN_BEHAVIORAL of FA_322 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U4 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => n4, B2 => Ci, ZN => n2);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_321 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_321;

architecture SYN_BEHAVIORAL of FA_321 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : CLKBUF_X1 port map( A => Ci, Z => n4);
   U4 : CLKBUF_X1 port map( A => n8, Z => n5);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n8);
   U7 : INV_X1 port map( A => n9, ZN => Co);
   U8 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => n5, B2 => n4, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_320 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_320;

architecture SYN_BEHAVIORAL of FA_320 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_319 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_319;

architecture SYN_BEHAVIORAL of FA_319 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_318 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_318;

architecture SYN_BEHAVIORAL of FA_318 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_317 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_317;

architecture SYN_BEHAVIORAL of FA_317 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_316 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_316;

architecture SYN_BEHAVIORAL of FA_316 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_315 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_315;

architecture SYN_BEHAVIORAL of FA_315 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_314 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_314;

architecture SYN_BEHAVIORAL of FA_314 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_313 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_313;

architecture SYN_BEHAVIORAL of FA_313 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_312 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_312;

architecture SYN_BEHAVIORAL of FA_312 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_311 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_311;

architecture SYN_BEHAVIORAL of FA_311 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_310 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_310;

architecture SYN_BEHAVIORAL of FA_310 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_309 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_309;

architecture SYN_BEHAVIORAL of FA_309 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_308 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_308;

architecture SYN_BEHAVIORAL of FA_308 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_307 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_307;

architecture SYN_BEHAVIORAL of FA_307 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_306 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_306;

architecture SYN_BEHAVIORAL of FA_306 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_305 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_305;

architecture SYN_BEHAVIORAL of FA_305 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_304 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_304;

architecture SYN_BEHAVIORAL of FA_304 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_303 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_303;

architecture SYN_BEHAVIORAL of FA_303 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_302 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_302;

architecture SYN_BEHAVIORAL of FA_302 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_301 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_301;

architecture SYN_BEHAVIORAL of FA_301 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_300 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_300;

architecture SYN_BEHAVIORAL of FA_300 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_299 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_299;

architecture SYN_BEHAVIORAL of FA_299 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_298 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_298;

architecture SYN_BEHAVIORAL of FA_298 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_297 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_297;

architecture SYN_BEHAVIORAL of FA_297 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_296 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_296;

architecture SYN_BEHAVIORAL of FA_296 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n5, B => Ci, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_295 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_295;

architecture SYN_BEHAVIORAL of FA_295 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n6, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_294 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_294;

architecture SYN_BEHAVIORAL of FA_294 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_293 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_293;

architecture SYN_BEHAVIORAL of FA_293 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n6, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_292 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_292;

architecture SYN_BEHAVIORAL of FA_292 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n2);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_291 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_291;

architecture SYN_BEHAVIORAL of FA_291 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_290 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_290;

architecture SYN_BEHAVIORAL of FA_290 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_289 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_289;

architecture SYN_BEHAVIORAL of FA_289 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_288 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_288;

architecture SYN_BEHAVIORAL of FA_288 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_287 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_287;

architecture SYN_BEHAVIORAL of FA_287 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_286 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_286;

architecture SYN_BEHAVIORAL of FA_286 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_285 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_285;

architecture SYN_BEHAVIORAL of FA_285 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_284 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_284;

architecture SYN_BEHAVIORAL of FA_284 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_283 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_283;

architecture SYN_BEHAVIORAL of FA_283 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_282 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_282;

architecture SYN_BEHAVIORAL of FA_282 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n8, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : INV_X1 port map( A => n7, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n8);
   U7 : XNOR2_X1 port map( A => B, B => n8, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_281 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_281;

architecture SYN_BEHAVIORAL of FA_281 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n7);
   U1 : NAND2_X1 port map( A1 => n8, A2 => A, ZN => n4);
   U2 : NAND2_X1 port map( A1 => n7, A2 => Ci, ZN => n5);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : CLKBUF_X1 port map( A => B, Z => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_280 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_280;

architecture SYN_BEHAVIORAL of FA_280 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => n5, B2 => Ci, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_279 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_279;

architecture SYN_BEHAVIORAL of FA_279 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n5, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_278 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_278;

architecture SYN_BEHAVIORAL of FA_278 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_277 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_277;

architecture SYN_BEHAVIORAL of FA_277 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_276 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_276;

architecture SYN_BEHAVIORAL of FA_276 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_275 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_275;

architecture SYN_BEHAVIORAL of FA_275 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_274 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_274;

architecture SYN_BEHAVIORAL of FA_274 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_273 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_273;

architecture SYN_BEHAVIORAL of FA_273 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_272 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_272;

architecture SYN_BEHAVIORAL of FA_272 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_271 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_271;

architecture SYN_BEHAVIORAL of FA_271 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : INV_X1 port map( A => n2, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_270 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_270;

architecture SYN_BEHAVIORAL of FA_270 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_269 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_269;

architecture SYN_BEHAVIORAL of FA_269 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n5, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_268 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_268;

architecture SYN_BEHAVIORAL of FA_268 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : XNOR2_X1 port map( A => B, B => n6, ZN => n4);
   U5 : CLKBUF_X1 port map( A => B, Z => n5);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_267 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_267;

architecture SYN_BEHAVIORAL of FA_267 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n8);
   U2 : NAND2_X1 port map( A1 => n7, A2 => A, ZN => n4);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n9, ZN => n5);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : CLKBUF_X1 port map( A => B, Z => n7);
   U7 : XNOR2_X1 port map( A => B, B => n8, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_266 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_266;

architecture SYN_BEHAVIORAL of FA_266 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_265 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_265;

architecture SYN_BEHAVIORAL of FA_265 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_264 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_264;

architecture SYN_BEHAVIORAL of FA_264 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n8);
   U2 : NAND2_X1 port map( A1 => n7, A2 => A, ZN => n4);
   U4 : NAND2_X1 port map( A1 => n9, A2 => Ci, ZN => n5);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : CLKBUF_X1 port map( A => B, Z => n7);
   U7 : XNOR2_X1 port map( A => B, B => n8, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_263 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_263;

architecture SYN_BEHAVIORAL of FA_263 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_262 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_262;

architecture SYN_BEHAVIORAL of FA_262 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : NAND2_X1 port map( A1 => n8, A2 => A, ZN => n4);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n9, ZN => n5);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n9);
   U7 : CLKBUF_X1 port map( A => B, Z => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_261 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_261;

architecture SYN_BEHAVIORAL of FA_261 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n6, B2 => Ci, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_260 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_260;

architecture SYN_BEHAVIORAL of FA_260 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_259 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_259;

architecture SYN_BEHAVIORAL of FA_259 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n6, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n6, B2 => Ci, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_258 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_258;

architecture SYN_BEHAVIORAL of FA_258 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U4 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => n4, B2 => Ci, ZN => n2);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_257 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_257;

architecture SYN_BEHAVIORAL of FA_257 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : CLKBUF_X1 port map( A => Ci, Z => n4);
   U4 : CLKBUF_X1 port map( A => n8, Z => n5);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n8);
   U7 : INV_X1 port map( A => n9, ZN => Co);
   U8 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => n5, B2 => n4, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_256 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_256;

architecture SYN_BEHAVIORAL of FA_256 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_255 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_255;

architecture SYN_BEHAVIORAL of FA_255 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_254 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_254;

architecture SYN_BEHAVIORAL of FA_254 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_253 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_253;

architecture SYN_BEHAVIORAL of FA_253 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_252 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_252;

architecture SYN_BEHAVIORAL of FA_252 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_251 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_251;

architecture SYN_BEHAVIORAL of FA_251 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_250 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_250;

architecture SYN_BEHAVIORAL of FA_250 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_249 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_249;

architecture SYN_BEHAVIORAL of FA_249 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_248 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_248;

architecture SYN_BEHAVIORAL of FA_248 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_247 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_247;

architecture SYN_BEHAVIORAL of FA_247 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_246 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_246;

architecture SYN_BEHAVIORAL of FA_246 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_245 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_245;

architecture SYN_BEHAVIORAL of FA_245 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_244 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_244;

architecture SYN_BEHAVIORAL of FA_244 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_243 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_243;

architecture SYN_BEHAVIORAL of FA_243 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_242 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_242;

architecture SYN_BEHAVIORAL of FA_242 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_241 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_241;

architecture SYN_BEHAVIORAL of FA_241 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_240 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_240;

architecture SYN_BEHAVIORAL of FA_240 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_239 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_239;

architecture SYN_BEHAVIORAL of FA_239 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_238 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_238;

architecture SYN_BEHAVIORAL of FA_238 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_237 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_237;

architecture SYN_BEHAVIORAL of FA_237 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_236 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_236;

architecture SYN_BEHAVIORAL of FA_236 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_235 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_235;

architecture SYN_BEHAVIORAL of FA_235 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_234 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_234;

architecture SYN_BEHAVIORAL of FA_234 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_233 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_233;

architecture SYN_BEHAVIORAL of FA_233 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_232 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_232;

architecture SYN_BEHAVIORAL of FA_232 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_231 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_231;

architecture SYN_BEHAVIORAL of FA_231 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_230 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_230;

architecture SYN_BEHAVIORAL of FA_230 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_229 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_229;

architecture SYN_BEHAVIORAL of FA_229 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n6, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n6, B2 => Ci, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_228 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_228;

architecture SYN_BEHAVIORAL of FA_228 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n6, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_227 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_227;

architecture SYN_BEHAVIORAL of FA_227 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_226 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_226;

architecture SYN_BEHAVIORAL of FA_226 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => n5, B => B, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_225 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_225;

architecture SYN_BEHAVIORAL of FA_225 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_224 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_224;

architecture SYN_BEHAVIORAL of FA_224 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n7, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : INV_X1 port map( A => n8, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n7);
   U7 : XNOR2_X1 port map( A => B, B => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_223 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_223;

architecture SYN_BEHAVIORAL of FA_223 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => n6, B2 => Ci, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_222 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_222;

architecture SYN_BEHAVIORAL of FA_222 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_221 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_221;

architecture SYN_BEHAVIORAL of FA_221 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_220 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_220;

architecture SYN_BEHAVIORAL of FA_220 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_219 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_219;

architecture SYN_BEHAVIORAL of FA_219 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => n5, B => B, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_218 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_218;

architecture SYN_BEHAVIORAL of FA_218 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_217 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_217;

architecture SYN_BEHAVIORAL of FA_217 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_216 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_216;

architecture SYN_BEHAVIORAL of FA_216 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_215 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_215;

architecture SYN_BEHAVIORAL of FA_215 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_214 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_214;

architecture SYN_BEHAVIORAL of FA_214 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_213 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_213;

architecture SYN_BEHAVIORAL of FA_213 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n4);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n8, ZN => n5);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_212 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_212;

architecture SYN_BEHAVIORAL of FA_212 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_211 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_211;

architecture SYN_BEHAVIORAL of FA_211 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_210 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_210;

architecture SYN_BEHAVIORAL of FA_210 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_209 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_209;

architecture SYN_BEHAVIORAL of FA_209 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_208 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_208;

architecture SYN_BEHAVIORAL of FA_208 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => n5, B => B, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_207 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_207;

architecture SYN_BEHAVIORAL of FA_207 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n2);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_206 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_206;

architecture SYN_BEHAVIORAL of FA_206 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_205 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_205;

architecture SYN_BEHAVIORAL of FA_205 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_204 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_204;

architecture SYN_BEHAVIORAL of FA_204 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n2);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_203 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_203;

architecture SYN_BEHAVIORAL of FA_203 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_202 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_202;

architecture SYN_BEHAVIORAL of FA_202 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : OAI22_X1 port map( A1 => n5, A2 => n9, B1 => n7, B2 => n6, ZN => Co);
   U4 : INV_X1 port map( A => n4, ZN => n5);
   U5 : INV_X1 port map( A => Ci, ZN => n6);
   U6 : INV_X1 port map( A => n8, ZN => n7);
   U7 : INV_X1 port map( A => A, ZN => n9);
   U8 : XNOR2_X1 port map( A => B, B => n9, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_201 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_201;

architecture SYN_BEHAVIORAL of FA_201 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_200 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_200;

architecture SYN_BEHAVIORAL of FA_200 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n5, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_199 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_199;

architecture SYN_BEHAVIORAL of FA_199 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_198 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_198;

architecture SYN_BEHAVIORAL of FA_198 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : XNOR2_X1 port map( A => B, B => n6, ZN => n4);
   U5 : CLKBUF_X1 port map( A => B, Z => n5);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_197 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_197;

architecture SYN_BEHAVIORAL of FA_197 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_196 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_196;

architecture SYN_BEHAVIORAL of FA_196 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n6, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_195 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_195;

architecture SYN_BEHAVIORAL of FA_195 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n6, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_194 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_194;

architecture SYN_BEHAVIORAL of FA_194 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : XNOR2_X1 port map( A => B, B => n6, ZN => n4);
   U4 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => n4, B2 => Ci, ZN => n2);
   U5 : CLKBUF_X1 port map( A => B, Z => n5);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_193 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_193;

architecture SYN_BEHAVIORAL of FA_193 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : CLKBUF_X1 port map( A => Ci, Z => n4);
   U4 : CLKBUF_X1 port map( A => n8, Z => n5);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n8);
   U7 : INV_X1 port map( A => n9, ZN => Co);
   U8 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => n5, B2 => n4, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_192 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_192;

architecture SYN_BEHAVIORAL of FA_192 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_191 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_191;

architecture SYN_BEHAVIORAL of FA_191 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_190 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_190;

architecture SYN_BEHAVIORAL of FA_190 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_189 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_189;

architecture SYN_BEHAVIORAL of FA_189 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_188 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_188;

architecture SYN_BEHAVIORAL of FA_188 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_187 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_187;

architecture SYN_BEHAVIORAL of FA_187 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_186 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_186;

architecture SYN_BEHAVIORAL of FA_186 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_185 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_185;

architecture SYN_BEHAVIORAL of FA_185 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_184 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_184;

architecture SYN_BEHAVIORAL of FA_184 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_183 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_183;

architecture SYN_BEHAVIORAL of FA_183 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_182 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_182;

architecture SYN_BEHAVIORAL of FA_182 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_181 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_181;

architecture SYN_BEHAVIORAL of FA_181 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_180 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_180;

architecture SYN_BEHAVIORAL of FA_180 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_179 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_179;

architecture SYN_BEHAVIORAL of FA_179 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_178 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_178;

architecture SYN_BEHAVIORAL of FA_178 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_177 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_177;

architecture SYN_BEHAVIORAL of FA_177 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_176 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_176;

architecture SYN_BEHAVIORAL of FA_176 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_175 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_175;

architecture SYN_BEHAVIORAL of FA_175 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_174 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_174;

architecture SYN_BEHAVIORAL of FA_174 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_173 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_173;

architecture SYN_BEHAVIORAL of FA_173 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_172 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_172;

architecture SYN_BEHAVIORAL of FA_172 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_171 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_171;

architecture SYN_BEHAVIORAL of FA_171 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_170 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_170;

architecture SYN_BEHAVIORAL of FA_170 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_169 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_169;

architecture SYN_BEHAVIORAL of FA_169 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_168 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_168;

architecture SYN_BEHAVIORAL of FA_168 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_167 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_167;

architecture SYN_BEHAVIORAL of FA_167 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_166 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_166;

architecture SYN_BEHAVIORAL of FA_166 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_165 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_165;

architecture SYN_BEHAVIORAL of FA_165 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => n7, Z => n5);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => n7, B2 => Ci, ZN => n8);
   U7 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_164 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_164;

architecture SYN_BEHAVIORAL of FA_164 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => n7, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n8, ZN => Co);
   U7 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => n7, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_163 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_163;

architecture SYN_BEHAVIORAL of FA_163 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n6, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_162 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_162;

architecture SYN_BEHAVIORAL of FA_162 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => n5, B => B, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n6, B2 => Ci, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_161 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_161;

architecture SYN_BEHAVIORAL of FA_161 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n6, B2 => Ci, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_160 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_160;

architecture SYN_BEHAVIORAL of FA_160 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_159 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_159;

architecture SYN_BEHAVIORAL of FA_159 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_158 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_158;

architecture SYN_BEHAVIORAL of FA_158 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_157 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_157;

architecture SYN_BEHAVIORAL of FA_157 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_156 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_156;

architecture SYN_BEHAVIORAL of FA_156 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_155 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_155;

architecture SYN_BEHAVIORAL of FA_155 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_154 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_154;

architecture SYN_BEHAVIORAL of FA_154 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_153 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_153;

architecture SYN_BEHAVIORAL of FA_153 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_152 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_152;

architecture SYN_BEHAVIORAL of FA_152 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_151 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_151;

architecture SYN_BEHAVIORAL of FA_151 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_150 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_150;

architecture SYN_BEHAVIORAL of FA_150 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U2 : INV_X1 port map( A => n5, ZN => Co);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_149 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_149;

architecture SYN_BEHAVIORAL of FA_149 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_148 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_148;

architecture SYN_BEHAVIORAL of FA_148 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : NAND2_X1 port map( A1 => n8, A2 => A, ZN => n4);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n9, ZN => n5);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n9);
   U7 : CLKBUF_X1 port map( A => B, Z => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_147 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_147;

architecture SYN_BEHAVIORAL of FA_147 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_146 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_146;

architecture SYN_BEHAVIORAL of FA_146 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_145 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_145;

architecture SYN_BEHAVIORAL of FA_145 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_144 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_144;

architecture SYN_BEHAVIORAL of FA_144 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_143 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_143;

architecture SYN_BEHAVIORAL of FA_143 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_142 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_142;

architecture SYN_BEHAVIORAL of FA_142 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_141 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_141;

architecture SYN_BEHAVIORAL of FA_141 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_140 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_140;

architecture SYN_BEHAVIORAL of FA_140 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_139 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_139;

architecture SYN_BEHAVIORAL of FA_139 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_138 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_138;

architecture SYN_BEHAVIORAL of FA_138 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n7, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : INV_X1 port map( A => n8, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n7);
   U7 : XNOR2_X1 port map( A => B, B => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_137 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_137;

architecture SYN_BEHAVIORAL of FA_137 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_136 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_136;

architecture SYN_BEHAVIORAL of FA_136 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_135 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_135;

architecture SYN_BEHAVIORAL of FA_135 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n2);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_134 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_134;

architecture SYN_BEHAVIORAL of FA_134 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : INV_X1 port map( A => n2, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n5);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_133 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_133;

architecture SYN_BEHAVIORAL of FA_133 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_132 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_132;

architecture SYN_BEHAVIORAL of FA_132 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => n4, B2 => Ci, ZN => n2);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_131 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_131;

architecture SYN_BEHAVIORAL of FA_131 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_130 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_130;

architecture SYN_BEHAVIORAL of FA_130 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_129 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_129;

architecture SYN_BEHAVIORAL of FA_129 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : CLKBUF_X1 port map( A => Ci, Z => n4);
   U4 : CLKBUF_X1 port map( A => n8, Z => n5);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n8);
   U7 : INV_X1 port map( A => n9, ZN => Co);
   U8 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => n5, B2 => n4, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_128 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_128;

architecture SYN_BEHAVIORAL of FA_128 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_127 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_127;

architecture SYN_BEHAVIORAL of FA_127 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_126 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_126;

architecture SYN_BEHAVIORAL of FA_126 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_125 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_125;

architecture SYN_BEHAVIORAL of FA_125 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_124 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_124;

architecture SYN_BEHAVIORAL of FA_124 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_123 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_123;

architecture SYN_BEHAVIORAL of FA_123 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_122 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_122;

architecture SYN_BEHAVIORAL of FA_122 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_121 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_121;

architecture SYN_BEHAVIORAL of FA_121 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_120 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_120;

architecture SYN_BEHAVIORAL of FA_120 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_119 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_119;

architecture SYN_BEHAVIORAL of FA_119 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_118 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_118;

architecture SYN_BEHAVIORAL of FA_118 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_117 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_117;

architecture SYN_BEHAVIORAL of FA_117 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_116 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_116;

architecture SYN_BEHAVIORAL of FA_116 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_115 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_115;

architecture SYN_BEHAVIORAL of FA_115 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_114 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_114;

architecture SYN_BEHAVIORAL of FA_114 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_113 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_113;

architecture SYN_BEHAVIORAL of FA_113 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_112 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_112;

architecture SYN_BEHAVIORAL of FA_112 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_111 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_111;

architecture SYN_BEHAVIORAL of FA_111 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_110 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_110;

architecture SYN_BEHAVIORAL of FA_110 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_109 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_109;

architecture SYN_BEHAVIORAL of FA_109 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_108 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_108;

architecture SYN_BEHAVIORAL of FA_108 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_107 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_107;

architecture SYN_BEHAVIORAL of FA_107 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_106 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_106;

architecture SYN_BEHAVIORAL of FA_106 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_105 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_105;

architecture SYN_BEHAVIORAL of FA_105 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_104 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_104;

architecture SYN_BEHAVIORAL of FA_104 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_103 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_103;

architecture SYN_BEHAVIORAL of FA_103 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_102 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_102;

architecture SYN_BEHAVIORAL of FA_102 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_101 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_101;

architecture SYN_BEHAVIORAL of FA_101 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_100 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_100;

architecture SYN_BEHAVIORAL of FA_100 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_99 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_99;

architecture SYN_BEHAVIORAL of FA_99 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_98 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_98;

architecture SYN_BEHAVIORAL of FA_98 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_97 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_97;

architecture SYN_BEHAVIORAL of FA_97 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => Ci, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_96 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_96;

architecture SYN_BEHAVIORAL of FA_96 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_95 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_95;

architecture SYN_BEHAVIORAL of FA_95 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_94 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_94;

architecture SYN_BEHAVIORAL of FA_94 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_93 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_93;

architecture SYN_BEHAVIORAL of FA_93 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n5, B => Ci, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_92 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_92;

architecture SYN_BEHAVIORAL of FA_92 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => Ci, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_91 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_91;

architecture SYN_BEHAVIORAL of FA_91 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_90 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_90;

architecture SYN_BEHAVIORAL of FA_90 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_89 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_89;

architecture SYN_BEHAVIORAL of FA_89 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n5, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_88 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_88;

architecture SYN_BEHAVIORAL of FA_88 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_87 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_87;

architecture SYN_BEHAVIORAL of FA_87 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_86 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_86;

architecture SYN_BEHAVIORAL of FA_86 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_85 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_85;

architecture SYN_BEHAVIORAL of FA_85 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_84 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_84;

architecture SYN_BEHAVIORAL of FA_84 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_83 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_83;

architecture SYN_BEHAVIORAL of FA_83 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n5, B => Ci, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_82 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_82;

architecture SYN_BEHAVIORAL of FA_82 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_81 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_81;

architecture SYN_BEHAVIORAL of FA_81 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n7, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : INV_X1 port map( A => n8, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n7);
   U7 : XNOR2_X1 port map( A => B, B => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_80 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_80;

architecture SYN_BEHAVIORAL of FA_80 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_79 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_79;

architecture SYN_BEHAVIORAL of FA_79 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_78 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_78;

architecture SYN_BEHAVIORAL of FA_78 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_77 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_77;

architecture SYN_BEHAVIORAL of FA_77 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_76 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_76;

architecture SYN_BEHAVIORAL of FA_76 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_75 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_75;

architecture SYN_BEHAVIORAL of FA_75 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_74 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_74;

architecture SYN_BEHAVIORAL of FA_74 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_73 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_73;

architecture SYN_BEHAVIORAL of FA_73 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_72 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_72;

architecture SYN_BEHAVIORAL of FA_72 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_71 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_71;

architecture SYN_BEHAVIORAL of FA_71 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_70 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_70;

architecture SYN_BEHAVIORAL of FA_70 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_69 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_69;

architecture SYN_BEHAVIORAL of FA_69 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n5, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => Ci, Z => n5);
   U5 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n6, ZN => n2);
   U6 : CLKBUF_X1 port map( A => B, Z => n7);
   U7 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_68 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_68;

architecture SYN_BEHAVIORAL of FA_68 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : INV_X1 port map( A => n2, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n5);
   U6 : CLKBUF_X1 port map( A => Ci, Z => n7);
   U7 : XNOR2_X1 port map( A => B, B => n6, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_67 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_67;

architecture SYN_BEHAVIORAL of FA_67 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : INV_X1 port map( A => n2, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_66 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_66;

architecture SYN_BEHAVIORAL of FA_66 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U4 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_65 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_65;

architecture SYN_BEHAVIORAL of FA_65 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n6, n7, n8, n9, n10, n11 : std_logic;

begin
   
   U1 : OR2_X1 port map( A1 => n8, A2 => n5, ZN => Co);
   U2 : AND2_X1 port map( A1 => A, A2 => n11, ZN => n5);
   U3 : CLKBUF_X1 port map( A => Ci, Z => n6);
   U4 : INV_X1 port map( A => n6, ZN => n9);
   U5 : CLKBUF_X1 port map( A => n10, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => A, ZN => n10);
   U7 : XNOR2_X1 port map( A => Ci, B => n10, ZN => S);
   U8 : NOR2_X1 port map( A1 => n9, A2 => n7, ZN => n8);
   U9 : CLKBUF_X1 port map( A => B, Z => n11);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_64 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_64;

architecture SYN_BEHAVIORAL of FA_64 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_63 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_63;

architecture SYN_BEHAVIORAL of FA_63 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_62 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_62;

architecture SYN_BEHAVIORAL of FA_62 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_61 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_61;

architecture SYN_BEHAVIORAL of FA_61 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_60 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_60;

architecture SYN_BEHAVIORAL of FA_60 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_59 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_59;

architecture SYN_BEHAVIORAL of FA_59 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_58 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_58;

architecture SYN_BEHAVIORAL of FA_58 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_57 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_57;

architecture SYN_BEHAVIORAL of FA_57 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_56 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_56;

architecture SYN_BEHAVIORAL of FA_56 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_55 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_55;

architecture SYN_BEHAVIORAL of FA_55 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_54 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_54;

architecture SYN_BEHAVIORAL of FA_54 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_53 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_53;

architecture SYN_BEHAVIORAL of FA_53 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_52 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_52;

architecture SYN_BEHAVIORAL of FA_52 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_51 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_51;

architecture SYN_BEHAVIORAL of FA_51 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_50 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_50;

architecture SYN_BEHAVIORAL of FA_50 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_49 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_49;

architecture SYN_BEHAVIORAL of FA_49 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_48 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_48;

architecture SYN_BEHAVIORAL of FA_48 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_47 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_47;

architecture SYN_BEHAVIORAL of FA_47 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_46 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_46;

architecture SYN_BEHAVIORAL of FA_46 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_45 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_45;

architecture SYN_BEHAVIORAL of FA_45 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_44 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_44;

architecture SYN_BEHAVIORAL of FA_44 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_43 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_43;

architecture SYN_BEHAVIORAL of FA_43 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_42 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_42;

architecture SYN_BEHAVIORAL of FA_42 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_41 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_41;

architecture SYN_BEHAVIORAL of FA_41 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_40 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_40;

architecture SYN_BEHAVIORAL of FA_40 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_39 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_39;

architecture SYN_BEHAVIORAL of FA_39 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_38 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_38;

architecture SYN_BEHAVIORAL of FA_38 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_37 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_37;

architecture SYN_BEHAVIORAL of FA_37 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_36 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_36;

architecture SYN_BEHAVIORAL of FA_36 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_35 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_35;

architecture SYN_BEHAVIORAL of FA_35 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_34 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_34;

architecture SYN_BEHAVIORAL of FA_34 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_33 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_33;

architecture SYN_BEHAVIORAL of FA_33 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_32 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_32;

architecture SYN_BEHAVIORAL of FA_32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_31 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_31;

architecture SYN_BEHAVIORAL of FA_31 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_30 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_30;

architecture SYN_BEHAVIORAL of FA_30 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_29 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_29;

architecture SYN_BEHAVIORAL of FA_29 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U1 : CLKBUF_X1 port map( A => Ci, Z => n4);
   U2 : CLKBUF_X1 port map( A => n6, Z => n5);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n6, B2 => Ci, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_28 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_28;

architecture SYN_BEHAVIORAL of FA_28 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : CLKBUF_X1 port map( A => n5, Z => n4);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_27 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_27;

architecture SYN_BEHAVIORAL of FA_27 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : CLKBUF_X1 port map( A => Ci, Z => n4);
   U2 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_26 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_26;

architecture SYN_BEHAVIORAL of FA_26 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n5, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => Ci, Z => n5);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_25 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_25;

architecture SYN_BEHAVIORAL of FA_25 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_24 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_24;

architecture SYN_BEHAVIORAL of FA_24 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => n6, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n6);
   U1 : CLKBUF_X1 port map( A => Ci, Z => n4);
   U2 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => n6, B2 => Ci, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_23 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_23;

architecture SYN_BEHAVIORAL of FA_23 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : CLKBUF_X1 port map( A => n5, Z => n4);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_22 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_22;

architecture SYN_BEHAVIORAL of FA_22 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_21 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_21;

architecture SYN_BEHAVIORAL of FA_21 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_20 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_20;

architecture SYN_BEHAVIORAL of FA_20 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : CLKBUF_X1 port map( A => Ci, Z => n4);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_19 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_19;

architecture SYN_BEHAVIORAL of FA_19 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n6);
   U4 : CLKBUF_X1 port map( A => n6, Z => n5);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_18 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_18;

architecture SYN_BEHAVIORAL of FA_18 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U1 : CLKBUF_X1 port map( A => Ci, Z => n4);
   U2 : CLKBUF_X1 port map( A => n6, Z => n5);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_17 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_17;

architecture SYN_BEHAVIORAL of FA_17 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : CLKBUF_X1 port map( A => Ci, Z => n4);
   U2 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_16 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_16;

architecture SYN_BEHAVIORAL of FA_16 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : CLKBUF_X1 port map( A => Ci, Z => n4);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_15 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_15;

architecture SYN_BEHAVIORAL of FA_15 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n6);
   U1 : CLKBUF_X1 port map( A => Ci, Z => n4);
   U2 : CLKBUF_X1 port map( A => n6, Z => n5);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n6, B2 => Ci, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_14 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_14;

architecture SYN_BEHAVIORAL of FA_14 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_13 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_13;

architecture SYN_BEHAVIORAL of FA_13 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : CLKBUF_X1 port map( A => n5, Z => n4);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_12 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_12;

architecture SYN_BEHAVIORAL of FA_12 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_11 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_11;

architecture SYN_BEHAVIORAL of FA_11 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n6, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U4 : XNOR2_X1 port map( A => n5, B => B, ZN => n8);
   U5 : CLKBUF_X1 port map( A => Ci, Z => n6);
   U6 : CLKBUF_X1 port map( A => B, Z => n7);
   U7 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n8, ZN => n9);
   U8 : INV_X1 port map( A => n9, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_10 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_10;

architecture SYN_BEHAVIORAL of FA_10 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : CLKBUF_X1 port map( A => Ci, Z => n4);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_9 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_9;

architecture SYN_BEHAVIORAL of FA_9 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n5, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n6);
   U1 : CLKBUF_X1 port map( A => n6, Z => n4);
   U2 : CLKBUF_X1 port map( A => Ci, Z => n5);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_8 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_8;

architecture SYN_BEHAVIORAL of FA_8 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n5, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : CLKBUF_X1 port map( A => Ci, Z => n4);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_7 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_7;

architecture SYN_BEHAVIORAL of FA_7 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n5, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => Ci, Z => n5);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_6 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_6;

architecture SYN_BEHAVIORAL of FA_6 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n7, n8, n9, n10 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => n8, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n10);
   U1 : NAND2_X1 port map( A1 => n9, A2 => A, ZN => n4);
   U2 : NAND2_X1 port map( A1 => Ci, A2 => n10, ZN => n5);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : CLKBUF_X1 port map( A => n10, Z => n7);
   U7 : CLKBUF_X1 port map( A => Ci, Z => n8);
   U8 : CLKBUF_X1 port map( A => B, Z => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_5 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_5;

architecture SYN_BEHAVIORAL of FA_5 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal net162483, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => net162483, Z => S);
   U1 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U2 : NOR2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : AOI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n6);
   U5 : NOR2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U6 : CLKBUF_X1 port map( A => Ci, Z => net162483);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_4 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_4;

architecture SYN_BEHAVIORAL of FA_4 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal net154226, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => net154226, B => n4, Z => S);
   U1 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U2 : NOR2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : AOI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n6);
   U5 : NOR2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U6 : CLKBUF_X1 port map( A => Ci, Z => net154226);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_3 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_3;

architecture SYN_BEHAVIORAL of FA_3 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal net154429, net154985, n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => net154429, B => net154985, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => n4, B2 => Ci, ZN => n2);
   U4 : INV_X1 port map( A => n2, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n5);
   U6 : CLKBUF_X1 port map( A => Ci, Z => net154429);
   U7 : XNOR2_X1 port map( A => B, B => n6, ZN => n4);
   U8 : CLKBUF_X1 port map( A => n4, Z => net154985);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_2 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2;

architecture SYN_BEHAVIORAL of FA_2 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal net155512, net156196, net156195, n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => net155512, B => n4, Z => S);
   U1 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U2 : AND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NOR2_X1 port map( A1 => n5, A2 => Ci, ZN => net156196);
   U5 : NOR2_X1 port map( A1 => A, A2 => B, ZN => net156195);
   U6 : NOR2_X1 port map( A1 => net156196, A2 => net156195, ZN => Co);
   U7 : CLKBUF_X1 port map( A => Ci, Z => net155512);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_1 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1;

architecture SYN_BEHAVIORAL of FA_1 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net150614, net177427, net177422, n5, n6, n7, n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => net150614, ZN => net177422);
   U2 : OR2_X1 port map( A1 => n8, A2 => n5, ZN => Co);
   U3 : AND2_X1 port map( A1 => A, A2 => n7, ZN => n5);
   U4 : XNOR2_X1 port map( A => n6, B => Ci, ZN => S);
   U5 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U6 : CLKBUF_X1 port map( A => n6, Z => net177427);
   U7 : CLKBUF_X1 port map( A => Ci, Z => net150614);
   U8 : CLKBUF_X1 port map( A => B, Z => n7);
   U9 : NOR2_X1 port map( A1 => net177427, A2 => net177422, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity MUX51_MuxNbit64_15 is

   port( zeroSignal, A_signal, A_neg, A_shifted, A_neg_shifted : in 
         std_logic_vector (63 downto 0);  Sel : in std_logic_vector (2 downto 
         0);  Y : out std_logic_vector (63 downto 0));

end MUX51_MuxNbit64_15;

architecture SYN_BEHAVIORAL_2 of MUX51_MuxNbit64_15 is

   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X3
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X4
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, 
      n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, 
      n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, 
      n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, 
      n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, 
      n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, 
      n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, 
      n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, 
      n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, 
      n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, 
      n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, 
      n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, 
      n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, 
      n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, 
      n308 : std_logic;

begin
   
   U1 : NOR3_X1 port map( A1 => n307, A2 => Sel(2), A3 => n308, ZN => n145);
   U2 : CLKBUF_X3 port map( A => n301, Z => n151);
   U3 : BUF_X1 port map( A => n145, Z => n173);
   U4 : BUF_X1 port map( A => n158, Z => n157);
   U5 : BUF_X1 port map( A => Sel(1), Z => n144);
   U6 : OR3_X1 port map( A1 => n307, A2 => Sel(2), A3 => Sel(1), ZN => n141);
   U7 : INV_X4 port map( A => n141, ZN => n150);
   U8 : NOR3_X2 port map( A1 => n307, A2 => Sel(2), A3 => n144, ZN => n301);
   U9 : CLKBUF_X1 port map( A => n172, Z => n170);
   U10 : BUF_X4 port map( A => n173, Z => n169);
   U11 : CLKBUF_X1 port map( A => n145, Z => n172);
   U12 : CLKBUF_X1 port map( A => n173, Z => n171);
   U13 : INV_X1 port map( A => n144, ZN => n142);
   U14 : INV_X1 port map( A => Sel(0), ZN => n143);
   U15 : CLKBUF_X3 port map( A => n157, Z => n156);
   U16 : CLKBUF_X1 port map( A => n157, Z => n155);
   U17 : CLKBUF_X3 port map( A => n157, Z => n154);
   U18 : CLKBUF_X1 port map( A => n303, Z => n148);
   U19 : BUF_X1 port map( A => n167, Z => n165);
   U20 : CLKBUF_X3 port map( A => n148, Z => n147);
   U21 : BUF_X1 port map( A => n166, Z => n161);
   U22 : BUF_X1 port map( A => n165, Z => n163);
   U23 : BUF_X1 port map( A => n166, Z => n160);
   U24 : BUF_X1 port map( A => n165, Z => n162);
   U25 : BUF_X1 port map( A => n166, Z => n159);
   U26 : BUF_X1 port map( A => n165, Z => n164);
   U27 : BUF_X1 port map( A => n167, Z => n166);
   U28 : BUF_X1 port map( A => n302, Z => n158);
   U29 : AND3_X1 port map( A1 => n307, A2 => n308, A3 => Sel(2), ZN => n303);
   U30 : BUF_X1 port map( A => n304, Z => n167);
   U31 : NOR2_X1 port map( A1 => n147, A2 => n174, ZN => n304);
   U32 : AOI222_X1 port map( A1 => A_shifted(2), A2 => n171, B1 => 
                           zeroSignal(2), B2 => n160, C1 => A_neg_shifted(2), 
                           C2 => n147, ZN => n219);
   U33 : AOI22_X1 port map( A1 => A_neg(39), A2 => n156, B1 => A_signal(39), B2
                           => n150, ZN => n240);
   U34 : AOI222_X1 port map( A1 => A_shifted(4), A2 => n172, B1 => 
                           zeroSignal(4), B2 => n162, C1 => A_neg_shifted(4), 
                           C2 => n303, ZN => n263);
   U35 : NAND2_X1 port map( A1 => n244, A2 => n243, ZN => Y(40));
   U36 : AOI22_X1 port map( A1 => A_neg(40), A2 => n156, B1 => A_signal(40), B2
                           => n151, ZN => n244);
   U37 : NAND2_X1 port map( A1 => n188, A2 => n187, ZN => Y(15));
   U38 : AOI22_X1 port map( A1 => A_neg(15), A2 => n154, B1 => A_signal(15), B2
                           => n150, ZN => n188);
   U39 : NAND2_X1 port map( A1 => n250, A2 => n249, ZN => Y(43));
   U40 : AOI22_X1 port map( A1 => A_neg(43), A2 => n154, B1 => A_signal(43), B2
                           => n151, ZN => n250);
   U41 : NAND2_X1 port map( A1 => n184, A2 => n183, ZN => Y(13));
   U42 : NAND2_X1 port map( A1 => n192, A2 => n191, ZN => Y(17));
   U43 : AOI222_X1 port map( A1 => A_shifted(17), A2 => n169, B1 => 
                           zeroSignal(17), B2 => n159, C1 => A_neg_shifted(17),
                           C2 => n147, ZN => n191);
   U44 : AOI22_X1 port map( A1 => A_neg(17), A2 => n154, B1 => A_signal(17), B2
                           => n150, ZN => n192);
   U45 : NAND2_X1 port map( A1 => n190, A2 => n189, ZN => Y(16));
   U46 : AOI222_X1 port map( A1 => A_shifted(16), A2 => n169, B1 => 
                           zeroSignal(16), B2 => n159, C1 => A_neg_shifted(16),
                           C2 => n147, ZN => n189);
   U47 : AOI22_X1 port map( A1 => A_neg(16), A2 => n154, B1 => A_signal(16), B2
                           => n151, ZN => n190);
   U48 : NAND2_X1 port map( A1 => n186, A2 => n185, ZN => Y(14));
   U49 : NAND2_X1 port map( A1 => n194, A2 => n193, ZN => Y(18));
   U50 : AOI222_X1 port map( A1 => A_shifted(18), A2 => n169, B1 => 
                           zeroSignal(18), B2 => n159, C1 => A_neg_shifted(18),
                           C2 => n147, ZN => n193);
   U51 : AOI22_X1 port map( A1 => A_neg(18), A2 => n154, B1 => A_signal(18), B2
                           => n150, ZN => n194);
   U52 : NAND2_X1 port map( A1 => n196, A2 => n195, ZN => Y(19));
   U53 : AOI222_X1 port map( A1 => A_shifted(19), A2 => n169, B1 => 
                           zeroSignal(19), B2 => n159, C1 => A_neg_shifted(19),
                           C2 => n147, ZN => n195);
   U54 : AOI22_X1 port map( A1 => A_neg(19), A2 => n154, B1 => A_signal(19), B2
                           => n151, ZN => n196);
   U55 : NAND2_X1 port map( A1 => n274, A2 => n273, ZN => Y(54));
   U56 : AOI222_X1 port map( A1 => A_shifted(54), A2 => n168, B1 => 
                           zeroSignal(54), B2 => n163, C1 => A_neg_shifted(54),
                           C2 => n147, ZN => n273);
   U57 : AOI22_X1 port map( A1 => A_neg(54), A2 => n154, B1 => A_signal(54), B2
                           => n150, ZN => n274);
   U58 : NAND2_X1 port map( A1 => n272, A2 => n271, ZN => Y(53));
   U59 : AOI222_X1 port map( A1 => A_shifted(53), A2 => n171, B1 => 
                           zeroSignal(53), B2 => n163, C1 => A_neg_shifted(53),
                           C2 => n147, ZN => n271);
   U60 : AOI22_X1 port map( A1 => A_neg(53), A2 => n156, B1 => A_signal(53), B2
                           => n150, ZN => n272);
   U61 : NAND2_X1 port map( A1 => n276, A2 => n275, ZN => Y(55));
   U62 : AOI222_X1 port map( A1 => A_shifted(55), A2 => n169, B1 => 
                           zeroSignal(55), B2 => n163, C1 => A_neg_shifted(55),
                           C2 => n147, ZN => n275);
   U63 : AOI22_X1 port map( A1 => A_neg(55), A2 => n156, B1 => A_signal(55), B2
                           => n151, ZN => n276);
   U64 : NAND2_X1 port map( A1 => n256, A2 => n255, ZN => Y(46));
   U65 : AOI222_X1 port map( A1 => A_shifted(46), A2 => n169, B1 => 
                           zeroSignal(46), B2 => n162, C1 => A_neg_shifted(46),
                           C2 => n147, ZN => n255);
   U66 : AOI22_X1 port map( A1 => A_neg(46), A2 => n154, B1 => A_signal(46), B2
                           => n151, ZN => n256);
   U67 : NAND2_X1 port map( A1 => n202, A2 => n201, ZN => Y(21));
   U68 : AOI22_X1 port map( A1 => A_neg(21), A2 => n154, B1 => A_signal(21), B2
                           => n150, ZN => n202);
   U69 : NAND2_X1 port map( A1 => n278, A2 => n277, ZN => Y(56));
   U70 : AOI222_X1 port map( A1 => A_shifted(56), A2 => n171, B1 => 
                           zeroSignal(56), B2 => n163, C1 => A_neg_shifted(56),
                           C2 => n147, ZN => n277);
   U71 : AOI22_X1 port map( A1 => A_neg(56), A2 => n156, B1 => A_signal(56), B2
                           => n150, ZN => n278);
   U72 : NAND2_X1 port map( A1 => n254, A2 => n253, ZN => Y(45));
   U73 : AOI22_X1 port map( A1 => A_neg(45), A2 => n156, B1 => A_signal(45), B2
                           => n150, ZN => n254);
   U74 : NAND2_X1 port map( A1 => n280, A2 => n279, ZN => Y(57));
   U75 : AOI222_X1 port map( A1 => A_shifted(57), A2 => n168, B1 => 
                           zeroSignal(57), B2 => n163, C1 => A_neg_shifted(57),
                           C2 => n147, ZN => n279);
   U76 : AOI22_X1 port map( A1 => A_neg(57), A2 => n154, B1 => A_signal(57), B2
                           => n150, ZN => n280);
   U77 : NAND2_X1 port map( A1 => n204, A2 => n203, ZN => Y(22));
   U78 : AOI222_X1 port map( A1 => A_shifted(22), A2 => n169, B1 => 
                           zeroSignal(22), B2 => n160, C1 => A_neg_shifted(22),
                           C2 => n147, ZN => n203);
   U79 : AOI22_X1 port map( A1 => A_neg(22), A2 => n154, B1 => A_signal(22), B2
                           => n151, ZN => n204);
   U80 : NAND2_X1 port map( A1 => n258, A2 => n257, ZN => Y(47));
   U81 : AOI222_X1 port map( A1 => A_shifted(47), A2 => n171, B1 => 
                           zeroSignal(47), B2 => n162, C1 => A_neg_shifted(47),
                           C2 => n147, ZN => n257);
   U82 : NAND2_X1 port map( A1 => n282, A2 => n281, ZN => Y(58));
   U83 : AOI222_X1 port map( A1 => A_shifted(58), A2 => n169, B1 => 
                           zeroSignal(58), B2 => n163, C1 => A_neg_shifted(58),
                           C2 => n147, ZN => n281);
   U84 : AOI22_X1 port map( A1 => A_neg(58), A2 => n156, B1 => A_signal(58), B2
                           => n151, ZN => n282);
   U85 : NAND2_X1 port map( A1 => n206, A2 => n205, ZN => Y(23));
   U86 : AOI222_X1 port map( A1 => A_shifted(23), A2 => n169, B1 => 
                           zeroSignal(23), B2 => n160, C1 => A_neg_shifted(23),
                           C2 => n147, ZN => n205);
   U87 : AOI22_X1 port map( A1 => A_neg(23), A2 => n154, B1 => A_signal(23), B2
                           => n150, ZN => n206);
   U88 : NAND2_X1 port map( A1 => n200, A2 => n199, ZN => Y(20));
   U89 : AOI222_X1 port map( A1 => A_shifted(20), A2 => n169, B1 => 
                           zeroSignal(20), B2 => n160, C1 => A_neg_shifted(20),
                           C2 => n147, ZN => n199);
   U90 : NAND2_X1 port map( A1 => n208, A2 => n207, ZN => Y(24));
   U91 : AOI222_X1 port map( A1 => A_shifted(24), A2 => n169, B1 => 
                           zeroSignal(24), B2 => n160, C1 => A_neg_shifted(24),
                           C2 => n147, ZN => n207);
   U92 : AOI22_X1 port map( A1 => A_neg(24), A2 => n156, B1 => A_signal(24), B2
                           => n150, ZN => n208);
   U93 : NAND2_X1 port map( A1 => n284, A2 => n283, ZN => Y(59));
   U94 : AOI222_X1 port map( A1 => A_shifted(59), A2 => n168, B1 => 
                           zeroSignal(59), B2 => n163, C1 => A_neg_shifted(59),
                           C2 => n147, ZN => n283);
   U95 : AOI22_X1 port map( A1 => A_neg(59), A2 => n155, B1 => A_signal(59), B2
                           => n150, ZN => n284);
   U96 : NAND2_X1 port map( A1 => n210, A2 => n209, ZN => Y(25));
   U97 : AOI222_X1 port map( A1 => A_shifted(25), A2 => n168, B1 => 
                           zeroSignal(25), B2 => n160, C1 => A_neg_shifted(25),
                           C2 => n147, ZN => n209);
   U98 : AOI22_X1 port map( A1 => A_neg(25), A2 => n156, B1 => A_signal(25), B2
                           => n151, ZN => n210);
   U99 : NAND2_X1 port map( A1 => n252, A2 => n251, ZN => Y(44));
   U100 : NAND2_X1 port map( A1 => n292, A2 => n291, ZN => Y(62));
   U101 : AOI222_X1 port map( A1 => A_shifted(62), A2 => n168, B1 => 
                           zeroSignal(62), B2 => n163, C1 => A_neg_shifted(62),
                           C2 => n147, ZN => n291);
   U102 : AOI22_X1 port map( A1 => A_neg(62), A2 => n156, B1 => A_signal(62), 
                           B2 => n150, ZN => n292);
   U103 : NAND2_X1 port map( A1 => n212, A2 => n211, ZN => Y(26));
   U104 : AOI222_X1 port map( A1 => A_shifted(26), A2 => n169, B1 => 
                           zeroSignal(26), B2 => n160, C1 => A_neg_shifted(26),
                           C2 => n147, ZN => n211);
   U105 : AOI22_X1 port map( A1 => A_neg(26), A2 => n154, B1 => A_signal(26), 
                           B2 => n150, ZN => n212);
   U106 : NAND2_X1 port map( A1 => n214, A2 => n213, ZN => Y(27));
   U107 : AOI222_X1 port map( A1 => A_shifted(27), A2 => n168, B1 => 
                           zeroSignal(27), B2 => n160, C1 => A_neg_shifted(27),
                           C2 => n147, ZN => n213);
   U108 : AOI22_X1 port map( A1 => A_neg(27), A2 => n156, B1 => A_signal(27), 
                           B2 => n150, ZN => n214);
   U109 : NAND2_X1 port map( A1 => n288, A2 => n287, ZN => Y(60));
   U110 : AOI222_X1 port map( A1 => A_shifted(60), A2 => n169, B1 => 
                           zeroSignal(60), B2 => n163, C1 => A_neg_shifted(60),
                           C2 => n147, ZN => n287);
   U111 : AOI22_X1 port map( A1 => A_neg(60), A2 => n156, B1 => A_signal(60), 
                           B2 => n150, ZN => n288);
   U112 : NAND2_X1 port map( A1 => n290, A2 => n289, ZN => Y(61));
   U113 : AOI222_X1 port map( A1 => A_shifted(61), A2 => n171, B1 => 
                           zeroSignal(61), B2 => n163, C1 => A_neg_shifted(61),
                           C2 => n147, ZN => n289);
   U114 : AOI22_X1 port map( A1 => A_neg(61), A2 => n154, B1 => A_signal(61), 
                           B2 => n151, ZN => n290);
   U115 : NAND2_X1 port map( A1 => n218, A2 => n217, ZN => Y(29));
   U116 : AOI222_X1 port map( A1 => A_shifted(29), A2 => n168, B1 => 
                           zeroSignal(29), B2 => n160, C1 => A_neg_shifted(29),
                           C2 => n147, ZN => n217);
   U117 : AOI22_X1 port map( A1 => A_neg(29), A2 => n154, B1 => A_signal(29), 
                           B2 => n150, ZN => n218);
   U118 : NAND2_X1 port map( A1 => n216, A2 => n215, ZN => Y(28));
   U119 : AOI222_X1 port map( A1 => A_shifted(28), A2 => n169, B1 => 
                           zeroSignal(28), B2 => n160, C1 => A_neg_shifted(28),
                           C2 => n147, ZN => n215);
   U120 : AOI22_X1 port map( A1 => A_neg(28), A2 => n156, B1 => A_signal(28), 
                           B2 => n151, ZN => n216);
   U121 : NAND2_X1 port map( A1 => n294, A2 => n293, ZN => Y(63));
   U122 : AOI222_X1 port map( A1 => A_shifted(63), A2 => n169, B1 => 
                           zeroSignal(63), B2 => n163, C1 => A_neg_shifted(63),
                           C2 => n147, ZN => n293);
   U123 : AOI22_X1 port map( A1 => A_neg(63), A2 => n155, B1 => A_signal(63), 
                           B2 => n150, ZN => n294);
   U124 : NAND2_X1 port map( A1 => n222, A2 => n221, ZN => Y(30));
   U125 : AOI222_X1 port map( A1 => A_shifted(30), A2 => n169, B1 => 
                           zeroSignal(30), B2 => n160, C1 => A_neg_shifted(30),
                           C2 => n147, ZN => n221);
   U126 : AOI22_X1 port map( A1 => A_neg(30), A2 => n156, B1 => A_signal(30), 
                           B2 => n150, ZN => n222);
   U127 : NAND2_X1 port map( A1 => n260, A2 => n259, ZN => Y(48));
   U128 : AOI22_X1 port map( A1 => A_neg(48), A2 => n156, B1 => A_signal(48), 
                           B2 => n150, ZN => n260);
   U129 : NAND2_X1 port map( A1 => n262, A2 => n261, ZN => Y(49));
   U130 : AOI222_X1 port map( A1 => A_shifted(49), A2 => n169, B1 => 
                           zeroSignal(49), B2 => n162, C1 => A_neg_shifted(49),
                           C2 => n147, ZN => n261);
   U131 : AOI22_X1 port map( A1 => A_neg(49), A2 => n154, B1 => A_signal(49), 
                           B2 => n151, ZN => n262);
   U132 : NAND2_X1 port map( A1 => n226, A2 => n225, ZN => Y(32));
   U133 : AOI22_X1 port map( A1 => A_neg(32), A2 => n156, B1 => A_signal(32), 
                           B2 => n150, ZN => n226);
   U134 : NAND2_X1 port map( A1 => n230, A2 => n229, ZN => Y(34));
   U135 : AOI222_X1 port map( A1 => A_shifted(34), A2 => n168, B1 => 
                           zeroSignal(34), B2 => n161, C1 => A_neg_shifted(34),
                           C2 => n147, ZN => n229);
   U136 : AOI22_X1 port map( A1 => A_neg(34), A2 => n156, B1 => A_signal(34), 
                           B2 => n151, ZN => n230);
   U137 : NAND2_X1 port map( A1 => n246, A2 => n245, ZN => Y(41));
   U138 : NAND2_X1 port map( A1 => n228, A2 => n227, ZN => Y(33));
   U139 : AOI222_X1 port map( A1 => A_shifted(33), A2 => n169, B1 => 
                           zeroSignal(33), B2 => n161, C1 => A_neg_shifted(33),
                           C2 => n147, ZN => n227);
   U140 : AOI22_X1 port map( A1 => A_neg(33), A2 => n154, B1 => A_signal(33), 
                           B2 => n150, ZN => n228);
   U141 : NAND2_X1 port map( A1 => n224, A2 => n223, ZN => Y(31));
   U142 : AOI222_X1 port map( A1 => A_shifted(31), A2 => n168, B1 => 
                           zeroSignal(31), B2 => n161, C1 => A_neg_shifted(31),
                           C2 => n147, ZN => n223);
   U143 : NAND2_X1 port map( A1 => n268, A2 => n267, ZN => Y(51));
   U144 : AOI222_X1 port map( A1 => A_shifted(51), A2 => n168, B1 => 
                           zeroSignal(51), B2 => n162, C1 => A_neg_shifted(51),
                           C2 => n147, ZN => n267);
   U145 : AOI22_X1 port map( A1 => A_neg(51), A2 => n156, B1 => A_signal(51), 
                           B2 => n150, ZN => n268);
   U146 : NAND2_X1 port map( A1 => n232, A2 => n231, ZN => Y(35));
   U147 : AOI22_X1 port map( A1 => A_neg(35), A2 => n154, B1 => A_signal(35), 
                           B2 => n150, ZN => n232);
   U148 : NAND2_X1 port map( A1 => n266, A2 => n265, ZN => Y(50));
   U149 : AOI222_X1 port map( A1 => A_shifted(50), A2 => n171, B1 => 
                           zeroSignal(50), B2 => n162, C1 => A_neg_shifted(50),
                           C2 => n147, ZN => n265);
   U150 : NAND2_X1 port map( A1 => n270, A2 => n269, ZN => Y(52));
   U151 : AOI222_X1 port map( A1 => A_shifted(52), A2 => n169, B1 => 
                           zeroSignal(52), B2 => n162, C1 => A_neg_shifted(52),
                           C2 => n147, ZN => n269);
   U152 : AOI22_X1 port map( A1 => A_neg(52), A2 => n154, B1 => A_signal(52), 
                           B2 => n151, ZN => n270);
   U153 : NAND2_X1 port map( A1 => n234, A2 => n233, ZN => Y(36));
   U154 : AOI22_X1 port map( A1 => A_neg(36), A2 => n156, B1 => A_signal(36), 
                           B2 => n150, ZN => n234);
   U155 : NAND2_X1 port map( A1 => n236, A2 => n235, ZN => Y(37));
   U156 : AOI22_X1 port map( A1 => A_neg(37), A2 => n156, B1 => A_signal(37), 
                           B2 => n151, ZN => n236);
   U157 : NAND2_X1 port map( A1 => n248, A2 => n247, ZN => Y(42));
   U158 : AOI22_X1 port map( A1 => A_neg(42), A2 => n156, B1 => A_signal(42), 
                           B2 => n150, ZN => n248);
   U159 : NAND2_X1 port map( A1 => n238, A2 => n237, ZN => Y(38));
   U160 : AOI22_X1 port map( A1 => A_neg(38), A2 => n154, B1 => A_signal(38), 
                           B2 => n150, ZN => n238);
   U161 : NAND2_X1 port map( A1 => n176, A2 => n175, ZN => Y(0));
   U162 : AOI22_X1 port map( A1 => A_neg(0), A2 => n156, B1 => A_signal(0), B2 
                           => n150, ZN => n176);
   U163 : AOI222_X1 port map( A1 => A_shifted(0), A2 => n168, B1 => 
                           zeroSignal(0), B2 => n159, C1 => A_neg_shifted(0), 
                           C2 => n147, ZN => n175);
   U164 : NAND2_X1 port map( A1 => n198, A2 => n197, ZN => Y(1));
   U165 : AOI22_X1 port map( A1 => A_neg(1), A2 => n154, B1 => A_signal(1), B2 
                           => n151, ZN => n198);
   U166 : AOI222_X1 port map( A1 => A_shifted(1), A2 => n169, B1 => 
                           zeroSignal(1), B2 => n159, C1 => A_neg_shifted(1), 
                           C2 => n147, ZN => n197);
   U167 : AOI222_X1 port map( A1 => A_shifted(13), A2 => n169, B1 => 
                           zeroSignal(13), B2 => n159, C1 => A_neg_shifted(13),
                           C2 => n146, ZN => n183);
   U168 : AOI22_X1 port map( A1 => A_neg(12), A2 => n156, B1 => A_signal(12), 
                           B2 => n150, ZN => n182);
   U169 : NAND2_X1 port map( A1 => n178, A2 => n177, ZN => Y(10));
   U170 : AOI222_X1 port map( A1 => A_shifted(5), A2 => n173, B1 => 
                           zeroSignal(5), B2 => n163, C1 => A_neg_shifted(5), 
                           C2 => n303, ZN => n285);
   U171 : AOI222_X1 port map( A1 => A_shifted(15), A2 => n169, B1 => 
                           zeroSignal(15), B2 => n159, C1 => A_neg_shifted(15),
                           C2 => n147, ZN => n187);
   U172 : AOI22_X1 port map( A1 => A_neg(14), A2 => n154, B1 => A_signal(14), 
                           B2 => n150, ZN => n186);
   U173 : NAND2_X1 port map( A1 => n182, A2 => n181, ZN => Y(12));
   U174 : CLKBUF_X1 port map( A => n303, Z => n149);
   U175 : BUF_X1 port map( A => n149, Z => n146);
   U176 : AOI22_X1 port map( A1 => A_neg(50), A2 => n156, B1 => A_signal(50), 
                           B2 => n150, ZN => n266);
   U177 : AOI222_X1 port map( A1 => A_shifted(14), A2 => n169, B1 => 
                           zeroSignal(14), B2 => n159, C1 => A_neg_shifted(14),
                           C2 => n147, ZN => n185);
   U178 : AOI22_X1 port map( A1 => A_neg(13), A2 => n154, B1 => A_signal(13), 
                           B2 => n151, ZN => n184);
   U179 : NAND2_X1 port map( A1 => n180, A2 => n179, ZN => Y(11));
   U180 : AOI222_X1 port map( A1 => A_shifted(11), A2 => n169, B1 => 
                           zeroSignal(11), B2 => n159, C1 => A_neg_shifted(11),
                           C2 => n146, ZN => n179);
   U181 : AOI22_X1 port map( A1 => A_neg(10), A2 => n155, B1 => A_signal(10), 
                           B2 => n151, ZN => n178);
   U182 : NAND2_X1 port map( A1 => n300, A2 => n299, ZN => Y(8));
   U183 : AOI222_X1 port map( A1 => A_shifted(12), A2 => n169, B1 => 
                           zeroSignal(12), B2 => n159, C1 => A_neg_shifted(12),
                           C2 => n146, ZN => n181);
   U184 : AOI22_X1 port map( A1 => A_neg(11), A2 => n155, B1 => A_signal(11), 
                           B2 => n150, ZN => n180);
   U185 : NAND2_X1 port map( A1 => n306, A2 => n305, ZN => Y(9));
   U186 : AOI222_X1 port map( A1 => A_shifted(10), A2 => n168, B1 => 
                           zeroSignal(10), B2 => n159, C1 => A_neg_shifted(10),
                           C2 => n148, ZN => n177);
   U187 : AOI22_X1 port map( A1 => A_neg(9), A2 => n155, B1 => A_signal(9), B2 
                           => n150, ZN => n306);
   U188 : NAND2_X1 port map( A1 => n298, A2 => n297, ZN => Y(7));
   U189 : AOI222_X1 port map( A1 => A_shifted(9), A2 => n171, B1 => 
                           zeroSignal(9), B2 => n164, C1 => A_neg_shifted(9), 
                           C2 => n148, ZN => n305);
   U190 : AOI22_X1 port map( A1 => A_neg(8), A2 => n155, B1 => A_signal(8), B2 
                           => n150, ZN => n300);
   U191 : NAND2_X1 port map( A1 => n296, A2 => n295, ZN => Y(6));
   U192 : AOI222_X1 port map( A1 => A_shifted(6), A2 => n170, B1 => 
                           zeroSignal(6), B2 => n164, C1 => A_neg_shifted(6), 
                           C2 => n303, ZN => n295);
   U193 : NAND2_X1 port map( A1 => n286, A2 => n285, ZN => Y(5));
   U194 : AOI222_X1 port map( A1 => A_shifted(44), A2 => n169, B1 => 
                           zeroSignal(44), B2 => n162, C1 => A_neg_shifted(44),
                           C2 => n147, ZN => n251);
   U195 : AOI222_X1 port map( A1 => A_shifted(43), A2 => n168, B1 => 
                           zeroSignal(43), B2 => n162, C1 => A_neg_shifted(43),
                           C2 => n147, ZN => n249);
   U196 : AOI222_X1 port map( A1 => A_shifted(41), A2 => n168, B1 => 
                           zeroSignal(41), B2 => n161, C1 => A_neg_shifted(41),
                           C2 => n147, ZN => n245);
   U197 : AOI222_X1 port map( A1 => A_shifted(40), A2 => n169, B1 => 
                           zeroSignal(40), B2 => n161, C1 => A_neg_shifted(40),
                           C2 => n147, ZN => n243);
   U198 : AOI222_X1 port map( A1 => A_shifted(38), A2 => n169, B1 => 
                           zeroSignal(38), B2 => n161, C1 => A_neg_shifted(38),
                           C2 => n147, ZN => n237);
   U199 : AOI222_X1 port map( A1 => A_shifted(37), A2 => n169, B1 => 
                           zeroSignal(37), B2 => n161, C1 => A_neg_shifted(37),
                           C2 => n147, ZN => n235);
   U200 : AOI222_X1 port map( A1 => A_shifted(36), A2 => n168, B1 => 
                           zeroSignal(36), B2 => n161, C1 => A_neg_shifted(36),
                           C2 => n147, ZN => n233);
   U201 : AOI222_X1 port map( A1 => A_shifted(35), A2 => n169, B1 => 
                           zeroSignal(35), B2 => n161, C1 => A_neg_shifted(35),
                           C2 => n147, ZN => n231);
   U202 : AOI22_X1 port map( A1 => A_neg(2), A2 => n302, B1 => A_signal(2), B2 
                           => n301, ZN => n220);
   U203 : AOI22_X1 port map( A1 => A_neg(5), A2 => n157, B1 => A_signal(5), B2 
                           => n150, ZN => n286);
   U204 : AOI222_X1 port map( A1 => A_shifted(7), A2 => n170, B1 => 
                           zeroSignal(7), B2 => n164, C1 => A_neg_shifted(7), 
                           C2 => n149, ZN => n297);
   U205 : AOI22_X1 port map( A1 => A_neg(6), A2 => n157, B1 => A_signal(6), B2 
                           => n150, ZN => n296);
   U206 : AOI22_X1 port map( A1 => A_neg(4), A2 => n158, B1 => A_signal(4), B2 
                           => n151, ZN => n264);
   U207 : NAND2_X1 port map( A1 => n264, A2 => n263, ZN => Y(4));
   U208 : AOI222_X1 port map( A1 => A_shifted(39), A2 => n168, B1 => 
                           zeroSignal(39), B2 => n161, C1 => A_neg_shifted(39),
                           C2 => n147, ZN => n239);
   U209 : NAND2_X1 port map( A1 => n240, A2 => n239, ZN => Y(39));
   U210 : AOI22_X1 port map( A1 => A_neg(3), A2 => n302, B1 => A_signal(3), B2 
                           => n153, ZN => n242);
   U211 : AOI222_X1 port map( A1 => A_shifted(48), A2 => n168, B1 => 
                           zeroSignal(48), B2 => n162, C1 => A_neg_shifted(48),
                           C2 => n147, ZN => n259);
   U212 : AOI22_X1 port map( A1 => A_neg(47), A2 => n156, B1 => A_signal(47), 
                           B2 => n150, ZN => n258);
   U213 : AOI222_X1 port map( A1 => A_shifted(45), A2 => n168, B1 => 
                           zeroSignal(45), B2 => n162, C1 => A_neg_shifted(45),
                           C2 => n147, ZN => n253);
   U214 : AOI22_X1 port map( A1 => A_neg(44), A2 => n156, B1 => A_signal(44), 
                           B2 => n150, ZN => n252);
   U215 : AOI222_X1 port map( A1 => A_shifted(32), A2 => n169, B1 => 
                           zeroSignal(32), B2 => n161, C1 => A_neg_shifted(32),
                           C2 => n147, ZN => n225);
   U216 : AOI22_X1 port map( A1 => A_neg(31), A2 => n154, B1 => A_signal(31), 
                           B2 => n151, ZN => n224);
   U217 : AOI222_X1 port map( A1 => A_shifted(42), A2 => n169, B1 => 
                           zeroSignal(42), B2 => n162, C1 => A_neg_shifted(42),
                           C2 => n147, ZN => n247);
   U218 : AOI22_X1 port map( A1 => A_neg(41), A2 => n154, B1 => A_signal(41), 
                           B2 => n150, ZN => n246);
   U219 : AOI222_X1 port map( A1 => A_shifted(21), A2 => n169, B1 => 
                           zeroSignal(21), B2 => n160, C1 => A_neg_shifted(21),
                           C2 => n147, ZN => n201);
   U220 : AOI22_X1 port map( A1 => A_neg(20), A2 => n154, B1 => A_signal(20), 
                           B2 => n150, ZN => n200);
   U221 : AOI21_X1 port map( B1 => n143, B2 => n142, A => Sel(2), ZN => n174);
   U222 : NOR3_X1 port map( A1 => n152, A2 => Sel(2), A3 => n308, ZN => n302);
   U223 : CLKBUF_X1 port map( A => n173, Z => n168);
   U224 : BUF_X1 port map( A => n301, Z => n153);
   U225 : INV_X1 port map( A => Sel(1), ZN => n308);
   U226 : INV_X1 port map( A => n143, ZN => n152);
   U227 : AOI222_X1 port map( A1 => A_shifted(3), A2 => n145, B1 => 
                           zeroSignal(3), B2 => n161, C1 => A_neg_shifted(3), 
                           C2 => n303, ZN => n241);
   U228 : INV_X1 port map( A => Sel(0), ZN => n307);
   U229 : NAND2_X1 port map( A1 => n220, A2 => n219, ZN => Y(2));
   U230 : NAND2_X1 port map( A1 => n242, A2 => n241, ZN => Y(3));
   U231 : AOI22_X1 port map( A1 => A_neg(7), A2 => n157, B1 => A_signal(7), B2 
                           => n151, ZN => n298);
   U232 : AOI222_X1 port map( A1 => A_shifted(8), A2 => n171, B1 => 
                           zeroSignal(8), B2 => n164, C1 => A_neg_shifted(8), 
                           C2 => n148, ZN => n299);

end SYN_BEHAVIORAL_2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity MUX51_MuxNbit64_14 is

   port( zeroSignal, A_signal, A_neg, A_shifted, A_neg_shifted : in 
         std_logic_vector (63 downto 0);  Sel : in std_logic_vector (2 downto 
         0);  Y : out std_logic_vector (63 downto 0));

end MUX51_MuxNbit64_14;

architecture SYN_BEHAVIORAL_2 of MUX51_MuxNbit64_14 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X3
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, 
      n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, 
      n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, 
      n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, 
      n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, 
      n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, 
      n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, 
      n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, 
      n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, 
      n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, 
      n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, 
      n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, 
      n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, 
      n296, n297, n298, n299, n300, n301, n302, n303, n304, n305 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n178, A2 => n177, ZN => Y(12));
   U2 : NAND2_X1 port map( A1 => n250, A2 => n249, ZN => Y(45));
   U3 : NAND2_X1 port map( A1 => n268, A2 => n267, ZN => Y(53));
   U4 : OR3_X1 port map( A1 => Sel(1), A2 => Sel(2), A3 => n304, ZN => n141);
   U5 : BUF_X2 port map( A => n301, Z => n144);
   U6 : NAND2_X2 port map( A1 => n184, A2 => n183, ZN => Y(15));
   U7 : CLKBUF_X1 port map( A => n155, Z => n154);
   U8 : CLKBUF_X1 port map( A => n156, Z => n159);
   U9 : BUF_X1 port map( A => n169, Z => n168);
   U10 : BUF_X1 port map( A => n298, Z => n155);
   U11 : CLKBUF_X3 port map( A => n159, Z => n157);
   U12 : BUF_X1 port map( A => n154, Z => n147);
   U13 : CLKBUF_X1 port map( A => n153, Z => n152);
   U14 : BUF_X1 port map( A => n154, Z => n148);
   U15 : BUF_X1 port map( A => n154, Z => n149);
   U16 : BUF_X1 port map( A => n167, Z => n165);
   U17 : BUF_X1 port map( A => n168, Z => n162);
   U18 : BUF_X1 port map( A => n168, Z => n163);
   U19 : BUF_X1 port map( A => n167, Z => n164);
   U20 : BUF_X1 port map( A => n168, Z => n161);
   U21 : BUF_X1 port map( A => n167, Z => n166);
   U22 : CLKBUF_X1 port map( A => n299, Z => n156);
   U23 : BUF_X1 port map( A => n169, Z => n167);
   U24 : NOR3_X1 port map( A1 => Sel(0), A2 => Sel(2), A3 => n305, ZN => n298);
   U25 : INV_X4 port map( A => n141, ZN => n297);
   U26 : BUF_X1 port map( A => n300, Z => n169);
   U27 : NOR2_X1 port map( A1 => n157, A2 => n170, ZN => n300);
   U28 : AOI222_X1 port map( A1 => A_shifted(45), A2 => n144, B1 => 
                           zeroSignal(45), B2 => n164, C1 => A_neg_shifted(45),
                           C2 => n157, ZN => n249);
   U29 : AOI22_X1 port map( A1 => A_neg(45), A2 => n150, B1 => A_signal(45), B2
                           => n297, ZN => n250);
   U30 : NAND2_X1 port map( A1 => n290, A2 => n289, ZN => Y(63));
   U31 : AOI222_X1 port map( A1 => A_shifted(63), A2 => n144, B1 => 
                           zeroSignal(63), B2 => n165, C1 => A_neg_shifted(63),
                           C2 => n157, ZN => n289);
   U32 : AOI22_X1 port map( A1 => A_neg(63), A2 => n151, B1 => A_signal(63), B2
                           => n297, ZN => n290);
   U33 : AOI22_X1 port map( A1 => A_neg(53), A2 => n151, B1 => A_signal(53), B2
                           => n297, ZN => n268);
   U34 : NAND2_X1 port map( A1 => n236, A2 => n235, ZN => Y(39));
   U35 : AOI222_X1 port map( A1 => A_shifted(39), A2 => n144, B1 => 
                           zeroSignal(39), B2 => n163, C1 => A_neg_shifted(39),
                           C2 => n157, ZN => n235);
   U36 : AOI22_X1 port map( A1 => A_neg(39), A2 => n149, B1 => A_signal(39), B2
                           => n297, ZN => n236);
   U37 : NAND2_X1 port map( A1 => n240, A2 => n239, ZN => Y(40));
   U38 : AOI222_X1 port map( A1 => A_shifted(40), A2 => n145, B1 => 
                           zeroSignal(40), B2 => n163, C1 => A_neg_shifted(40),
                           C2 => n157, ZN => n239);
   U39 : AOI22_X1 port map( A1 => A_neg(40), A2 => n149, B1 => A_signal(40), B2
                           => n297, ZN => n240);
   U40 : NAND2_X1 port map( A1 => n242, A2 => n241, ZN => Y(41));
   U41 : AOI222_X1 port map( A1 => A_shifted(41), A2 => n146, B1 => 
                           zeroSignal(41), B2 => n163, C1 => A_neg_shifted(41),
                           C2 => n157, ZN => n241);
   U42 : AOI22_X1 port map( A1 => A_neg(41), A2 => n149, B1 => A_signal(41), B2
                           => n297, ZN => n242);
   U43 : NAND2_X1 port map( A1 => n180, A2 => n179, ZN => Y(13));
   U44 : NAND2_X1 port map( A1 => n244, A2 => n243, ZN => Y(42));
   U45 : AOI22_X1 port map( A1 => A_neg(42), A2 => n150, B1 => A_signal(42), B2
                           => n297, ZN => n244);
   U46 : AOI222_X1 port map( A1 => A_shifted(42), A2 => n144, B1 => 
                           zeroSignal(42), B2 => n164, C1 => A_neg_shifted(42),
                           C2 => n157, ZN => n243);
   U47 : NAND2_X1 port map( A1 => n188, A2 => n187, ZN => Y(17));
   U48 : AOI22_X1 port map( A1 => A_neg(17), A2 => n147, B1 => A_signal(17), B2
                           => n297, ZN => n188);
   U49 : NAND2_X1 port map( A1 => n182, A2 => n181, ZN => Y(14));
   U50 : NAND2_X1 port map( A1 => n192, A2 => n191, ZN => Y(19));
   U51 : AOI222_X1 port map( A1 => A_shifted(19), A2 => n145, B1 => 
                           zeroSignal(19), B2 => n161, C1 => A_neg_shifted(19),
                           C2 => n158, ZN => n191);
   U52 : AOI22_X1 port map( A1 => A_neg(19), A2 => n147, B1 => A_signal(19), B2
                           => n297, ZN => n192);
   U53 : NAND2_X1 port map( A1 => n190, A2 => n189, ZN => Y(18));
   U54 : AOI222_X1 port map( A1 => A_shifted(18), A2 => n144, B1 => 
                           zeroSignal(18), B2 => n161, C1 => A_neg_shifted(18),
                           C2 => n158, ZN => n189);
   U55 : AOI22_X1 port map( A1 => A_neg(18), A2 => n147, B1 => A_signal(18), B2
                           => n297, ZN => n190);
   U56 : NAND2_X1 port map( A1 => n272, A2 => n271, ZN => Y(55));
   U57 : AOI222_X1 port map( A1 => A_shifted(55), A2 => n145, B1 => 
                           zeroSignal(55), B2 => n165, C1 => A_neg_shifted(55),
                           C2 => n157, ZN => n271);
   U58 : AOI22_X1 port map( A1 => A_neg(55), A2 => n151, B1 => A_signal(55), B2
                           => n297, ZN => n272);
   U59 : NAND2_X1 port map( A1 => n186, A2 => n185, ZN => Y(16));
   U60 : NAND2_X1 port map( A1 => n274, A2 => n273, ZN => Y(56));
   U61 : AOI222_X1 port map( A1 => A_shifted(56), A2 => n146, B1 => 
                           zeroSignal(56), B2 => n165, C1 => A_neg_shifted(56),
                           C2 => n157, ZN => n273);
   U62 : AOI22_X1 port map( A1 => A_neg(56), A2 => n151, B1 => A_signal(56), B2
                           => n297, ZN => n274);
   U63 : NAND2_X1 port map( A1 => n196, A2 => n195, ZN => Y(20));
   U64 : AOI222_X1 port map( A1 => A_shifted(20), A2 => n146, B1 => 
                           zeroSignal(20), B2 => n162, C1 => A_neg_shifted(20),
                           C2 => n157, ZN => n195);
   U65 : AOI22_X1 port map( A1 => A_neg(20), A2 => n148, B1 => A_signal(20), B2
                           => n297, ZN => n196);
   U66 : NAND2_X1 port map( A1 => n276, A2 => n275, ZN => Y(57));
   U67 : AOI222_X1 port map( A1 => A_shifted(57), A2 => n144, B1 => 
                           zeroSignal(57), B2 => n165, C1 => A_neg_shifted(57),
                           C2 => n157, ZN => n275);
   U68 : AOI22_X1 port map( A1 => A_neg(57), A2 => n151, B1 => A_signal(57), B2
                           => n297, ZN => n276);
   U69 : NAND2_X1 port map( A1 => n198, A2 => n197, ZN => Y(21));
   U70 : AOI222_X1 port map( A1 => A_shifted(21), A2 => n144, B1 => 
                           zeroSignal(21), B2 => n162, C1 => A_neg_shifted(21),
                           C2 => n157, ZN => n197);
   U71 : AOI22_X1 port map( A1 => A_neg(21), A2 => n148, B1 => A_signal(21), B2
                           => n297, ZN => n198);
   U72 : NAND2_X1 port map( A1 => n278, A2 => n277, ZN => Y(58));
   U73 : AOI222_X1 port map( A1 => A_shifted(58), A2 => n145, B1 => 
                           zeroSignal(58), B2 => n165, C1 => A_neg_shifted(58),
                           C2 => n157, ZN => n277);
   U74 : AOI22_X1 port map( A1 => A_neg(58), A2 => n151, B1 => A_signal(58), B2
                           => n297, ZN => n278);
   U75 : NAND2_X1 port map( A1 => n254, A2 => n253, ZN => Y(47));
   U76 : AOI22_X1 port map( A1 => A_neg(47), A2 => n150, B1 => A_signal(47), B2
                           => n297, ZN => n254);
   U77 : NAND2_X1 port map( A1 => n280, A2 => n279, ZN => Y(59));
   U78 : AOI222_X1 port map( A1 => A_shifted(59), A2 => n146, B1 => 
                           zeroSignal(59), B2 => n165, C1 => A_neg_shifted(59),
                           C2 => n157, ZN => n279);
   U79 : AOI22_X1 port map( A1 => A_neg(59), A2 => n151, B1 => A_signal(59), B2
                           => n297, ZN => n280);
   U80 : NAND2_X1 port map( A1 => n202, A2 => n201, ZN => Y(23));
   U81 : AOI22_X1 port map( A1 => A_neg(23), A2 => n148, B1 => A_signal(23), B2
                           => n297, ZN => n202);
   U82 : NAND2_X1 port map( A1 => n258, A2 => n257, ZN => Y(49));
   U83 : AOI222_X1 port map( A1 => A_shifted(49), A2 => n145, B1 => 
                           zeroSignal(49), B2 => n164, C1 => A_neg_shifted(49),
                           C2 => n157, ZN => n257);
   U84 : NAND2_X1 port map( A1 => n284, A2 => n283, ZN => Y(60));
   U85 : AOI222_X1 port map( A1 => A_shifted(60), A2 => n144, B1 => 
                           zeroSignal(60), B2 => n165, C1 => A_neg_shifted(60),
                           C2 => n157, ZN => n283);
   U86 : AOI22_X1 port map( A1 => A_neg(60), A2 => n151, B1 => A_signal(60), B2
                           => n297, ZN => n284);
   U87 : NAND2_X1 port map( A1 => n204, A2 => n203, ZN => Y(24));
   U88 : AOI222_X1 port map( A1 => A_shifted(24), A2 => n144, B1 => 
                           zeroSignal(24), B2 => n162, C1 => A_neg_shifted(24),
                           C2 => n157, ZN => n203);
   U89 : AOI22_X1 port map( A1 => A_neg(24), A2 => n148, B1 => A_signal(24), B2
                           => n297, ZN => n204);
   U90 : NAND2_X1 port map( A1 => n288, A2 => n287, ZN => Y(62));
   U91 : AOI222_X1 port map( A1 => A_shifted(62), A2 => n145, B1 => 
                           zeroSignal(62), B2 => n165, C1 => A_neg_shifted(62),
                           C2 => n157, ZN => n287);
   U92 : AOI22_X1 port map( A1 => A_neg(62), A2 => n151, B1 => A_signal(62), B2
                           => n297, ZN => n288);
   U93 : NAND2_X1 port map( A1 => n252, A2 => n251, ZN => Y(46));
   U94 : AOI222_X1 port map( A1 => A_shifted(46), A2 => n145, B1 => 
                           zeroSignal(46), B2 => n164, C1 => A_neg_shifted(46),
                           C2 => n157, ZN => n251);
   U95 : NAND2_X1 port map( A1 => n256, A2 => n255, ZN => Y(48));
   U96 : AOI222_X1 port map( A1 => A_shifted(48), A2 => n144, B1 => 
                           zeroSignal(48), B2 => n164, C1 => A_neg_shifted(48),
                           C2 => n157, ZN => n255);
   U97 : AOI22_X1 port map( A1 => A_neg(48), A2 => n150, B1 => A_signal(48), B2
                           => n297, ZN => n256);
   U98 : NAND2_X1 port map( A1 => n286, A2 => n285, ZN => Y(61));
   U99 : AOI222_X1 port map( A1 => A_shifted(61), A2 => n145, B1 => 
                           zeroSignal(61), B2 => n165, C1 => A_neg_shifted(61),
                           C2 => n157, ZN => n285);
   U100 : AOI22_X1 port map( A1 => A_neg(61), A2 => n151, B1 => A_signal(61), 
                           B2 => n297, ZN => n286);
   U101 : NAND2_X1 port map( A1 => n206, A2 => n205, ZN => Y(25));
   U102 : AOI222_X1 port map( A1 => A_shifted(25), A2 => n145, B1 => 
                           zeroSignal(25), B2 => n162, C1 => A_neg_shifted(25),
                           C2 => n157, ZN => n205);
   U103 : AOI22_X1 port map( A1 => A_neg(25), A2 => n148, B1 => A_signal(25), 
                           B2 => n297, ZN => n206);
   U104 : NAND2_X1 port map( A1 => n200, A2 => n199, ZN => Y(22));
   U105 : AOI222_X1 port map( A1 => A_shifted(22), A2 => n145, B1 => 
                           zeroSignal(22), B2 => n162, C1 => A_neg_shifted(22),
                           C2 => n157, ZN => n199);
   U106 : NAND2_X1 port map( A1 => n210, A2 => n209, ZN => Y(27));
   U107 : AOI222_X1 port map( A1 => A_shifted(27), A2 => n144, B1 => 
                           zeroSignal(27), B2 => n162, C1 => A_neg_shifted(27),
                           C2 => n157, ZN => n209);
   U108 : AOI22_X1 port map( A1 => A_neg(27), A2 => n148, B1 => A_signal(27), 
                           B2 => n297, ZN => n210);
   U109 : NAND2_X1 port map( A1 => n208, A2 => n207, ZN => Y(26));
   U110 : AOI222_X1 port map( A1 => A_shifted(26), A2 => n146, B1 => 
                           zeroSignal(26), B2 => n162, C1 => A_neg_shifted(26),
                           C2 => n157, ZN => n207);
   U111 : AOI22_X1 port map( A1 => A_neg(26), A2 => n148, B1 => A_signal(26), 
                           B2 => n297, ZN => n208);
   U112 : NAND2_X1 port map( A1 => n214, A2 => n213, ZN => Y(29));
   U113 : AOI222_X1 port map( A1 => A_shifted(29), A2 => n146, B1 => 
                           zeroSignal(29), B2 => n162, C1 => A_neg_shifted(29),
                           C2 => n157, ZN => n213);
   U114 : AOI22_X1 port map( A1 => A_neg(29), A2 => n148, B1 => A_signal(29), 
                           B2 => n297, ZN => n214);
   U115 : NAND2_X1 port map( A1 => n212, A2 => n211, ZN => Y(28));
   U116 : AOI222_X1 port map( A1 => A_shifted(28), A2 => n145, B1 => 
                           zeroSignal(28), B2 => n162, C1 => A_neg_shifted(28),
                           C2 => n157, ZN => n211);
   U117 : AOI22_X1 port map( A1 => A_neg(28), A2 => n148, B1 => A_signal(28), 
                           B2 => n297, ZN => n212);
   U118 : NAND2_X1 port map( A1 => n218, A2 => n217, ZN => Y(30));
   U119 : AOI222_X1 port map( A1 => A_shifted(30), A2 => n144, B1 => 
                           zeroSignal(30), B2 => n162, C1 => A_neg_shifted(30),
                           C2 => n157, ZN => n217);
   U120 : AOI22_X1 port map( A1 => A_neg(30), A2 => n148, B1 => A_signal(30), 
                           B2 => n297, ZN => n218);
   U121 : NAND2_X1 port map( A1 => n220, A2 => n219, ZN => Y(31));
   U122 : AOI222_X1 port map( A1 => A_shifted(31), A2 => n145, B1 => 
                           zeroSignal(31), B2 => n163, C1 => A_neg_shifted(31),
                           C2 => n157, ZN => n219);
   U123 : AOI22_X1 port map( A1 => A_neg(31), A2 => n149, B1 => A_signal(31), 
                           B2 => n297, ZN => n220);
   U124 : NAND2_X1 port map( A1 => n222, A2 => n221, ZN => Y(32));
   U125 : AOI222_X1 port map( A1 => A_shifted(32), A2 => n146, B1 => 
                           zeroSignal(32), B2 => n163, C1 => A_neg_shifted(32),
                           C2 => n157, ZN => n221);
   U126 : AOI22_X1 port map( A1 => A_neg(32), A2 => n149, B1 => A_signal(32), 
                           B2 => n297, ZN => n222);
   U127 : NAND2_X1 port map( A1 => n226, A2 => n225, ZN => Y(34));
   U128 : AOI22_X1 port map( A1 => A_neg(34), A2 => n149, B1 => A_signal(34), 
                           B2 => n297, ZN => n226);
   U129 : NAND2_X1 port map( A1 => n262, A2 => n261, ZN => Y(50));
   U130 : AOI22_X1 port map( A1 => A_neg(50), A2 => n150, B1 => A_signal(50), 
                           B2 => n297, ZN => n262);
   U131 : NAND2_X1 port map( A1 => n264, A2 => n263, ZN => Y(51));
   U132 : AOI222_X1 port map( A1 => A_shifted(51), A2 => n144, B1 => 
                           zeroSignal(51), B2 => n164, C1 => A_neg_shifted(51),
                           C2 => n157, ZN => n263);
   U133 : AOI22_X1 port map( A1 => A_neg(51), A2 => n150, B1 => A_signal(51), 
                           B2 => n297, ZN => n264);
   U134 : NAND2_X1 port map( A1 => n228, A2 => n227, ZN => Y(35));
   U135 : AOI222_X1 port map( A1 => A_shifted(35), A2 => n146, B1 => 
                           zeroSignal(35), B2 => n163, C1 => A_neg_shifted(35),
                           C2 => n157, ZN => n227);
   U136 : AOI22_X1 port map( A1 => A_neg(35), A2 => n149, B1 => A_signal(35), 
                           B2 => n297, ZN => n228);
   U137 : NAND2_X1 port map( A1 => n230, A2 => n229, ZN => Y(36));
   U138 : AOI222_X1 port map( A1 => A_shifted(36), A2 => n144, B1 => 
                           zeroSignal(36), B2 => n163, C1 => A_neg_shifted(36),
                           C2 => n157, ZN => n229);
   U139 : AOI22_X1 port map( A1 => A_neg(36), A2 => n149, B1 => A_signal(36), 
                           B2 => n297, ZN => n230);
   U140 : NAND2_X1 port map( A1 => n246, A2 => n245, ZN => Y(43));
   U141 : AOI222_X1 port map( A1 => A_shifted(43), A2 => n145, B1 => 
                           zeroSignal(43), B2 => n164, C1 => A_neg_shifted(43),
                           C2 => n157, ZN => n245);
   U142 : NAND2_X1 port map( A1 => n266, A2 => n265, ZN => Y(52));
   U143 : AOI222_X1 port map( A1 => A_shifted(52), A2 => n145, B1 => 
                           zeroSignal(52), B2 => n164, C1 => A_neg_shifted(52),
                           C2 => n157, ZN => n265);
   U144 : AOI22_X1 port map( A1 => A_neg(52), A2 => n150, B1 => A_signal(52), 
                           B2 => n297, ZN => n266);
   U145 : NAND2_X1 port map( A1 => n232, A2 => n231, ZN => Y(37));
   U146 : AOI222_X1 port map( A1 => A_shifted(37), A2 => n145, B1 => 
                           zeroSignal(37), B2 => n163, C1 => A_neg_shifted(37),
                           C2 => n157, ZN => n231);
   U147 : AOI22_X1 port map( A1 => A_neg(37), A2 => n149, B1 => A_signal(37), 
                           B2 => n297, ZN => n232);
   U148 : NAND2_X1 port map( A1 => n224, A2 => n223, ZN => Y(33));
   U149 : AOI222_X1 port map( A1 => A_shifted(33), A2 => n144, B1 => 
                           zeroSignal(33), B2 => n163, C1 => A_neg_shifted(33),
                           C2 => n157, ZN => n223);
   U150 : NAND2_X1 port map( A1 => n270, A2 => n269, ZN => Y(54));
   U151 : AOI222_X1 port map( A1 => A_shifted(54), A2 => n144, B1 => 
                           zeroSignal(54), B2 => n165, C1 => A_neg_shifted(54),
                           C2 => n157, ZN => n269);
   U152 : AOI22_X1 port map( A1 => A_neg(54), A2 => n151, B1 => A_signal(54), 
                           B2 => n297, ZN => n270);
   U153 : NAND2_X1 port map( A1 => n234, A2 => n233, ZN => Y(38));
   U154 : AOI222_X1 port map( A1 => A_shifted(38), A2 => n146, B1 => 
                           zeroSignal(38), B2 => n163, C1 => A_neg_shifted(38),
                           C2 => n157, ZN => n233);
   U155 : AOI22_X1 port map( A1 => A_neg(38), A2 => n149, B1 => A_signal(38), 
                           B2 => n297, ZN => n234);
   U156 : NAND2_X1 port map( A1 => n248, A2 => n247, ZN => Y(44));
   U157 : AOI22_X1 port map( A1 => A_neg(44), A2 => n150, B1 => A_signal(44), 
                           B2 => n297, ZN => n248);
   U158 : NAND2_X1 port map( A1 => n172, A2 => n171, ZN => Y(0));
   U159 : AOI22_X1 port map( A1 => A_neg(0), A2 => n147, B1 => A_signal(0), B2 
                           => n297, ZN => n172);
   U160 : AOI222_X1 port map( A1 => A_shifted(0), A2 => n146, B1 => 
                           zeroSignal(0), B2 => n161, C1 => A_neg_shifted(0), 
                           C2 => n157, ZN => n171);
   U161 : NAND2_X1 port map( A1 => n194, A2 => n193, ZN => Y(1));
   U162 : AOI22_X1 port map( A1 => A_neg(1), A2 => n147, B1 => A_signal(1), B2 
                           => n297, ZN => n194);
   U163 : AOI222_X1 port map( A1 => A_shifted(1), A2 => n145, B1 => 
                           zeroSignal(1), B2 => n161, C1 => A_neg_shifted(1), 
                           C2 => n157, ZN => n193);
   U164 : NAND2_X1 port map( A1 => n216, A2 => n215, ZN => Y(2));
   U165 : AOI22_X1 port map( A1 => A_neg(2), A2 => n148, B1 => A_signal(2), B2 
                           => n297, ZN => n216);
   U166 : AOI222_X1 port map( A1 => A_shifted(2), A2 => n144, B1 => 
                           zeroSignal(2), B2 => n162, C1 => A_neg_shifted(2), 
                           C2 => n157, ZN => n215);
   U167 : NAND2_X1 port map( A1 => n238, A2 => n237, ZN => Y(3));
   U168 : AOI22_X1 port map( A1 => A_neg(3), A2 => n149, B1 => A_signal(3), B2 
                           => n297, ZN => n238);
   U169 : AOI222_X1 port map( A1 => A_shifted(3), A2 => n144, B1 => 
                           zeroSignal(3), B2 => n163, C1 => A_neg_shifted(3), 
                           C2 => n157, ZN => n237);
   U170 : CLKBUF_X1 port map( A => n156, Z => n160);
   U171 : CLKBUF_X1 port map( A => n159, Z => n158);
   U172 : AOI222_X1 port map( A1 => A_shifted(15), A2 => n144, B1 => 
                           zeroSignal(15), B2 => n161, C1 => A_neg_shifted(15),
                           C2 => n160, ZN => n183);
   U173 : AOI22_X1 port map( A1 => A_neg(14), A2 => n147, B1 => A_signal(14), 
                           B2 => n297, ZN => n182);
   U174 : AOI222_X1 port map( A1 => A_shifted(7), A2 => n145, B1 => 
                           zeroSignal(7), B2 => n166, C1 => A_neg_shifted(7), 
                           C2 => n156, ZN => n293);
   U175 : AOI222_X1 port map( A1 => A_shifted(17), A2 => n146, B1 => 
                           zeroSignal(17), B2 => n161, C1 => A_neg_shifted(17),
                           C2 => n158, ZN => n187);
   U176 : AOI22_X1 port map( A1 => A_neg(16), A2 => n147, B1 => A_signal(16), 
                           B2 => n297, ZN => n186);
   U177 : AOI222_X1 port map( A1 => A_shifted(53), A2 => n146, B1 => 
                           zeroSignal(53), B2 => n165, C1 => A_neg_shifted(53),
                           C2 => n157, ZN => n267);
   U178 : NAND2_X1 port map( A1 => n176, A2 => n175, ZN => Y(11));
   U179 : AOI222_X1 port map( A1 => A_shifted(16), A2 => n145, B1 => 
                           zeroSignal(16), B2 => n161, C1 => A_neg_shifted(16),
                           C2 => n158, ZN => n185);
   U180 : AOI22_X1 port map( A1 => A_neg(15), A2 => n147, B1 => A_signal(15), 
                           B2 => n297, ZN => n184);
   U181 : NAND2_X1 port map( A1 => n174, A2 => n173, ZN => Y(10));
   U182 : NAND2_X1 port map( A1 => n303, A2 => n302, ZN => Y(9));
   U183 : AOI222_X1 port map( A1 => A_shifted(13), A2 => n145, B1 => 
                           zeroSignal(13), B2 => n161, C1 => A_neg_shifted(13),
                           C2 => n159, ZN => n179);
   U184 : AOI22_X1 port map( A1 => A_neg(12), A2 => n147, B1 => A_signal(12), 
                           B2 => n297, ZN => n178);
   U185 : AOI222_X1 port map( A1 => A_shifted(14), A2 => n146, B1 => 
                           zeroSignal(14), B2 => n161, C1 => A_neg_shifted(14),
                           C2 => n159, ZN => n181);
   U186 : AOI22_X1 port map( A1 => A_neg(13), A2 => n147, B1 => A_signal(13), 
                           B2 => n297, ZN => n180);
   U187 : AOI222_X1 port map( A1 => A_shifted(12), A2 => n144, B1 => 
                           zeroSignal(12), B2 => n161, C1 => A_neg_shifted(12),
                           C2 => n159, ZN => n177);
   U188 : AOI22_X1 port map( A1 => A_neg(11), A2 => n147, B1 => A_signal(11), 
                           B2 => n297, ZN => n176);
   U189 : AOI222_X1 port map( A1 => A_shifted(11), A2 => n146, B1 => 
                           zeroSignal(11), B2 => n161, C1 => A_neg_shifted(11),
                           C2 => n160, ZN => n175);
   U190 : AOI22_X1 port map( A1 => A_neg(10), A2 => n147, B1 => A_signal(10), 
                           B2 => n297, ZN => n174);
   U191 : NAND2_X1 port map( A1 => n296, A2 => n295, ZN => Y(8));
   U192 : NAND2_X1 port map( A1 => n294, A2 => n293, ZN => Y(7));
   U193 : AOI222_X1 port map( A1 => A_shifted(10), A2 => n145, B1 => 
                           zeroSignal(10), B2 => n161, C1 => A_neg_shifted(10),
                           C2 => n156, ZN => n173);
   U194 : AOI222_X1 port map( A1 => A_shifted(8), A2 => n146, B1 => 
                           zeroSignal(8), B2 => n166, C1 => A_neg_shifted(8), 
                           C2 => n156, ZN => n295);
   U195 : AOI22_X1 port map( A1 => A_neg(7), A2 => n152, B1 => A_signal(7), B2 
                           => n297, ZN => n294);
   U196 : AOI222_X1 port map( A1 => A_shifted(9), A2 => n144, B1 => 
                           zeroSignal(9), B2 => n166, C1 => A_neg_shifted(9), 
                           C2 => n156, ZN => n302);
   U197 : AOI22_X1 port map( A1 => A_neg(8), A2 => n152, B1 => A_signal(8), B2 
                           => n297, ZN => n296);
   U198 : CLKBUF_X1 port map( A => n153, Z => n151);
   U199 : BUF_X1 port map( A => n155, Z => n153);
   U200 : AOI222_X1 port map( A1 => A_shifted(6), A2 => n144, B1 => 
                           zeroSignal(6), B2 => n166, C1 => A_neg_shifted(6), 
                           C2 => n299, ZN => n291);
   U201 : AOI22_X1 port map( A1 => A_neg(6), A2 => n152, B1 => A_signal(6), B2 
                           => n297, ZN => n292);
   U202 : NAND2_X1 port map( A1 => n292, A2 => n291, ZN => Y(6));
   U203 : AOI222_X1 port map( A1 => A_shifted(50), A2 => n146, B1 => 
                           zeroSignal(50), B2 => n164, C1 => A_neg_shifted(50),
                           C2 => n157, ZN => n261);
   U204 : AOI22_X1 port map( A1 => A_neg(49), A2 => n150, B1 => A_signal(49), 
                           B2 => n297, ZN => n258);
   U205 : AOI222_X1 port map( A1 => A_shifted(47), A2 => n146, B1 => 
                           zeroSignal(47), B2 => n164, C1 => A_neg_shifted(47),
                           C2 => n157, ZN => n253);
   U206 : AOI22_X1 port map( A1 => A_neg(46), A2 => n150, B1 => A_signal(46), 
                           B2 => n297, ZN => n252);
   U207 : AOI222_X1 port map( A1 => A_shifted(34), A2 => n145, B1 => 
                           zeroSignal(34), B2 => n163, C1 => A_neg_shifted(34),
                           C2 => n157, ZN => n225);
   U208 : AOI22_X1 port map( A1 => A_neg(33), A2 => n149, B1 => A_signal(33), 
                           B2 => n297, ZN => n224);
   U209 : AOI22_X1 port map( A1 => A_neg(4), A2 => n150, B1 => A_signal(4), B2 
                           => n297, ZN => n260);
   U210 : BUF_X1 port map( A => n153, Z => n150);
   U211 : AOI222_X1 port map( A1 => A_shifted(44), A2 => n146, B1 => 
                           zeroSignal(44), B2 => n164, C1 => A_neg_shifted(44),
                           C2 => n157, ZN => n247);
   U212 : AOI22_X1 port map( A1 => A_neg(43), A2 => n150, B1 => A_signal(43), 
                           B2 => n297, ZN => n246);
   U213 : BUF_X1 port map( A => n301, Z => n142);
   U214 : BUF_X1 port map( A => n301, Z => n143);
   U215 : BUF_X2 port map( A => n142, Z => n145);
   U216 : BUF_X2 port map( A => n143, Z => n146);
   U217 : NOR3_X1 port map( A1 => n304, A2 => Sel(2), A3 => n305, ZN => n301);
   U218 : AOI222_X1 port map( A1 => A_shifted(23), A2 => n146, B1 => 
                           zeroSignal(23), B2 => n162, C1 => A_neg_shifted(23),
                           C2 => n157, ZN => n201);
   U219 : AOI22_X1 port map( A1 => A_neg(22), A2 => n148, B1 => A_signal(22), 
                           B2 => n297, ZN => n200);
   U220 : INV_X1 port map( A => Sel(0), ZN => n304);
   U221 : AOI21_X1 port map( B1 => n304, B2 => n305, A => Sel(2), ZN => n170);
   U222 : AND3_X1 port map( A1 => n304, A2 => n305, A3 => Sel(2), ZN => n299);
   U223 : NAND2_X1 port map( A1 => n260, A2 => n259, ZN => Y(4));
   U224 : AOI222_X1 port map( A1 => A_shifted(4), A2 => n146, B1 => 
                           zeroSignal(4), B2 => n164, C1 => A_neg_shifted(4), 
                           C2 => n157, ZN => n259);
   U225 : AOI222_X1 port map( A1 => A_shifted(5), A2 => n146, B1 => 
                           zeroSignal(5), B2 => n165, C1 => A_neg_shifted(5), 
                           C2 => n299, ZN => n281);
   U226 : AOI22_X1 port map( A1 => A_neg(5), A2 => n151, B1 => A_signal(5), B2 
                           => n297, ZN => n282);
   U227 : INV_X1 port map( A => Sel(1), ZN => n305);
   U228 : NAND2_X1 port map( A1 => n282, A2 => n281, ZN => Y(5));
   U229 : AOI22_X1 port map( A1 => A_neg(9), A2 => n152, B1 => A_signal(9), B2 
                           => n297, ZN => n303);

end SYN_BEHAVIORAL_2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity MUX51_MuxNbit64_13 is

   port( zeroSignal, A_signal, A_neg, A_shifted, A_neg_shifted : in 
         std_logic_vector (63 downto 0);  Sel : in std_logic_vector (2 downto 
         0);  Y : out std_logic_vector (63 downto 0));

end MUX51_MuxNbit64_13;

architecture SYN_BEHAVIORAL_2 of MUX51_MuxNbit64_13 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, 
      n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, 
      n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, 
      n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, 
      n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, 
      n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, 
      n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, 
      n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, 
      n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, 
      n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, 
      n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, 
      n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, 
      n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, 
      n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, 
      n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319 : 
      std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => n167, Z => n161);
   U2 : CLKBUF_X1 port map( A => n141, Z => n166);
   U3 : BUF_X1 port map( A => n141, Z => n167);
   U4 : BUF_X1 port map( A => n185, Z => n183);
   U5 : BUF_X1 port map( A => n142, Z => n158);
   U6 : BUF_X1 port map( A => n151, Z => n149);
   U7 : BUF_X1 port map( A => n142, Z => n159);
   U8 : BUF_X1 port map( A => n185, Z => n184);
   U9 : BUF_X1 port map( A => n151, Z => n150);
   U10 : BUF_X1 port map( A => n176, Z => n175);
   U11 : BUF_X1 port map( A => n176, Z => n174);
   U12 : AND3_X1 port map( A1 => n318, A2 => n319, A3 => Sel(2), ZN => n141);
   U13 : BUF_X1 port map( A => n315, Z => n185);
   U14 : NOR3_X1 port map( A1 => Sel(0), A2 => Sel(2), A3 => n319, ZN => n142);
   U15 : BUF_X1 port map( A => n183, Z => n182);
   U16 : BUF_X1 port map( A => n158, Z => n157);
   U17 : BUF_X1 port map( A => n149, Z => n148);
   U18 : BUF_X1 port map( A => n167, Z => n160);
   U19 : BUF_X1 port map( A => n184, Z => n177);
   U20 : BUF_X1 port map( A => n159, Z => n152);
   U21 : BUF_X1 port map( A => n150, Z => n143);
   U22 : BUF_X1 port map( A => n166, Z => n165);
   U23 : BUF_X1 port map( A => n166, Z => n164);
   U24 : BUF_X1 port map( A => n184, Z => n178);
   U25 : BUF_X1 port map( A => n159, Z => n153);
   U26 : BUF_X1 port map( A => n150, Z => n144);
   U27 : BUF_X1 port map( A => n166, Z => n163);
   U28 : BUF_X1 port map( A => n184, Z => n179);
   U29 : BUF_X1 port map( A => n159, Z => n154);
   U30 : BUF_X1 port map( A => n150, Z => n145);
   U31 : BUF_X1 port map( A => n167, Z => n162);
   U32 : BUF_X1 port map( A => n183, Z => n180);
   U33 : BUF_X1 port map( A => n158, Z => n155);
   U34 : BUF_X1 port map( A => n149, Z => n146);
   U35 : BUF_X1 port map( A => n183, Z => n181);
   U36 : BUF_X1 port map( A => n158, Z => n156);
   U37 : BUF_X1 port map( A => n149, Z => n147);
   U38 : BUF_X1 port map( A => n175, Z => n169);
   U39 : BUF_X1 port map( A => n175, Z => n170);
   U40 : BUF_X1 port map( A => n174, Z => n172);
   U41 : BUF_X1 port map( A => n175, Z => n168);
   U42 : BUF_X1 port map( A => n174, Z => n171);
   U43 : BUF_X1 port map( A => n174, Z => n173);
   U44 : INV_X1 port map( A => Sel(1), ZN => n319);
   U45 : NOR3_X1 port map( A1 => n318, A2 => Sel(2), A3 => n319, ZN => n315);
   U46 : BUF_X1 port map( A => n313, Z => n151);
   U47 : NOR3_X1 port map( A1 => Sel(1), A2 => Sel(2), A3 => n318, ZN => n313);
   U48 : INV_X1 port map( A => Sel(0), ZN => n318);
   U49 : BUF_X1 port map( A => n314, Z => n176);
   U50 : NOR2_X1 port map( A1 => n165, A2 => n186, ZN => n314);
   U51 : AOI21_X1 port map( B1 => n318, B2 => n319, A => Sel(2), ZN => n186);
   U52 : NAND2_X1 port map( A1 => n310, A2 => n309, ZN => Y(7));
   U53 : AOI22_X1 port map( A1 => A_neg(7), A2 => n157, B1 => A_signal(7), B2 
                           => n148, ZN => n310);
   U54 : AOI222_X1 port map( A1 => A_shifted(6), A2 => n182, B1 => 
                           zeroSignal(6), B2 => n173, C1 => A_neg_shifted(6), 
                           C2 => n160, ZN => n307);
   U55 : NAND2_X1 port map( A1 => n312, A2 => n311, ZN => Y(8));
   U56 : AOI222_X1 port map( A1 => A_shifted(8), A2 => n182, B1 => 
                           zeroSignal(8), B2 => n173, C1 => A_neg_shifted(8), 
                           C2 => n160, ZN => n311);
   U57 : AOI222_X1 port map( A1 => A_shifted(9), A2 => n182, B1 => 
                           zeroSignal(9), B2 => n173, C1 => A_neg_shifted(9), 
                           C2 => n160, ZN => n316);
   U58 : AOI222_X1 port map( A1 => A_shifted(11), A2 => n177, B1 => 
                           zeroSignal(11), B2 => n168, C1 => A_neg_shifted(11),
                           C2 => n165, ZN => n191);
   U59 : NAND2_X1 port map( A1 => n212, A2 => n211, ZN => Y(20));
   U60 : AOI22_X1 port map( A1 => A_neg(20), A2 => n153, B1 => A_signal(20), B2
                           => n144, ZN => n212);
   U61 : AOI222_X1 port map( A1 => A_shifted(20), A2 => n178, B1 => 
                           zeroSignal(20), B2 => n169, C1 => A_neg_shifted(20),
                           C2 => n164, ZN => n211);
   U62 : NAND2_X1 port map( A1 => n216, A2 => n215, ZN => Y(22));
   U63 : AOI22_X1 port map( A1 => A_neg(22), A2 => n153, B1 => A_signal(22), B2
                           => n144, ZN => n216);
   U64 : AOI222_X1 port map( A1 => A_shifted(22), A2 => n178, B1 => 
                           zeroSignal(22), B2 => n169, C1 => A_neg_shifted(22),
                           C2 => n164, ZN => n215);
   U65 : NAND2_X1 port map( A1 => n214, A2 => n213, ZN => Y(21));
   U66 : AOI22_X1 port map( A1 => A_neg(21), A2 => n153, B1 => A_signal(21), B2
                           => n144, ZN => n214);
   U67 : AOI222_X1 port map( A1 => A_shifted(21), A2 => n178, B1 => 
                           zeroSignal(21), B2 => n169, C1 => A_neg_shifted(21),
                           C2 => n164, ZN => n213);
   U68 : NAND2_X1 port map( A1 => n218, A2 => n217, ZN => Y(23));
   U69 : AOI22_X1 port map( A1 => A_neg(23), A2 => n153, B1 => A_signal(23), B2
                           => n144, ZN => n218);
   U70 : AOI222_X1 port map( A1 => A_shifted(23), A2 => n178, B1 => 
                           zeroSignal(23), B2 => n169, C1 => A_neg_shifted(23),
                           C2 => n164, ZN => n217);
   U71 : NAND2_X1 port map( A1 => n220, A2 => n219, ZN => Y(24));
   U72 : AOI222_X1 port map( A1 => A_shifted(24), A2 => n178, B1 => 
                           zeroSignal(24), B2 => n169, C1 => A_neg_shifted(24),
                           C2 => n163, ZN => n219);
   U73 : NAND2_X1 port map( A1 => n224, A2 => n223, ZN => Y(26));
   U74 : AOI22_X1 port map( A1 => A_neg(26), A2 => n153, B1 => A_signal(26), B2
                           => n144, ZN => n224);
   U75 : AOI222_X1 port map( A1 => A_shifted(26), A2 => n178, B1 => 
                           zeroSignal(26), B2 => n169, C1 => A_neg_shifted(26),
                           C2 => n163, ZN => n223);
   U76 : NAND2_X1 port map( A1 => n228, A2 => n227, ZN => Y(28));
   U77 : AOI22_X1 port map( A1 => A_neg(28), A2 => n153, B1 => A_signal(28), B2
                           => n144, ZN => n228);
   U78 : AOI222_X1 port map( A1 => A_shifted(28), A2 => n178, B1 => 
                           zeroSignal(28), B2 => n169, C1 => A_neg_shifted(28),
                           C2 => n163, ZN => n227);
   U79 : NAND2_X1 port map( A1 => n226, A2 => n225, ZN => Y(27));
   U80 : AOI22_X1 port map( A1 => A_neg(27), A2 => n153, B1 => A_signal(27), B2
                           => n144, ZN => n226);
   U81 : AOI222_X1 port map( A1 => A_shifted(27), A2 => n178, B1 => 
                           zeroSignal(27), B2 => n169, C1 => A_neg_shifted(27),
                           C2 => n163, ZN => n225);
   U82 : NAND2_X1 port map( A1 => n230, A2 => n229, ZN => Y(29));
   U83 : AOI22_X1 port map( A1 => A_neg(29), A2 => n153, B1 => A_signal(29), B2
                           => n144, ZN => n230);
   U84 : AOI222_X1 port map( A1 => A_shifted(29), A2 => n178, B1 => 
                           zeroSignal(29), B2 => n169, C1 => A_neg_shifted(29),
                           C2 => n163, ZN => n229);
   U85 : NAND2_X1 port map( A1 => n234, A2 => n233, ZN => Y(30));
   U86 : AOI22_X1 port map( A1 => A_neg(30), A2 => n153, B1 => A_signal(30), B2
                           => n144, ZN => n234);
   U87 : AOI222_X1 port map( A1 => A_shifted(30), A2 => n179, B1 => 
                           zeroSignal(30), B2 => n169, C1 => A_neg_shifted(30),
                           C2 => n163, ZN => n233);
   U88 : NAND2_X1 port map( A1 => n236, A2 => n235, ZN => Y(31));
   U89 : AOI22_X1 port map( A1 => A_neg(31), A2 => n154, B1 => A_signal(31), B2
                           => n145, ZN => n236);
   U90 : AOI222_X1 port map( A1 => A_shifted(31), A2 => n179, B1 => 
                           zeroSignal(31), B2 => n170, C1 => A_neg_shifted(31),
                           C2 => n163, ZN => n235);
   U91 : NAND2_X1 port map( A1 => n238, A2 => n237, ZN => Y(32));
   U92 : AOI22_X1 port map( A1 => A_neg(32), A2 => n154, B1 => A_signal(32), B2
                           => n145, ZN => n238);
   U93 : AOI222_X1 port map( A1 => A_shifted(32), A2 => n179, B1 => 
                           zeroSignal(32), B2 => n170, C1 => A_neg_shifted(32),
                           C2 => n163, ZN => n237);
   U94 : NAND2_X1 port map( A1 => n242, A2 => n241, ZN => Y(34));
   U95 : AOI22_X1 port map( A1 => A_neg(34), A2 => n154, B1 => A_signal(34), B2
                           => n145, ZN => n242);
   U96 : AOI222_X1 port map( A1 => A_shifted(34), A2 => n179, B1 => 
                           zeroSignal(34), B2 => n170, C1 => A_neg_shifted(34),
                           C2 => n163, ZN => n241);
   U97 : NAND2_X1 port map( A1 => n240, A2 => n239, ZN => Y(33));
   U98 : AOI22_X1 port map( A1 => A_neg(33), A2 => n154, B1 => A_signal(33), B2
                           => n145, ZN => n240);
   U99 : AOI222_X1 port map( A1 => A_shifted(33), A2 => n179, B1 => 
                           zeroSignal(33), B2 => n170, C1 => A_neg_shifted(33),
                           C2 => n163, ZN => n239);
   U100 : NAND2_X1 port map( A1 => n252, A2 => n251, ZN => Y(39));
   U101 : AOI222_X1 port map( A1 => A_shifted(39), A2 => n179, B1 => 
                           zeroSignal(39), B2 => n170, C1 => A_neg_shifted(39),
                           C2 => n162, ZN => n251);
   U102 : AOI22_X1 port map( A1 => A_neg(39), A2 => n154, B1 => A_signal(39), 
                           B2 => n145, ZN => n252);
   U103 : NAND2_X1 port map( A1 => n244, A2 => n243, ZN => Y(35));
   U104 : AOI222_X1 port map( A1 => A_shifted(35), A2 => n179, B1 => 
                           zeroSignal(35), B2 => n170, C1 => A_neg_shifted(35),
                           C2 => n162, ZN => n243);
   U105 : NAND2_X1 port map( A1 => n198, A2 => n197, ZN => Y(14));
   U106 : AOI222_X1 port map( A1 => A_shifted(14), A2 => n177, B1 => 
                           zeroSignal(14), B2 => n168, C1 => A_neg_shifted(14),
                           C2 => n164, ZN => n197);
   U107 : NAND2_X1 port map( A1 => n248, A2 => n247, ZN => Y(37));
   U108 : AOI22_X1 port map( A1 => A_neg(37), A2 => n154, B1 => A_signal(37), 
                           B2 => n145, ZN => n248);
   U109 : AOI222_X1 port map( A1 => A_shifted(37), A2 => n179, B1 => 
                           zeroSignal(37), B2 => n170, C1 => A_neg_shifted(37),
                           C2 => n162, ZN => n247);
   U110 : NAND2_X1 port map( A1 => n250, A2 => n249, ZN => Y(38));
   U111 : AOI22_X1 port map( A1 => A_neg(38), A2 => n154, B1 => A_signal(38), 
                           B2 => n145, ZN => n250);
   U112 : AOI222_X1 port map( A1 => A_shifted(38), A2 => n179, B1 => 
                           zeroSignal(38), B2 => n170, C1 => A_neg_shifted(38),
                           C2 => n162, ZN => n249);
   U113 : NAND2_X1 port map( A1 => n204, A2 => n203, ZN => Y(17));
   U114 : AOI222_X1 port map( A1 => A_shifted(17), A2 => n177, B1 => 
                           zeroSignal(17), B2 => n168, C1 => A_neg_shifted(17),
                           C2 => n164, ZN => n203);
   U115 : NAND2_X1 port map( A1 => n256, A2 => n255, ZN => Y(40));
   U116 : AOI222_X1 port map( A1 => A_shifted(40), A2 => n180, B1 => 
                           zeroSignal(40), B2 => n170, C1 => A_neg_shifted(40),
                           C2 => n162, ZN => n255);
   U117 : AOI22_X1 port map( A1 => A_neg(40), A2 => n154, B1 => A_signal(40), 
                           B2 => n145, ZN => n256);
   U118 : NAND2_X1 port map( A1 => n208, A2 => n207, ZN => Y(19));
   U119 : AOI22_X1 port map( A1 => A_neg(19), A2 => n152, B1 => A_signal(19), 
                           B2 => n143, ZN => n208);
   U120 : AOI222_X1 port map( A1 => A_shifted(19), A2 => n177, B1 => 
                           zeroSignal(19), B2 => n168, C1 => A_neg_shifted(19),
                           C2 => n164, ZN => n207);
   U121 : NAND2_X1 port map( A1 => n258, A2 => n257, ZN => Y(41));
   U122 : AOI222_X1 port map( A1 => A_shifted(41), A2 => n180, B1 => 
                           zeroSignal(41), B2 => n170, C1 => A_neg_shifted(41),
                           C2 => n162, ZN => n257);
   U123 : AOI22_X1 port map( A1 => A_neg(41), A2 => n154, B1 => A_signal(41), 
                           B2 => n145, ZN => n258);
   U124 : NAND2_X1 port map( A1 => n200, A2 => n199, ZN => Y(15));
   U125 : AOI222_X1 port map( A1 => A_shifted(15), A2 => n177, B1 => 
                           zeroSignal(15), B2 => n168, C1 => A_neg_shifted(15),
                           C2 => n164, ZN => n199);
   U126 : NAND2_X1 port map( A1 => n260, A2 => n259, ZN => Y(42));
   U127 : AOI222_X1 port map( A1 => A_shifted(42), A2 => n180, B1 => 
                           zeroSignal(42), B2 => n171, C1 => A_neg_shifted(42),
                           C2 => n162, ZN => n259);
   U128 : AOI22_X1 port map( A1 => A_neg(42), A2 => n155, B1 => A_signal(42), 
                           B2 => n146, ZN => n260);
   U129 : NAND2_X1 port map( A1 => n262, A2 => n261, ZN => Y(43));
   U130 : AOI222_X1 port map( A1 => A_shifted(43), A2 => n180, B1 => 
                           zeroSignal(43), B2 => n171, C1 => A_neg_shifted(43),
                           C2 => n162, ZN => n261);
   U131 : AOI22_X1 port map( A1 => A_neg(43), A2 => n155, B1 => A_signal(43), 
                           B2 => n146, ZN => n262);
   U132 : NAND2_X1 port map( A1 => n202, A2 => n201, ZN => Y(16));
   U133 : AOI222_X1 port map( A1 => A_shifted(16), A2 => n177, B1 => 
                           zeroSignal(16), B2 => n168, C1 => A_neg_shifted(16),
                           C2 => n164, ZN => n201);
   U134 : NAND2_X1 port map( A1 => n206, A2 => n205, ZN => Y(18));
   U135 : AOI222_X1 port map( A1 => A_shifted(18), A2 => n177, B1 => 
                           zeroSignal(18), B2 => n168, C1 => A_neg_shifted(18),
                           C2 => n164, ZN => n205);
   U136 : NAND2_X1 port map( A1 => n264, A2 => n263, ZN => Y(44));
   U137 : AOI22_X1 port map( A1 => A_neg(44), A2 => n155, B1 => A_signal(44), 
                           B2 => n146, ZN => n264);
   U138 : AOI222_X1 port map( A1 => A_shifted(44), A2 => n180, B1 => 
                           zeroSignal(44), B2 => n171, C1 => A_neg_shifted(44),
                           C2 => n162, ZN => n263);
   U139 : NAND2_X1 port map( A1 => n222, A2 => n221, ZN => Y(25));
   U140 : AOI22_X1 port map( A1 => A_neg(25), A2 => n153, B1 => A_signal(25), 
                           B2 => n144, ZN => n222);
   U141 : AOI222_X1 port map( A1 => A_shifted(25), A2 => n178, B1 => 
                           zeroSignal(25), B2 => n169, C1 => A_neg_shifted(25),
                           C2 => n163, ZN => n221);
   U142 : NAND2_X1 port map( A1 => n270, A2 => n269, ZN => Y(47));
   U143 : AOI222_X1 port map( A1 => A_shifted(47), A2 => n180, B1 => 
                           zeroSignal(47), B2 => n171, C1 => A_neg_shifted(47),
                           C2 => n161, ZN => n269);
   U144 : AOI22_X1 port map( A1 => A_neg(47), A2 => n155, B1 => A_signal(47), 
                           B2 => n146, ZN => n270);
   U145 : NAND2_X1 port map( A1 => n292, A2 => n291, ZN => Y(57));
   U146 : AOI222_X1 port map( A1 => A_shifted(57), A2 => n181, B1 => 
                           zeroSignal(57), B2 => n172, C1 => A_neg_shifted(57),
                           C2 => n160, ZN => n291);
   U147 : AOI22_X1 port map( A1 => A_neg(57), A2 => n156, B1 => A_signal(57), 
                           B2 => n147, ZN => n292);
   U148 : NAND2_X1 port map( A1 => n304, A2 => n303, ZN => Y(62));
   U149 : AOI222_X1 port map( A1 => A_shifted(62), A2 => n182, B1 => 
                           zeroSignal(62), B2 => n172, C1 => A_neg_shifted(62),
                           C2 => n160, ZN => n303);
   U150 : AOI22_X1 port map( A1 => A_neg(62), A2 => n156, B1 => A_signal(62), 
                           B2 => n147, ZN => n304);
   U151 : NAND2_X1 port map( A1 => n294, A2 => n293, ZN => Y(58));
   U152 : AOI222_X1 port map( A1 => A_shifted(58), A2 => n181, B1 => 
                           zeroSignal(58), B2 => n172, C1 => A_neg_shifted(58),
                           C2 => n160, ZN => n293);
   U153 : AOI22_X1 port map( A1 => A_neg(58), A2 => n156, B1 => A_signal(58), 
                           B2 => n147, ZN => n294);
   U154 : NAND2_X1 port map( A1 => n306, A2 => n305, ZN => Y(63));
   U155 : AOI222_X1 port map( A1 => A_shifted(63), A2 => n182, B1 => 
                           zeroSignal(63), B2 => n172, C1 => A_neg_shifted(63),
                           C2 => n160, ZN => n305);
   U156 : AOI22_X1 port map( A1 => A_neg(63), A2 => n156, B1 => A_signal(63), 
                           B2 => n147, ZN => n306);
   U157 : NAND2_X1 port map( A1 => n296, A2 => n295, ZN => Y(59));
   U158 : AOI222_X1 port map( A1 => A_shifted(59), A2 => n181, B1 => 
                           zeroSignal(59), B2 => n172, C1 => A_neg_shifted(59),
                           C2 => n160, ZN => n295);
   U159 : AOI22_X1 port map( A1 => A_neg(59), A2 => n156, B1 => A_signal(59), 
                           B2 => n147, ZN => n296);
   U160 : NAND2_X1 port map( A1 => n302, A2 => n301, ZN => Y(61));
   U161 : AOI222_X1 port map( A1 => A_shifted(61), A2 => n182, B1 => 
                           zeroSignal(61), B2 => n172, C1 => A_neg_shifted(61),
                           C2 => n160, ZN => n301);
   U162 : AOI22_X1 port map( A1 => A_neg(61), A2 => n156, B1 => A_signal(61), 
                           B2 => n147, ZN => n302);
   U163 : NAND2_X1 port map( A1 => n300, A2 => n299, ZN => Y(60));
   U164 : AOI222_X1 port map( A1 => A_shifted(60), A2 => n182, B1 => 
                           zeroSignal(60), B2 => n172, C1 => A_neg_shifted(60),
                           C2 => n160, ZN => n299);
   U165 : AOI22_X1 port map( A1 => A_neg(60), A2 => n156, B1 => A_signal(60), 
                           B2 => n147, ZN => n300);
   U166 : NAND2_X1 port map( A1 => n274, A2 => n273, ZN => Y(49));
   U167 : AOI22_X1 port map( A1 => A_neg(49), A2 => n155, B1 => A_signal(49), 
                           B2 => n146, ZN => n274);
   U168 : NAND2_X1 port map( A1 => n280, A2 => n279, ZN => Y(51));
   U169 : AOI222_X1 port map( A1 => A_shifted(51), A2 => n181, B1 => 
                           zeroSignal(51), B2 => n171, C1 => A_neg_shifted(51),
                           C2 => n161, ZN => n279);
   U170 : NAND2_X1 port map( A1 => n246, A2 => n245, ZN => Y(36));
   U171 : AOI22_X1 port map( A1 => A_neg(36), A2 => n154, B1 => A_signal(36), 
                           B2 => n145, ZN => n246);
   U172 : AOI222_X1 port map( A1 => A_shifted(36), A2 => n179, B1 => 
                           zeroSignal(36), B2 => n170, C1 => A_neg_shifted(36),
                           C2 => n162, ZN => n245);
   U173 : NAND2_X1 port map( A1 => n278, A2 => n277, ZN => Y(50));
   U174 : AOI222_X1 port map( A1 => A_shifted(50), A2 => n181, B1 => 
                           zeroSignal(50), B2 => n171, C1 => A_neg_shifted(50),
                           C2 => n161, ZN => n277);
   U175 : AOI22_X1 port map( A1 => A_neg(50), A2 => n155, B1 => A_signal(50), 
                           B2 => n146, ZN => n278);
   U176 : NAND2_X1 port map( A1 => n272, A2 => n271, ZN => Y(48));
   U177 : AOI222_X1 port map( A1 => A_shifted(48), A2 => n180, B1 => 
                           zeroSignal(48), B2 => n171, C1 => A_neg_shifted(48),
                           C2 => n161, ZN => n271);
   U178 : NAND2_X1 port map( A1 => n282, A2 => n281, ZN => Y(52));
   U179 : AOI22_X1 port map( A1 => A_neg(52), A2 => n155, B1 => A_signal(52), 
                           B2 => n146, ZN => n282);
   U180 : NAND2_X1 port map( A1 => n284, A2 => n283, ZN => Y(53));
   U181 : AOI222_X1 port map( A1 => A_shifted(53), A2 => n181, B1 => 
                           zeroSignal(53), B2 => n172, C1 => A_neg_shifted(53),
                           C2 => n161, ZN => n283);
   U182 : AOI22_X1 port map( A1 => A_neg(53), A2 => n156, B1 => A_signal(53), 
                           B2 => n147, ZN => n284);
   U183 : NAND2_X1 port map( A1 => n266, A2 => n265, ZN => Y(45));
   U184 : AOI222_X1 port map( A1 => A_shifted(45), A2 => n180, B1 => 
                           zeroSignal(45), B2 => n171, C1 => A_neg_shifted(45),
                           C2 => n162, ZN => n265);
   U185 : NAND2_X1 port map( A1 => n286, A2 => n285, ZN => Y(54));
   U186 : AOI222_X1 port map( A1 => A_shifted(54), A2 => n181, B1 => 
                           zeroSignal(54), B2 => n172, C1 => A_neg_shifted(54),
                           C2 => n161, ZN => n285);
   U187 : AOI22_X1 port map( A1 => A_neg(54), A2 => n156, B1 => A_signal(54), 
                           B2 => n147, ZN => n286);
   U188 : NAND2_X1 port map( A1 => n288, A2 => n287, ZN => Y(55));
   U189 : AOI222_X1 port map( A1 => A_shifted(55), A2 => n181, B1 => 
                           zeroSignal(55), B2 => n172, C1 => A_neg_shifted(55),
                           C2 => n161, ZN => n287);
   U190 : AOI22_X1 port map( A1 => A_neg(55), A2 => n156, B1 => A_signal(55), 
                           B2 => n147, ZN => n288);
   U191 : NAND2_X1 port map( A1 => n290, A2 => n289, ZN => Y(56));
   U192 : AOI222_X1 port map( A1 => A_shifted(56), A2 => n181, B1 => 
                           zeroSignal(56), B2 => n172, C1 => A_neg_shifted(56),
                           C2 => n161, ZN => n289);
   U193 : AOI22_X1 port map( A1 => A_neg(56), A2 => n156, B1 => A_signal(56), 
                           B2 => n147, ZN => n290);
   U194 : NAND2_X1 port map( A1 => n268, A2 => n267, ZN => Y(46));
   U195 : AOI22_X1 port map( A1 => A_neg(46), A2 => n155, B1 => A_signal(46), 
                           B2 => n146, ZN => n268);
   U196 : NAND2_X1 port map( A1 => n188, A2 => n187, ZN => Y(0));
   U197 : AOI22_X1 port map( A1 => A_neg(0), A2 => n152, B1 => A_signal(0), B2 
                           => n143, ZN => n188);
   U198 : AOI222_X1 port map( A1 => A_shifted(0), A2 => n177, B1 => 
                           zeroSignal(0), B2 => n168, C1 => A_neg_shifted(0), 
                           C2 => n165, ZN => n187);
   U199 : NAND2_X1 port map( A1 => n210, A2 => n209, ZN => Y(1));
   U200 : AOI22_X1 port map( A1 => A_neg(1), A2 => n152, B1 => A_signal(1), B2 
                           => n143, ZN => n210);
   U201 : AOI222_X1 port map( A1 => A_shifted(1), A2 => n178, B1 => 
                           zeroSignal(1), B2 => n168, C1 => A_neg_shifted(1), 
                           C2 => n164, ZN => n209);
   U202 : NAND2_X1 port map( A1 => n232, A2 => n231, ZN => Y(2));
   U203 : AOI22_X1 port map( A1 => A_neg(2), A2 => n153, B1 => A_signal(2), B2 
                           => n144, ZN => n232);
   U204 : AOI222_X1 port map( A1 => A_shifted(2), A2 => n179, B1 => 
                           zeroSignal(2), B2 => n169, C1 => A_neg_shifted(2), 
                           C2 => n163, ZN => n231);
   U205 : NAND2_X1 port map( A1 => n254, A2 => n253, ZN => Y(3));
   U206 : AOI22_X1 port map( A1 => A_neg(3), A2 => n154, B1 => A_signal(3), B2 
                           => n145, ZN => n254);
   U207 : AOI222_X1 port map( A1 => A_shifted(3), A2 => n180, B1 => 
                           zeroSignal(3), B2 => n170, C1 => A_neg_shifted(3), 
                           C2 => n162, ZN => n253);
   U208 : NAND2_X1 port map( A1 => n276, A2 => n275, ZN => Y(4));
   U209 : AOI22_X1 port map( A1 => A_neg(4), A2 => n155, B1 => A_signal(4), B2 
                           => n146, ZN => n276);
   U210 : AOI222_X1 port map( A1 => A_shifted(4), A2 => n181, B1 => 
                           zeroSignal(4), B2 => n171, C1 => A_neg_shifted(4), 
                           C2 => n161, ZN => n275);
   U211 : NAND2_X1 port map( A1 => n298, A2 => n297, ZN => Y(5));
   U212 : AOI22_X1 port map( A1 => A_neg(5), A2 => n156, B1 => A_signal(5), B2 
                           => n147, ZN => n298);
   U213 : AOI222_X1 port map( A1 => A_shifted(5), A2 => n182, B1 => 
                           zeroSignal(5), B2 => n172, C1 => A_neg_shifted(5), 
                           C2 => n160, ZN => n297);
   U214 : AOI22_X1 port map( A1 => A_neg(16), A2 => n152, B1 => A_signal(16), 
                           B2 => n143, ZN => n202);
   U215 : AOI22_X1 port map( A1 => A_neg(8), A2 => n157, B1 => A_signal(8), B2 
                           => n148, ZN => n312);
   U216 : AOI22_X1 port map( A1 => A_neg(18), A2 => n152, B1 => A_signal(18), 
                           B2 => n143, ZN => n206);
   U217 : AOI222_X1 port map( A1 => A_shifted(7), A2 => n182, B1 => 
                           zeroSignal(7), B2 => n173, C1 => A_neg_shifted(7), 
                           C2 => n160, ZN => n309);
   U218 : NAND2_X1 port map( A1 => n308, A2 => n307, ZN => Y(6));
   U219 : AOI222_X1 port map( A1 => A_shifted(13), A2 => n177, B1 => 
                           zeroSignal(13), B2 => n168, C1 => A_neg_shifted(13),
                           C2 => n164, ZN => n195);
   U220 : NAND2_X1 port map( A1 => n196, A2 => n195, ZN => Y(13));
   U221 : AOI22_X1 port map( A1 => A_neg(17), A2 => n152, B1 => A_signal(17), 
                           B2 => n143, ZN => n204);
   U222 : AOI222_X1 port map( A1 => A_shifted(12), A2 => n177, B1 => 
                           zeroSignal(12), B2 => n168, C1 => A_neg_shifted(12),
                           C2 => n165, ZN => n193);
   U223 : NAND2_X1 port map( A1 => n192, A2 => n191, ZN => Y(11));
   U224 : NAND2_X1 port map( A1 => n194, A2 => n193, ZN => Y(12));
   U225 : AOI22_X1 port map( A1 => A_neg(14), A2 => n152, B1 => A_signal(14), 
                           B2 => n143, ZN => n198);
   U226 : AOI22_X1 port map( A1 => A_neg(15), A2 => n152, B1 => A_signal(15), 
                           B2 => n143, ZN => n200);
   U227 : AOI22_X1 port map( A1 => A_neg(13), A2 => n152, B1 => A_signal(13), 
                           B2 => n143, ZN => n196);
   U228 : AOI22_X1 port map( A1 => A_neg(12), A2 => n152, B1 => A_signal(12), 
                           B2 => n143, ZN => n194);
   U229 : AOI222_X1 port map( A1 => A_shifted(10), A2 => n177, B1 => 
                           zeroSignal(10), B2 => n168, C1 => A_neg_shifted(10),
                           C2 => n165, ZN => n189);
   U230 : NAND2_X1 port map( A1 => n317, A2 => n316, ZN => Y(9));
   U231 : NAND2_X1 port map( A1 => n190, A2 => n189, ZN => Y(10));
   U232 : AOI22_X1 port map( A1 => A_neg(11), A2 => n152, B1 => A_signal(11), 
                           B2 => n143, ZN => n192);
   U233 : AOI22_X1 port map( A1 => A_neg(6), A2 => n157, B1 => A_signal(6), B2 
                           => n148, ZN => n308);
   U234 : AOI22_X1 port map( A1 => A_neg(9), A2 => n157, B1 => A_signal(9), B2 
                           => n148, ZN => n317);
   U235 : AOI22_X1 port map( A1 => A_neg(10), A2 => n152, B1 => A_signal(10), 
                           B2 => n143, ZN => n190);
   U236 : AOI222_X1 port map( A1 => A_shifted(52), A2 => n181, B1 => 
                           zeroSignal(52), B2 => n171, C1 => A_neg_shifted(52),
                           C2 => n161, ZN => n281);
   U237 : AOI22_X1 port map( A1 => A_neg(51), A2 => n155, B1 => A_signal(51), 
                           B2 => n146, ZN => n280);
   U238 : AOI222_X1 port map( A1 => A_shifted(49), A2 => n180, B1 => 
                           zeroSignal(49), B2 => n171, C1 => A_neg_shifted(49),
                           C2 => n161, ZN => n273);
   U239 : AOI22_X1 port map( A1 => A_neg(48), A2 => n155, B1 => A_signal(48), 
                           B2 => n146, ZN => n272);
   U240 : AOI22_X1 port map( A1 => A_neg(35), A2 => n154, B1 => A_signal(35), 
                           B2 => n145, ZN => n244);
   U241 : AOI222_X1 port map( A1 => A_shifted(46), A2 => n180, B1 => 
                           zeroSignal(46), B2 => n171, C1 => A_neg_shifted(46),
                           C2 => n161, ZN => n267);
   U242 : AOI22_X1 port map( A1 => A_neg(45), A2 => n155, B1 => A_signal(45), 
                           B2 => n146, ZN => n266);
   U243 : AOI22_X1 port map( A1 => A_neg(24), A2 => n153, B1 => A_signal(24), 
                           B2 => n144, ZN => n220);

end SYN_BEHAVIORAL_2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity MUX51_MuxNbit64_12 is

   port( zeroSignal, A_signal, A_neg, A_shifted, A_neg_shifted : in 
         std_logic_vector (63 downto 0);  Sel : in std_logic_vector (2 downto 
         0);  Y : out std_logic_vector (63 downto 0));

end MUX51_MuxNbit64_12;

architecture SYN_BEHAVIORAL_2 of MUX51_MuxNbit64_12 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, 
      n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, 
      n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, 
      n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, 
      n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, 
      n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, 
      n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, 
      n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, 
      n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, 
      n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, 
      n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, 
      n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, 
      n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, 
      n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, 
      n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319 : 
      std_logic;

begin
   
   U1 : BUF_X1 port map( A => n141, Z => n167);
   U2 : BUF_X1 port map( A => n185, Z => n183);
   U3 : BUF_X1 port map( A => n142, Z => n158);
   U4 : BUF_X1 port map( A => n151, Z => n149);
   U5 : BUF_X1 port map( A => n142, Z => n159);
   U6 : BUF_X1 port map( A => n141, Z => n166);
   U7 : BUF_X1 port map( A => n185, Z => n184);
   U8 : BUF_X1 port map( A => n151, Z => n150);
   U9 : BUF_X1 port map( A => n176, Z => n175);
   U10 : BUF_X1 port map( A => n176, Z => n174);
   U11 : AND3_X1 port map( A1 => n318, A2 => n319, A3 => Sel(2), ZN => n141);
   U12 : NOR3_X1 port map( A1 => Sel(0), A2 => Sel(2), A3 => n319, ZN => n142);
   U13 : BUF_X1 port map( A => n183, Z => n182);
   U14 : BUF_X1 port map( A => n158, Z => n157);
   U15 : BUF_X1 port map( A => n149, Z => n148);
   U16 : BUF_X1 port map( A => n159, Z => n152);
   U17 : BUF_X1 port map( A => n167, Z => n160);
   U18 : BUF_X1 port map( A => n184, Z => n177);
   U19 : BUF_X1 port map( A => n150, Z => n143);
   U20 : BUF_X1 port map( A => n166, Z => n165);
   U21 : BUF_X1 port map( A => n166, Z => n164);
   U22 : BUF_X1 port map( A => n159, Z => n153);
   U23 : BUF_X1 port map( A => n184, Z => n178);
   U24 : BUF_X1 port map( A => n150, Z => n144);
   U25 : BUF_X1 port map( A => n166, Z => n163);
   U26 : BUF_X1 port map( A => n184, Z => n179);
   U27 : BUF_X1 port map( A => n159, Z => n154);
   U28 : BUF_X1 port map( A => n150, Z => n145);
   U29 : BUF_X1 port map( A => n167, Z => n162);
   U30 : BUF_X1 port map( A => n183, Z => n180);
   U31 : BUF_X1 port map( A => n158, Z => n155);
   U32 : BUF_X1 port map( A => n149, Z => n146);
   U33 : BUF_X1 port map( A => n167, Z => n161);
   U34 : BUF_X1 port map( A => n183, Z => n181);
   U35 : BUF_X1 port map( A => n158, Z => n156);
   U36 : BUF_X1 port map( A => n149, Z => n147);
   U37 : BUF_X1 port map( A => n175, Z => n169);
   U38 : BUF_X1 port map( A => n175, Z => n170);
   U39 : BUF_X1 port map( A => n174, Z => n171);
   U40 : BUF_X1 port map( A => n174, Z => n172);
   U41 : BUF_X1 port map( A => n175, Z => n168);
   U42 : BUF_X1 port map( A => n174, Z => n173);
   U43 : BUF_X1 port map( A => n315, Z => n185);
   U44 : NOR3_X1 port map( A1 => n318, A2 => Sel(2), A3 => n319, ZN => n315);
   U45 : INV_X1 port map( A => Sel(1), ZN => n319);
   U46 : BUF_X1 port map( A => n313, Z => n151);
   U47 : NOR3_X1 port map( A1 => Sel(1), A2 => Sel(2), A3 => n318, ZN => n313);
   U48 : INV_X1 port map( A => Sel(0), ZN => n318);
   U49 : BUF_X1 port map( A => n314, Z => n176);
   U50 : NOR2_X1 port map( A1 => n165, A2 => n186, ZN => n314);
   U51 : AOI21_X1 port map( B1 => n318, B2 => n319, A => Sel(2), ZN => n186);
   U52 : NAND2_X1 port map( A1 => n317, A2 => n316, ZN => Y(9));
   U53 : AOI22_X1 port map( A1 => A_neg(9), A2 => n157, B1 => A_signal(9), B2 
                           => n148, ZN => n317);
   U54 : NAND2_X1 port map( A1 => n312, A2 => n311, ZN => Y(8));
   U55 : AOI222_X1 port map( A1 => A_shifted(8), A2 => n182, B1 => 
                           zeroSignal(8), B2 => n173, C1 => A_neg_shifted(8), 
                           C2 => n160, ZN => n311);
   U56 : NAND2_X1 port map( A1 => n190, A2 => n189, ZN => Y(10));
   U57 : AOI222_X1 port map( A1 => A_shifted(10), A2 => n177, B1 => 
                           zeroSignal(10), B2 => n168, C1 => A_neg_shifted(10),
                           C2 => n165, ZN => n189);
   U58 : AOI22_X1 port map( A1 => A_neg(10), A2 => n152, B1 => A_signal(10), B2
                           => n143, ZN => n190);
   U59 : AOI222_X1 port map( A1 => A_shifted(11), A2 => n177, B1 => 
                           zeroSignal(11), B2 => n168, C1 => A_neg_shifted(11),
                           C2 => n165, ZN => n191);
   U60 : AOI22_X1 port map( A1 => A_neg(12), A2 => n152, B1 => A_signal(12), B2
                           => n143, ZN => n194);
   U61 : AOI222_X1 port map( A1 => A_shifted(13), A2 => n177, B1 => 
                           zeroSignal(13), B2 => n168, C1 => A_neg_shifted(13),
                           C2 => n164, ZN => n195);
   U62 : NAND2_X1 port map( A1 => n218, A2 => n217, ZN => Y(23));
   U63 : AOI222_X1 port map( A1 => A_shifted(23), A2 => n178, B1 => 
                           zeroSignal(23), B2 => n169, C1 => A_neg_shifted(23),
                           C2 => n164, ZN => n217);
   U64 : AOI22_X1 port map( A1 => A_neg(23), A2 => n153, B1 => A_signal(23), B2
                           => n144, ZN => n218);
   U65 : NAND2_X1 port map( A1 => n214, A2 => n213, ZN => Y(21));
   U66 : AOI222_X1 port map( A1 => A_shifted(21), A2 => n178, B1 => 
                           zeroSignal(21), B2 => n169, C1 => A_neg_shifted(21),
                           C2 => n164, ZN => n213);
   U67 : AOI22_X1 port map( A1 => A_neg(21), A2 => n153, B1 => A_signal(21), B2
                           => n144, ZN => n214);
   U68 : NAND2_X1 port map( A1 => n216, A2 => n215, ZN => Y(22));
   U69 : AOI222_X1 port map( A1 => A_shifted(22), A2 => n178, B1 => 
                           zeroSignal(22), B2 => n169, C1 => A_neg_shifted(22),
                           C2 => n164, ZN => n215);
   U70 : AOI22_X1 port map( A1 => A_neg(22), A2 => n153, B1 => A_signal(22), B2
                           => n144, ZN => n216);
   U71 : NAND2_X1 port map( A1 => n222, A2 => n221, ZN => Y(25));
   U72 : AOI222_X1 port map( A1 => A_shifted(25), A2 => n178, B1 => 
                           zeroSignal(25), B2 => n169, C1 => A_neg_shifted(25),
                           C2 => n163, ZN => n221);
   U73 : AOI22_X1 port map( A1 => A_neg(25), A2 => n153, B1 => A_signal(25), B2
                           => n144, ZN => n222);
   U74 : NAND2_X1 port map( A1 => n220, A2 => n219, ZN => Y(24));
   U75 : AOI222_X1 port map( A1 => A_shifted(24), A2 => n178, B1 => 
                           zeroSignal(24), B2 => n169, C1 => A_neg_shifted(24),
                           C2 => n163, ZN => n219);
   U76 : AOI22_X1 port map( A1 => A_neg(24), A2 => n153, B1 => A_signal(24), B2
                           => n144, ZN => n220);
   U77 : NAND2_X1 port map( A1 => n226, A2 => n225, ZN => Y(27));
   U78 : AOI222_X1 port map( A1 => A_shifted(27), A2 => n178, B1 => 
                           zeroSignal(27), B2 => n169, C1 => A_neg_shifted(27),
                           C2 => n163, ZN => n225);
   U79 : AOI22_X1 port map( A1 => A_neg(27), A2 => n153, B1 => A_signal(27), B2
                           => n144, ZN => n226);
   U80 : NAND2_X1 port map( A1 => n230, A2 => n229, ZN => Y(29));
   U81 : AOI222_X1 port map( A1 => A_shifted(29), A2 => n178, B1 => 
                           zeroSignal(29), B2 => n169, C1 => A_neg_shifted(29),
                           C2 => n163, ZN => n229);
   U82 : AOI22_X1 port map( A1 => A_neg(29), A2 => n153, B1 => A_signal(29), B2
                           => n144, ZN => n230);
   U83 : NAND2_X1 port map( A1 => n228, A2 => n227, ZN => Y(28));
   U84 : AOI222_X1 port map( A1 => A_shifted(28), A2 => n178, B1 => 
                           zeroSignal(28), B2 => n169, C1 => A_neg_shifted(28),
                           C2 => n163, ZN => n227);
   U85 : AOI22_X1 port map( A1 => A_neg(28), A2 => n153, B1 => A_signal(28), B2
                           => n144, ZN => n228);
   U86 : NAND2_X1 port map( A1 => n234, A2 => n233, ZN => Y(30));
   U87 : AOI222_X1 port map( A1 => A_shifted(30), A2 => n179, B1 => 
                           zeroSignal(30), B2 => n169, C1 => A_neg_shifted(30),
                           C2 => n163, ZN => n233);
   U88 : AOI22_X1 port map( A1 => A_neg(30), A2 => n153, B1 => A_signal(30), B2
                           => n144, ZN => n234);
   U89 : NAND2_X1 port map( A1 => n236, A2 => n235, ZN => Y(31));
   U90 : AOI222_X1 port map( A1 => A_shifted(31), A2 => n179, B1 => 
                           zeroSignal(31), B2 => n170, C1 => A_neg_shifted(31),
                           C2 => n163, ZN => n235);
   U91 : AOI22_X1 port map( A1 => A_neg(31), A2 => n154, B1 => A_signal(31), B2
                           => n145, ZN => n236);
   U92 : NAND2_X1 port map( A1 => n238, A2 => n237, ZN => Y(32));
   U93 : AOI222_X1 port map( A1 => A_shifted(32), A2 => n179, B1 => 
                           zeroSignal(32), B2 => n170, C1 => A_neg_shifted(32),
                           C2 => n163, ZN => n237);
   U94 : AOI22_X1 port map( A1 => A_neg(32), A2 => n154, B1 => A_signal(32), B2
                           => n145, ZN => n238);
   U95 : NAND2_X1 port map( A1 => n242, A2 => n241, ZN => Y(34));
   U96 : AOI222_X1 port map( A1 => A_shifted(34), A2 => n179, B1 => 
                           zeroSignal(34), B2 => n170, C1 => A_neg_shifted(34),
                           C2 => n163, ZN => n241);
   U97 : AOI22_X1 port map( A1 => A_neg(34), A2 => n154, B1 => A_signal(34), B2
                           => n145, ZN => n242);
   U98 : NAND2_X1 port map( A1 => n240, A2 => n239, ZN => Y(33));
   U99 : AOI222_X1 port map( A1 => A_shifted(33), A2 => n179, B1 => 
                           zeroSignal(33), B2 => n170, C1 => A_neg_shifted(33),
                           C2 => n163, ZN => n239);
   U100 : AOI22_X1 port map( A1 => A_neg(33), A2 => n154, B1 => A_signal(33), 
                           B2 => n145, ZN => n240);
   U101 : NAND2_X1 port map( A1 => n244, A2 => n243, ZN => Y(35));
   U102 : AOI222_X1 port map( A1 => A_shifted(35), A2 => n179, B1 => 
                           zeroSignal(35), B2 => n170, C1 => A_neg_shifted(35),
                           C2 => n162, ZN => n243);
   U103 : AOI22_X1 port map( A1 => A_neg(35), A2 => n154, B1 => A_signal(35), 
                           B2 => n145, ZN => n244);
   U104 : NAND2_X1 port map( A1 => n246, A2 => n245, ZN => Y(36));
   U105 : AOI222_X1 port map( A1 => A_shifted(36), A2 => n179, B1 => 
                           zeroSignal(36), B2 => n170, C1 => A_neg_shifted(36),
                           C2 => n162, ZN => n245);
   U106 : AOI22_X1 port map( A1 => A_neg(36), A2 => n154, B1 => A_signal(36), 
                           B2 => n145, ZN => n246);
   U107 : AOI22_X1 port map( A1 => A_neg(15), A2 => n152, B1 => A_signal(15), 
                           B2 => n143, ZN => n200);
   U108 : NAND2_X1 port map( A1 => n250, A2 => n249, ZN => Y(38));
   U109 : AOI222_X1 port map( A1 => A_shifted(38), A2 => n179, B1 => 
                           zeroSignal(38), B2 => n170, C1 => A_neg_shifted(38),
                           C2 => n162, ZN => n249);
   U110 : AOI22_X1 port map( A1 => A_neg(38), A2 => n154, B1 => A_signal(38), 
                           B2 => n145, ZN => n250);
   U111 : NAND2_X1 port map( A1 => n224, A2 => n223, ZN => Y(26));
   U112 : AOI22_X1 port map( A1 => A_neg(26), A2 => n153, B1 => A_signal(26), 
                           B2 => n144, ZN => n224);
   U113 : AOI222_X1 port map( A1 => A_shifted(26), A2 => n178, B1 => 
                           zeroSignal(26), B2 => n169, C1 => A_neg_shifted(26),
                           C2 => n163, ZN => n223);
   U114 : NAND2_X1 port map( A1 => n252, A2 => n251, ZN => Y(39));
   U115 : AOI222_X1 port map( A1 => A_shifted(39), A2 => n179, B1 => 
                           zeroSignal(39), B2 => n170, C1 => A_neg_shifted(39),
                           C2 => n162, ZN => n251);
   U116 : AOI22_X1 port map( A1 => A_neg(39), A2 => n154, B1 => A_signal(39), 
                           B2 => n145, ZN => n252);
   U117 : NAND2_X1 port map( A1 => n256, A2 => n255, ZN => Y(40));
   U118 : AOI222_X1 port map( A1 => A_shifted(40), A2 => n180, B1 => 
                           zeroSignal(40), B2 => n170, C1 => A_neg_shifted(40),
                           C2 => n162, ZN => n255);
   U119 : AOI22_X1 port map( A1 => A_neg(40), A2 => n154, B1 => A_signal(40), 
                           B2 => n145, ZN => n256);
   U120 : NAND2_X1 port map( A1 => n206, A2 => n205, ZN => Y(18));
   U121 : AOI222_X1 port map( A1 => A_shifted(18), A2 => n177, B1 => 
                           zeroSignal(18), B2 => n168, C1 => A_neg_shifted(18),
                           C2 => n164, ZN => n205);
   U122 : AOI22_X1 port map( A1 => A_neg(18), A2 => n152, B1 => A_signal(18), 
                           B2 => n143, ZN => n206);
   U123 : NAND2_X1 port map( A1 => n272, A2 => n271, ZN => Y(48));
   U124 : AOI222_X1 port map( A1 => A_shifted(48), A2 => n180, B1 => 
                           zeroSignal(48), B2 => n171, C1 => A_neg_shifted(48),
                           C2 => n161, ZN => n271);
   U125 : AOI22_X1 port map( A1 => A_neg(48), A2 => n155, B1 => A_signal(48), 
                           B2 => n146, ZN => n272);
   U126 : NAND2_X1 port map( A1 => n258, A2 => n257, ZN => Y(41));
   U127 : AOI222_X1 port map( A1 => A_shifted(41), A2 => n180, B1 => 
                           zeroSignal(41), B2 => n170, C1 => A_neg_shifted(41),
                           C2 => n162, ZN => n257);
   U128 : AOI22_X1 port map( A1 => A_neg(41), A2 => n154, B1 => A_signal(41), 
                           B2 => n145, ZN => n258);
   U129 : NAND2_X1 port map( A1 => n212, A2 => n211, ZN => Y(20));
   U130 : AOI222_X1 port map( A1 => A_shifted(20), A2 => n178, B1 => 
                           zeroSignal(20), B2 => n169, C1 => A_neg_shifted(20),
                           C2 => n164, ZN => n211);
   U131 : AOI22_X1 port map( A1 => A_neg(20), A2 => n153, B1 => A_signal(20), 
                           B2 => n144, ZN => n212);
   U132 : NAND2_X1 port map( A1 => n248, A2 => n247, ZN => Y(37));
   U133 : AOI22_X1 port map( A1 => A_neg(37), A2 => n154, B1 => A_signal(37), 
                           B2 => n145, ZN => n248);
   U134 : AOI222_X1 port map( A1 => A_shifted(37), A2 => n179, B1 => 
                           zeroSignal(37), B2 => n170, C1 => A_neg_shifted(37),
                           C2 => n162, ZN => n247);
   U135 : NAND2_X1 port map( A1 => n202, A2 => n201, ZN => Y(16));
   U136 : AOI22_X1 port map( A1 => A_neg(16), A2 => n152, B1 => A_signal(16), 
                           B2 => n143, ZN => n202);
   U137 : AOI222_X1 port map( A1 => A_shifted(16), A2 => n177, B1 => 
                           zeroSignal(16), B2 => n168, C1 => A_neg_shifted(16),
                           C2 => n164, ZN => n201);
   U138 : NAND2_X1 port map( A1 => n208, A2 => n207, ZN => Y(19));
   U139 : AOI22_X1 port map( A1 => A_neg(19), A2 => n152, B1 => A_signal(19), 
                           B2 => n143, ZN => n208);
   U140 : AOI222_X1 port map( A1 => A_shifted(19), A2 => n177, B1 => 
                           zeroSignal(19), B2 => n168, C1 => A_neg_shifted(19),
                           C2 => n164, ZN => n207);
   U141 : NAND2_X1 port map( A1 => n274, A2 => n273, ZN => Y(49));
   U142 : AOI22_X1 port map( A1 => A_neg(49), A2 => n155, B1 => A_signal(49), 
                           B2 => n146, ZN => n274);
   U143 : AOI222_X1 port map( A1 => A_shifted(49), A2 => n180, B1 => 
                           zeroSignal(49), B2 => n171, C1 => A_neg_shifted(49),
                           C2 => n161, ZN => n273);
   U144 : NAND2_X1 port map( A1 => n260, A2 => n259, ZN => Y(42));
   U145 : AOI222_X1 port map( A1 => A_shifted(42), A2 => n180, B1 => 
                           zeroSignal(42), B2 => n171, C1 => A_neg_shifted(42),
                           C2 => n162, ZN => n259);
   U146 : AOI22_X1 port map( A1 => A_neg(42), A2 => n155, B1 => A_signal(42), 
                           B2 => n146, ZN => n260);
   U147 : NAND2_X1 port map( A1 => n262, A2 => n261, ZN => Y(43));
   U148 : AOI222_X1 port map( A1 => A_shifted(43), A2 => n180, B1 => 
                           zeroSignal(43), B2 => n171, C1 => A_neg_shifted(43),
                           C2 => n162, ZN => n261);
   U149 : AOI22_X1 port map( A1 => A_neg(43), A2 => n155, B1 => A_signal(43), 
                           B2 => n146, ZN => n262);
   U150 : NAND2_X1 port map( A1 => n264, A2 => n263, ZN => Y(44));
   U151 : AOI222_X1 port map( A1 => A_shifted(44), A2 => n180, B1 => 
                           zeroSignal(44), B2 => n171, C1 => A_neg_shifted(44),
                           C2 => n162, ZN => n263);
   U152 : AOI22_X1 port map( A1 => A_neg(44), A2 => n155, B1 => A_signal(44), 
                           B2 => n146, ZN => n264);
   U153 : NAND2_X1 port map( A1 => n204, A2 => n203, ZN => Y(17));
   U154 : AOI22_X1 port map( A1 => A_neg(17), A2 => n152, B1 => A_signal(17), 
                           B2 => n143, ZN => n204);
   U155 : AOI222_X1 port map( A1 => A_shifted(17), A2 => n177, B1 => 
                           zeroSignal(17), B2 => n168, C1 => A_neg_shifted(17),
                           C2 => n164, ZN => n203);
   U156 : NAND2_X1 port map( A1 => n266, A2 => n265, ZN => Y(45));
   U157 : AOI222_X1 port map( A1 => A_shifted(45), A2 => n180, B1 => 
                           zeroSignal(45), B2 => n171, C1 => A_neg_shifted(45),
                           C2 => n162, ZN => n265);
   U158 : AOI22_X1 port map( A1 => A_neg(45), A2 => n155, B1 => A_signal(45), 
                           B2 => n146, ZN => n266);
   U159 : NAND2_X1 port map( A1 => n268, A2 => n267, ZN => Y(46));
   U160 : AOI22_X1 port map( A1 => A_neg(46), A2 => n155, B1 => A_signal(46), 
                           B2 => n146, ZN => n268);
   U161 : AOI222_X1 port map( A1 => A_shifted(46), A2 => n180, B1 => 
                           zeroSignal(46), B2 => n171, C1 => A_neg_shifted(46),
                           C2 => n161, ZN => n267);
   U162 : NAND2_X1 port map( A1 => n306, A2 => n305, ZN => Y(63));
   U163 : AOI222_X1 port map( A1 => A_shifted(63), A2 => n182, B1 => 
                           zeroSignal(63), B2 => n172, C1 => A_neg_shifted(63),
                           C2 => n160, ZN => n305);
   U164 : AOI22_X1 port map( A1 => A_neg(63), A2 => n156, B1 => A_signal(63), 
                           B2 => n147, ZN => n306);
   U165 : NAND2_X1 port map( A1 => n304, A2 => n303, ZN => Y(62));
   U166 : AOI222_X1 port map( A1 => A_shifted(62), A2 => n182, B1 => 
                           zeroSignal(62), B2 => n172, C1 => A_neg_shifted(62),
                           C2 => n160, ZN => n303);
   U167 : AOI22_X1 port map( A1 => A_neg(62), A2 => n156, B1 => A_signal(62), 
                           B2 => n147, ZN => n304);
   U168 : NAND2_X1 port map( A1 => n296, A2 => n295, ZN => Y(59));
   U169 : AOI222_X1 port map( A1 => A_shifted(59), A2 => n181, B1 => 
                           zeroSignal(59), B2 => n172, C1 => A_neg_shifted(59),
                           C2 => n160, ZN => n295);
   U170 : AOI22_X1 port map( A1 => A_neg(59), A2 => n156, B1 => A_signal(59), 
                           B2 => n147, ZN => n296);
   U171 : NAND2_X1 port map( A1 => n302, A2 => n301, ZN => Y(61));
   U172 : AOI222_X1 port map( A1 => A_shifted(61), A2 => n182, B1 => 
                           zeroSignal(61), B2 => n172, C1 => A_neg_shifted(61),
                           C2 => n160, ZN => n301);
   U173 : AOI22_X1 port map( A1 => A_neg(61), A2 => n156, B1 => A_signal(61), 
                           B2 => n147, ZN => n302);
   U174 : NAND2_X1 port map( A1 => n300, A2 => n299, ZN => Y(60));
   U175 : AOI222_X1 port map( A1 => A_shifted(60), A2 => n182, B1 => 
                           zeroSignal(60), B2 => n172, C1 => A_neg_shifted(60),
                           C2 => n160, ZN => n299);
   U176 : AOI22_X1 port map( A1 => A_neg(60), A2 => n156, B1 => A_signal(60), 
                           B2 => n147, ZN => n300);
   U177 : NAND2_X1 port map( A1 => n280, A2 => n279, ZN => Y(51));
   U178 : AOI22_X1 port map( A1 => A_neg(51), A2 => n155, B1 => A_signal(51), 
                           B2 => n146, ZN => n280);
   U179 : NAND2_X1 port map( A1 => n284, A2 => n283, ZN => Y(53));
   U180 : AOI222_X1 port map( A1 => A_shifted(53), A2 => n181, B1 => 
                           zeroSignal(53), B2 => n172, C1 => A_neg_shifted(53),
                           C2 => n161, ZN => n283);
   U181 : NAND2_X1 port map( A1 => n282, A2 => n281, ZN => Y(52));
   U182 : AOI222_X1 port map( A1 => A_shifted(52), A2 => n181, B1 => 
                           zeroSignal(52), B2 => n171, C1 => A_neg_shifted(52),
                           C2 => n161, ZN => n281);
   U183 : AOI22_X1 port map( A1 => A_neg(52), A2 => n155, B1 => A_signal(52), 
                           B2 => n146, ZN => n282);
   U184 : NAND2_X1 port map( A1 => n278, A2 => n277, ZN => Y(50));
   U185 : AOI222_X1 port map( A1 => A_shifted(50), A2 => n181, B1 => 
                           zeroSignal(50), B2 => n171, C1 => A_neg_shifted(50),
                           C2 => n161, ZN => n277);
   U186 : NAND2_X1 port map( A1 => n286, A2 => n285, ZN => Y(54));
   U187 : AOI22_X1 port map( A1 => A_neg(54), A2 => n156, B1 => A_signal(54), 
                           B2 => n147, ZN => n286);
   U188 : NAND2_X1 port map( A1 => n288, A2 => n287, ZN => Y(55));
   U189 : AOI222_X1 port map( A1 => A_shifted(55), A2 => n181, B1 => 
                           zeroSignal(55), B2 => n172, C1 => A_neg_shifted(55),
                           C2 => n161, ZN => n287);
   U190 : AOI22_X1 port map( A1 => A_neg(55), A2 => n156, B1 => A_signal(55), 
                           B2 => n147, ZN => n288);
   U191 : NAND2_X1 port map( A1 => n270, A2 => n269, ZN => Y(47));
   U192 : AOI222_X1 port map( A1 => A_shifted(47), A2 => n180, B1 => 
                           zeroSignal(47), B2 => n171, C1 => A_neg_shifted(47),
                           C2 => n161, ZN => n269);
   U193 : NAND2_X1 port map( A1 => n290, A2 => n289, ZN => Y(56));
   U194 : AOI222_X1 port map( A1 => A_shifted(56), A2 => n181, B1 => 
                           zeroSignal(56), B2 => n172, C1 => A_neg_shifted(56),
                           C2 => n161, ZN => n289);
   U195 : AOI22_X1 port map( A1 => A_neg(56), A2 => n156, B1 => A_signal(56), 
                           B2 => n147, ZN => n290);
   U196 : NAND2_X1 port map( A1 => n292, A2 => n291, ZN => Y(57));
   U197 : AOI222_X1 port map( A1 => A_shifted(57), A2 => n181, B1 => 
                           zeroSignal(57), B2 => n172, C1 => A_neg_shifted(57),
                           C2 => n160, ZN => n291);
   U198 : AOI22_X1 port map( A1 => A_neg(57), A2 => n156, B1 => A_signal(57), 
                           B2 => n147, ZN => n292);
   U199 : NAND2_X1 port map( A1 => n294, A2 => n293, ZN => Y(58));
   U200 : AOI222_X1 port map( A1 => A_shifted(58), A2 => n181, B1 => 
                           zeroSignal(58), B2 => n172, C1 => A_neg_shifted(58),
                           C2 => n160, ZN => n293);
   U201 : AOI22_X1 port map( A1 => A_neg(58), A2 => n156, B1 => A_signal(58), 
                           B2 => n147, ZN => n294);
   U202 : NAND2_X1 port map( A1 => n188, A2 => n187, ZN => Y(0));
   U203 : AOI22_X1 port map( A1 => A_neg(0), A2 => n152, B1 => A_signal(0), B2 
                           => n143, ZN => n188);
   U204 : AOI222_X1 port map( A1 => A_shifted(0), A2 => n177, B1 => 
                           zeroSignal(0), B2 => n168, C1 => A_neg_shifted(0), 
                           C2 => n165, ZN => n187);
   U205 : NAND2_X1 port map( A1 => n210, A2 => n209, ZN => Y(1));
   U206 : AOI22_X1 port map( A1 => A_neg(1), A2 => n152, B1 => A_signal(1), B2 
                           => n143, ZN => n210);
   U207 : AOI222_X1 port map( A1 => A_shifted(1), A2 => n178, B1 => 
                           zeroSignal(1), B2 => n168, C1 => A_neg_shifted(1), 
                           C2 => n164, ZN => n209);
   U208 : NAND2_X1 port map( A1 => n232, A2 => n231, ZN => Y(2));
   U209 : AOI22_X1 port map( A1 => A_neg(2), A2 => n153, B1 => A_signal(2), B2 
                           => n144, ZN => n232);
   U210 : AOI222_X1 port map( A1 => A_shifted(2), A2 => n179, B1 => 
                           zeroSignal(2), B2 => n169, C1 => A_neg_shifted(2), 
                           C2 => n163, ZN => n231);
   U211 : NAND2_X1 port map( A1 => n254, A2 => n253, ZN => Y(3));
   U212 : AOI22_X1 port map( A1 => A_neg(3), A2 => n154, B1 => A_signal(3), B2 
                           => n145, ZN => n254);
   U213 : AOI222_X1 port map( A1 => A_shifted(3), A2 => n180, B1 => 
                           zeroSignal(3), B2 => n170, C1 => A_neg_shifted(3), 
                           C2 => n162, ZN => n253);
   U214 : NAND2_X1 port map( A1 => n276, A2 => n275, ZN => Y(4));
   U215 : AOI22_X1 port map( A1 => A_neg(4), A2 => n155, B1 => A_signal(4), B2 
                           => n146, ZN => n276);
   U216 : AOI222_X1 port map( A1 => A_shifted(4), A2 => n181, B1 => 
                           zeroSignal(4), B2 => n171, C1 => A_neg_shifted(4), 
                           C2 => n161, ZN => n275);
   U217 : NAND2_X1 port map( A1 => n298, A2 => n297, ZN => Y(5));
   U218 : AOI22_X1 port map( A1 => A_neg(5), A2 => n156, B1 => A_signal(5), B2 
                           => n147, ZN => n298);
   U219 : AOI222_X1 port map( A1 => A_shifted(5), A2 => n182, B1 => 
                           zeroSignal(5), B2 => n172, C1 => A_neg_shifted(5), 
                           C2 => n160, ZN => n297);
   U220 : NAND2_X1 port map( A1 => n308, A2 => n307, ZN => Y(6));
   U221 : AOI22_X1 port map( A1 => A_neg(6), A2 => n157, B1 => A_signal(6), B2 
                           => n148, ZN => n308);
   U222 : AOI222_X1 port map( A1 => A_shifted(6), A2 => n182, B1 => 
                           zeroSignal(6), B2 => n173, C1 => A_neg_shifted(6), 
                           C2 => n160, ZN => n307);
   U223 : NAND2_X1 port map( A1 => n310, A2 => n309, ZN => Y(7));
   U224 : AOI22_X1 port map( A1 => A_neg(7), A2 => n157, B1 => A_signal(7), B2 
                           => n148, ZN => n310);
   U225 : AOI222_X1 port map( A1 => A_shifted(7), A2 => n182, B1 => 
                           zeroSignal(7), B2 => n173, C1 => A_neg_shifted(7), 
                           C2 => n160, ZN => n309);
   U226 : AOI222_X1 port map( A1 => A_shifted(9), A2 => n182, B1 => 
                           zeroSignal(9), B2 => n173, C1 => A_neg_shifted(9), 
                           C2 => n160, ZN => n316);
   U227 : AOI22_X1 port map( A1 => A_neg(8), A2 => n157, B1 => A_signal(8), B2 
                           => n148, ZN => n312);
   U228 : AOI222_X1 port map( A1 => A_shifted(15), A2 => n177, B1 => 
                           zeroSignal(15), B2 => n168, C1 => A_neg_shifted(15),
                           C2 => n164, ZN => n199);
   U229 : AOI22_X1 port map( A1 => A_neg(14), A2 => n152, B1 => A_signal(14), 
                           B2 => n143, ZN => n198);
   U230 : NAND2_X1 port map( A1 => n200, A2 => n199, ZN => Y(15));
   U231 : AOI222_X1 port map( A1 => A_shifted(14), A2 => n177, B1 => 
                           zeroSignal(14), B2 => n168, C1 => A_neg_shifted(14),
                           C2 => n164, ZN => n197);
   U232 : AOI22_X1 port map( A1 => A_neg(13), A2 => n152, B1 => A_signal(13), 
                           B2 => n143, ZN => n196);
   U233 : NAND2_X1 port map( A1 => n198, A2 => n197, ZN => Y(14));
   U234 : NAND2_X1 port map( A1 => n196, A2 => n195, ZN => Y(13));
   U235 : AOI222_X1 port map( A1 => A_shifted(12), A2 => n177, B1 => 
                           zeroSignal(12), B2 => n168, C1 => A_neg_shifted(12),
                           C2 => n165, ZN => n193);
   U236 : AOI22_X1 port map( A1 => A_neg(11), A2 => n152, B1 => A_signal(11), 
                           B2 => n143, ZN => n192);
   U237 : NAND2_X1 port map( A1 => n194, A2 => n193, ZN => Y(12));
   U238 : NAND2_X1 port map( A1 => n192, A2 => n191, ZN => Y(11));
   U239 : AOI222_X1 port map( A1 => A_shifted(54), A2 => n181, B1 => 
                           zeroSignal(54), B2 => n172, C1 => A_neg_shifted(54),
                           C2 => n161, ZN => n285);
   U240 : AOI22_X1 port map( A1 => A_neg(53), A2 => n156, B1 => A_signal(53), 
                           B2 => n147, ZN => n284);
   U241 : AOI222_X1 port map( A1 => A_shifted(51), A2 => n181, B1 => 
                           zeroSignal(51), B2 => n171, C1 => A_neg_shifted(51),
                           C2 => n161, ZN => n279);
   U242 : AOI22_X1 port map( A1 => A_neg(50), A2 => n155, B1 => A_signal(50), 
                           B2 => n146, ZN => n278);
   U243 : AOI22_X1 port map( A1 => A_neg(47), A2 => n155, B1 => A_signal(47), 
                           B2 => n146, ZN => n270);

end SYN_BEHAVIORAL_2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity MUX51_MuxNbit64_11 is

   port( zeroSignal, A_signal, A_neg, A_shifted, A_neg_shifted : in 
         std_logic_vector (63 downto 0);  Sel : in std_logic_vector (2 downto 
         0);  Y : out std_logic_vector (63 downto 0));

end MUX51_MuxNbit64_11;

architecture SYN_BEHAVIORAL_2 of MUX51_MuxNbit64_11 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, 
      n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, 
      n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, 
      n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, 
      n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, 
      n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, 
      n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, 
      n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, 
      n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, 
      n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, 
      n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, 
      n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, 
      n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, 
      n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, 
      n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319 : 
      std_logic;

begin
   
   U1 : BUF_X1 port map( A => n141, Z => n185);
   U2 : BUF_X1 port map( A => n151, Z => n150);
   U3 : BUF_X1 port map( A => n160, Z => n159);
   U4 : BUF_X1 port map( A => n142, Z => n167);
   U5 : BUF_X1 port map( A => n142, Z => n168);
   U6 : BUF_X1 port map( A => n141, Z => n184);
   U7 : BUF_X1 port map( A => n151, Z => n149);
   U8 : BUF_X1 port map( A => n160, Z => n158);
   U9 : BUF_X1 port map( A => n177, Z => n176);
   U10 : BUF_X1 port map( A => n177, Z => n175);
   U11 : NOR3_X1 port map( A1 => n318, A2 => Sel(2), A3 => n319, ZN => n141);
   U12 : BUF_X1 port map( A => n313, Z => n151);
   U13 : AND3_X1 port map( A1 => n318, A2 => n319, A3 => Sel(2), ZN => n142);
   U14 : BUF_X1 port map( A => n159, Z => n152);
   U15 : BUF_X1 port map( A => n150, Z => n143);
   U16 : BUF_X1 port map( A => n185, Z => n178);
   U17 : BUF_X1 port map( A => n167, Z => n166);
   U18 : BUF_X1 port map( A => n167, Z => n165);
   U19 : BUF_X1 port map( A => n159, Z => n153);
   U20 : BUF_X1 port map( A => n185, Z => n179);
   U21 : BUF_X1 port map( A => n150, Z => n144);
   U22 : BUF_X1 port map( A => n167, Z => n164);
   U23 : BUF_X1 port map( A => n185, Z => n180);
   U24 : BUF_X1 port map( A => n159, Z => n154);
   U25 : BUF_X1 port map( A => n150, Z => n145);
   U26 : BUF_X1 port map( A => n168, Z => n163);
   U27 : BUF_X1 port map( A => n184, Z => n181);
   U28 : BUF_X1 port map( A => n158, Z => n155);
   U29 : BUF_X1 port map( A => n149, Z => n146);
   U30 : BUF_X1 port map( A => n168, Z => n162);
   U31 : BUF_X1 port map( A => n184, Z => n182);
   U32 : BUF_X1 port map( A => n158, Z => n156);
   U33 : BUF_X1 port map( A => n149, Z => n147);
   U34 : BUF_X1 port map( A => n168, Z => n161);
   U35 : BUF_X1 port map( A => n184, Z => n183);
   U36 : BUF_X1 port map( A => n176, Z => n170);
   U37 : BUF_X1 port map( A => n176, Z => n171);
   U38 : BUF_X1 port map( A => n175, Z => n172);
   U39 : BUF_X1 port map( A => n175, Z => n173);
   U40 : BUF_X1 port map( A => n176, Z => n169);
   U41 : BUF_X1 port map( A => n158, Z => n157);
   U42 : BUF_X1 port map( A => n149, Z => n148);
   U43 : BUF_X1 port map( A => n175, Z => n174);
   U44 : BUF_X1 port map( A => n314, Z => n160);
   U45 : NOR3_X1 port map( A1 => Sel(0), A2 => Sel(2), A3 => n319, ZN => n314);
   U46 : INV_X1 port map( A => Sel(1), ZN => n319);
   U47 : INV_X1 port map( A => Sel(0), ZN => n318);
   U48 : NOR3_X1 port map( A1 => Sel(1), A2 => Sel(2), A3 => n318, ZN => n313);
   U49 : BUF_X1 port map( A => n315, Z => n177);
   U50 : NOR2_X1 port map( A1 => n166, A2 => n186, ZN => n315);
   U51 : AOI21_X1 port map( B1 => n318, B2 => n319, A => Sel(2), ZN => n186);
   U52 : NAND2_X1 port map( A1 => n192, A2 => n191, ZN => Y(11));
   U53 : AOI22_X1 port map( A1 => A_neg(11), A2 => n152, B1 => A_signal(11), B2
                           => n143, ZN => n192);
   U54 : NAND2_X1 port map( A1 => n190, A2 => n189, ZN => Y(10));
   U55 : AOI222_X1 port map( A1 => A_shifted(10), A2 => n178, B1 => 
                           zeroSignal(10), B2 => n169, C1 => A_neg_shifted(10),
                           C2 => n166, ZN => n189);
   U56 : NAND2_X1 port map( A1 => n194, A2 => n193, ZN => Y(12));
   U57 : AOI222_X1 port map( A1 => A_shifted(12), A2 => n178, B1 => 
                           zeroSignal(12), B2 => n169, C1 => A_neg_shifted(12),
                           C2 => n166, ZN => n193);
   U58 : AOI22_X1 port map( A1 => A_neg(12), A2 => n152, B1 => A_signal(12), B2
                           => n143, ZN => n194);
   U59 : AOI222_X1 port map( A1 => A_shifted(13), A2 => n178, B1 => 
                           zeroSignal(13), B2 => n169, C1 => A_neg_shifted(13),
                           C2 => n165, ZN => n195);
   U60 : AOI22_X1 port map( A1 => A_neg(14), A2 => n152, B1 => A_signal(14), B2
                           => n143, ZN => n198);
   U61 : AOI222_X1 port map( A1 => A_shifted(15), A2 => n178, B1 => 
                           zeroSignal(15), B2 => n169, C1 => A_neg_shifted(15),
                           C2 => n165, ZN => n199);
   U62 : NAND2_X1 port map( A1 => n272, A2 => n271, ZN => Y(48));
   U63 : AOI22_X1 port map( A1 => A_neg(48), A2 => n155, B1 => A_signal(48), B2
                           => n146, ZN => n272);
   U64 : AOI222_X1 port map( A1 => A_shifted(48), A2 => n181, B1 => 
                           zeroSignal(48), B2 => n172, C1 => A_neg_shifted(48),
                           C2 => n162, ZN => n271);
   U65 : NAND2_X1 port map( A1 => n222, A2 => n221, ZN => Y(25));
   U66 : AOI222_X1 port map( A1 => A_shifted(25), A2 => n179, B1 => 
                           zeroSignal(25), B2 => n170, C1 => A_neg_shifted(25),
                           C2 => n164, ZN => n221);
   U67 : AOI22_X1 port map( A1 => A_neg(25), A2 => n153, B1 => A_signal(25), B2
                           => n144, ZN => n222);
   U68 : NAND2_X1 port map( A1 => n218, A2 => n217, ZN => Y(23));
   U69 : AOI222_X1 port map( A1 => A_shifted(23), A2 => n179, B1 => 
                           zeroSignal(23), B2 => n170, C1 => A_neg_shifted(23),
                           C2 => n165, ZN => n217);
   U70 : AOI22_X1 port map( A1 => A_neg(23), A2 => n153, B1 => A_signal(23), B2
                           => n144, ZN => n218);
   U71 : NAND2_X1 port map( A1 => n220, A2 => n219, ZN => Y(24));
   U72 : AOI222_X1 port map( A1 => A_shifted(24), A2 => n179, B1 => 
                           zeroSignal(24), B2 => n170, C1 => A_neg_shifted(24),
                           C2 => n164, ZN => n219);
   U73 : AOI22_X1 port map( A1 => A_neg(24), A2 => n153, B1 => A_signal(24), B2
                           => n144, ZN => n220);
   U74 : NAND2_X1 port map( A1 => n226, A2 => n225, ZN => Y(27));
   U75 : AOI222_X1 port map( A1 => A_shifted(27), A2 => n179, B1 => 
                           zeroSignal(27), B2 => n170, C1 => A_neg_shifted(27),
                           C2 => n164, ZN => n225);
   U76 : AOI22_X1 port map( A1 => A_neg(27), A2 => n153, B1 => A_signal(27), B2
                           => n144, ZN => n226);
   U77 : NAND2_X1 port map( A1 => n224, A2 => n223, ZN => Y(26));
   U78 : AOI222_X1 port map( A1 => A_shifted(26), A2 => n179, B1 => 
                           zeroSignal(26), B2 => n170, C1 => A_neg_shifted(26),
                           C2 => n164, ZN => n223);
   U79 : AOI22_X1 port map( A1 => A_neg(26), A2 => n153, B1 => A_signal(26), B2
                           => n144, ZN => n224);
   U80 : NAND2_X1 port map( A1 => n230, A2 => n229, ZN => Y(29));
   U81 : AOI222_X1 port map( A1 => A_shifted(29), A2 => n179, B1 => 
                           zeroSignal(29), B2 => n170, C1 => A_neg_shifted(29),
                           C2 => n164, ZN => n229);
   U82 : AOI22_X1 port map( A1 => A_neg(29), A2 => n153, B1 => A_signal(29), B2
                           => n144, ZN => n230);
   U83 : NAND2_X1 port map( A1 => n234, A2 => n233, ZN => Y(30));
   U84 : AOI222_X1 port map( A1 => A_shifted(30), A2 => n180, B1 => 
                           zeroSignal(30), B2 => n170, C1 => A_neg_shifted(30),
                           C2 => n164, ZN => n233);
   U85 : AOI22_X1 port map( A1 => A_neg(30), A2 => n153, B1 => A_signal(30), B2
                           => n144, ZN => n234);
   U86 : NAND2_X1 port map( A1 => n236, A2 => n235, ZN => Y(31));
   U87 : AOI222_X1 port map( A1 => A_shifted(31), A2 => n180, B1 => 
                           zeroSignal(31), B2 => n171, C1 => A_neg_shifted(31),
                           C2 => n164, ZN => n235);
   U88 : AOI22_X1 port map( A1 => A_neg(31), A2 => n154, B1 => A_signal(31), B2
                           => n145, ZN => n236);
   U89 : NAND2_X1 port map( A1 => n238, A2 => n237, ZN => Y(32));
   U90 : AOI222_X1 port map( A1 => A_shifted(32), A2 => n180, B1 => 
                           zeroSignal(32), B2 => n171, C1 => A_neg_shifted(32),
                           C2 => n164, ZN => n237);
   U91 : AOI22_X1 port map( A1 => A_neg(32), A2 => n154, B1 => A_signal(32), B2
                           => n145, ZN => n238);
   U92 : NAND2_X1 port map( A1 => n242, A2 => n241, ZN => Y(34));
   U93 : AOI222_X1 port map( A1 => A_shifted(34), A2 => n180, B1 => 
                           zeroSignal(34), B2 => n171, C1 => A_neg_shifted(34),
                           C2 => n164, ZN => n241);
   U94 : AOI22_X1 port map( A1 => A_neg(34), A2 => n154, B1 => A_signal(34), B2
                           => n145, ZN => n242);
   U95 : NAND2_X1 port map( A1 => n240, A2 => n239, ZN => Y(33));
   U96 : AOI222_X1 port map( A1 => A_shifted(33), A2 => n180, B1 => 
                           zeroSignal(33), B2 => n171, C1 => A_neg_shifted(33),
                           C2 => n164, ZN => n239);
   U97 : AOI22_X1 port map( A1 => A_neg(33), A2 => n154, B1 => A_signal(33), B2
                           => n145, ZN => n240);
   U98 : NAND2_X1 port map( A1 => n244, A2 => n243, ZN => Y(35));
   U99 : AOI222_X1 port map( A1 => A_shifted(35), A2 => n180, B1 => 
                           zeroSignal(35), B2 => n171, C1 => A_neg_shifted(35),
                           C2 => n163, ZN => n243);
   U100 : AOI22_X1 port map( A1 => A_neg(35), A2 => n154, B1 => A_signal(35), 
                           B2 => n145, ZN => n244);
   U101 : NAND2_X1 port map( A1 => n246, A2 => n245, ZN => Y(36));
   U102 : AOI222_X1 port map( A1 => A_shifted(36), A2 => n180, B1 => 
                           zeroSignal(36), B2 => n171, C1 => A_neg_shifted(36),
                           C2 => n163, ZN => n245);
   U103 : AOI22_X1 port map( A1 => A_neg(36), A2 => n154, B1 => A_signal(36), 
                           B2 => n145, ZN => n246);
   U104 : NAND2_X1 port map( A1 => n248, A2 => n247, ZN => Y(37));
   U105 : AOI222_X1 port map( A1 => A_shifted(37), A2 => n180, B1 => 
                           zeroSignal(37), B2 => n171, C1 => A_neg_shifted(37),
                           C2 => n163, ZN => n247);
   U106 : AOI22_X1 port map( A1 => A_neg(37), A2 => n154, B1 => A_signal(37), 
                           B2 => n145, ZN => n248);
   U107 : NAND2_X1 port map( A1 => n250, A2 => n249, ZN => Y(38));
   U108 : AOI222_X1 port map( A1 => A_shifted(38), A2 => n180, B1 => 
                           zeroSignal(38), B2 => n171, C1 => A_neg_shifted(38),
                           C2 => n163, ZN => n249);
   U109 : AOI22_X1 port map( A1 => A_neg(38), A2 => n154, B1 => A_signal(38), 
                           B2 => n145, ZN => n250);
   U110 : AOI22_X1 port map( A1 => A_neg(17), A2 => n152, B1 => A_signal(17), 
                           B2 => n143, ZN => n204);
   U111 : NAND2_X1 port map( A1 => n228, A2 => n227, ZN => Y(28));
   U112 : AOI22_X1 port map( A1 => A_neg(28), A2 => n153, B1 => A_signal(28), 
                           B2 => n144, ZN => n228);
   U113 : AOI222_X1 port map( A1 => A_shifted(28), A2 => n179, B1 => 
                           zeroSignal(28), B2 => n170, C1 => A_neg_shifted(28),
                           C2 => n164, ZN => n227);
   U114 : NAND2_X1 port map( A1 => n256, A2 => n255, ZN => Y(40));
   U115 : AOI222_X1 port map( A1 => A_shifted(40), A2 => n181, B1 => 
                           zeroSignal(40), B2 => n171, C1 => A_neg_shifted(40),
                           C2 => n163, ZN => n255);
   U116 : AOI22_X1 port map( A1 => A_neg(40), A2 => n154, B1 => A_signal(40), 
                           B2 => n145, ZN => n256);
   U117 : NAND2_X1 port map( A1 => n258, A2 => n257, ZN => Y(41));
   U118 : AOI222_X1 port map( A1 => A_shifted(41), A2 => n181, B1 => 
                           zeroSignal(41), B2 => n171, C1 => A_neg_shifted(41),
                           C2 => n163, ZN => n257);
   U119 : AOI22_X1 port map( A1 => A_neg(41), A2 => n154, B1 => A_signal(41), 
                           B2 => n145, ZN => n258);
   U120 : NAND2_X1 port map( A1 => n260, A2 => n259, ZN => Y(42));
   U121 : AOI222_X1 port map( A1 => A_shifted(42), A2 => n181, B1 => 
                           zeroSignal(42), B2 => n172, C1 => A_neg_shifted(42),
                           C2 => n163, ZN => n259);
   U122 : AOI22_X1 port map( A1 => A_neg(42), A2 => n155, B1 => A_signal(42), 
                           B2 => n146, ZN => n260);
   U123 : NAND2_X1 port map( A1 => n212, A2 => n211, ZN => Y(20));
   U124 : AOI222_X1 port map( A1 => A_shifted(20), A2 => n179, B1 => 
                           zeroSignal(20), B2 => n170, C1 => A_neg_shifted(20),
                           C2 => n165, ZN => n211);
   U125 : AOI22_X1 port map( A1 => A_neg(20), A2 => n153, B1 => A_signal(20), 
                           B2 => n144, ZN => n212);
   U126 : NAND2_X1 port map( A1 => n216, A2 => n215, ZN => Y(22));
   U127 : AOI222_X1 port map( A1 => A_shifted(22), A2 => n179, B1 => 
                           zeroSignal(22), B2 => n170, C1 => A_neg_shifted(22),
                           C2 => n165, ZN => n215);
   U128 : AOI22_X1 port map( A1 => A_neg(22), A2 => n153, B1 => A_signal(22), 
                           B2 => n144, ZN => n216);
   U129 : NAND2_X1 port map( A1 => n252, A2 => n251, ZN => Y(39));
   U130 : AOI22_X1 port map( A1 => A_neg(39), A2 => n154, B1 => A_signal(39), 
                           B2 => n145, ZN => n252);
   U131 : AOI222_X1 port map( A1 => A_shifted(39), A2 => n180, B1 => 
                           zeroSignal(39), B2 => n171, C1 => A_neg_shifted(39),
                           C2 => n163, ZN => n251);
   U132 : NAND2_X1 port map( A1 => n278, A2 => n277, ZN => Y(50));
   U133 : AOI222_X1 port map( A1 => A_shifted(50), A2 => n182, B1 => 
                           zeroSignal(50), B2 => n172, C1 => A_neg_shifted(50),
                           C2 => n162, ZN => n277);
   U134 : AOI22_X1 port map( A1 => A_neg(50), A2 => n155, B1 => A_signal(50), 
                           B2 => n146, ZN => n278);
   U135 : NAND2_X1 port map( A1 => n262, A2 => n261, ZN => Y(43));
   U136 : AOI222_X1 port map( A1 => A_shifted(43), A2 => n181, B1 => 
                           zeroSignal(43), B2 => n172, C1 => A_neg_shifted(43),
                           C2 => n163, ZN => n261);
   U137 : AOI22_X1 port map( A1 => A_neg(43), A2 => n155, B1 => A_signal(43), 
                           B2 => n146, ZN => n262);
   U138 : NAND2_X1 port map( A1 => n274, A2 => n273, ZN => Y(49));
   U139 : AOI22_X1 port map( A1 => A_neg(49), A2 => n155, B1 => A_signal(49), 
                           B2 => n146, ZN => n274);
   U140 : AOI222_X1 port map( A1 => A_shifted(49), A2 => n181, B1 => 
                           zeroSignal(49), B2 => n172, C1 => A_neg_shifted(49),
                           C2 => n162, ZN => n273);
   U141 : NAND2_X1 port map( A1 => n206, A2 => n205, ZN => Y(18));
   U142 : AOI22_X1 port map( A1 => A_neg(18), A2 => n152, B1 => A_signal(18), 
                           B2 => n143, ZN => n206);
   U143 : AOI222_X1 port map( A1 => A_shifted(18), A2 => n178, B1 => 
                           zeroSignal(18), B2 => n169, C1 => A_neg_shifted(18),
                           C2 => n165, ZN => n205);
   U144 : NAND2_X1 port map( A1 => n214, A2 => n213, ZN => Y(21));
   U145 : AOI22_X1 port map( A1 => A_neg(21), A2 => n153, B1 => A_signal(21), 
                           B2 => n144, ZN => n214);
   U146 : AOI222_X1 port map( A1 => A_shifted(21), A2 => n179, B1 => 
                           zeroSignal(21), B2 => n170, C1 => A_neg_shifted(21),
                           C2 => n165, ZN => n213);
   U147 : NAND2_X1 port map( A1 => n264, A2 => n263, ZN => Y(44));
   U148 : AOI222_X1 port map( A1 => A_shifted(44), A2 => n181, B1 => 
                           zeroSignal(44), B2 => n172, C1 => A_neg_shifted(44),
                           C2 => n163, ZN => n263);
   U149 : AOI22_X1 port map( A1 => A_neg(44), A2 => n155, B1 => A_signal(44), 
                           B2 => n146, ZN => n264);
   U150 : NAND2_X1 port map( A1 => n280, A2 => n279, ZN => Y(51));
   U151 : AOI22_X1 port map( A1 => A_neg(51), A2 => n155, B1 => A_signal(51), 
                           B2 => n146, ZN => n280);
   U152 : AOI222_X1 port map( A1 => A_shifted(51), A2 => n182, B1 => 
                           zeroSignal(51), B2 => n172, C1 => A_neg_shifted(51),
                           C2 => n162, ZN => n279);
   U153 : NAND2_X1 port map( A1 => n266, A2 => n265, ZN => Y(45));
   U154 : AOI222_X1 port map( A1 => A_shifted(45), A2 => n181, B1 => 
                           zeroSignal(45), B2 => n172, C1 => A_neg_shifted(45),
                           C2 => n163, ZN => n265);
   U155 : AOI22_X1 port map( A1 => A_neg(45), A2 => n155, B1 => A_signal(45), 
                           B2 => n146, ZN => n266);
   U156 : NAND2_X1 port map( A1 => n268, A2 => n267, ZN => Y(46));
   U157 : AOI222_X1 port map( A1 => A_shifted(46), A2 => n181, B1 => 
                           zeroSignal(46), B2 => n172, C1 => A_neg_shifted(46),
                           C2 => n162, ZN => n267);
   U158 : AOI22_X1 port map( A1 => A_neg(46), A2 => n155, B1 => A_signal(46), 
                           B2 => n146, ZN => n268);
   U159 : NAND2_X1 port map( A1 => n208, A2 => n207, ZN => Y(19));
   U160 : AOI22_X1 port map( A1 => A_neg(19), A2 => n152, B1 => A_signal(19), 
                           B2 => n143, ZN => n208);
   U161 : AOI222_X1 port map( A1 => A_shifted(19), A2 => n178, B1 => 
                           zeroSignal(19), B2 => n169, C1 => A_neg_shifted(19),
                           C2 => n165, ZN => n207);
   U162 : NAND2_X1 port map( A1 => n270, A2 => n269, ZN => Y(47));
   U163 : AOI222_X1 port map( A1 => A_shifted(47), A2 => n181, B1 => 
                           zeroSignal(47), B2 => n172, C1 => A_neg_shifted(47),
                           C2 => n162, ZN => n269);
   U164 : AOI22_X1 port map( A1 => A_neg(47), A2 => n155, B1 => A_signal(47), 
                           B2 => n146, ZN => n270);
   U165 : NAND2_X1 port map( A1 => n306, A2 => n305, ZN => Y(63));
   U166 : AOI222_X1 port map( A1 => A_shifted(63), A2 => n183, B1 => 
                           zeroSignal(63), B2 => n173, C1 => A_neg_shifted(63),
                           C2 => n161, ZN => n305);
   U167 : AOI22_X1 port map( A1 => A_neg(63), A2 => n156, B1 => A_signal(63), 
                           B2 => n147, ZN => n306);
   U168 : NAND2_X1 port map( A1 => n304, A2 => n303, ZN => Y(62));
   U169 : AOI222_X1 port map( A1 => A_shifted(62), A2 => n183, B1 => 
                           zeroSignal(62), B2 => n173, C1 => A_neg_shifted(62),
                           C2 => n161, ZN => n303);
   U170 : AOI22_X1 port map( A1 => A_neg(62), A2 => n156, B1 => A_signal(62), 
                           B2 => n147, ZN => n304);
   U171 : NAND2_X1 port map( A1 => n302, A2 => n301, ZN => Y(61));
   U172 : AOI222_X1 port map( A1 => A_shifted(61), A2 => n183, B1 => 
                           zeroSignal(61), B2 => n173, C1 => A_neg_shifted(61),
                           C2 => n161, ZN => n301);
   U173 : AOI22_X1 port map( A1 => A_neg(61), A2 => n156, B1 => A_signal(61), 
                           B2 => n147, ZN => n302);
   U174 : NAND2_X1 port map( A1 => n284, A2 => n283, ZN => Y(53));
   U175 : AOI22_X1 port map( A1 => A_neg(53), A2 => n156, B1 => A_signal(53), 
                           B2 => n147, ZN => n284);
   U176 : NAND2_X1 port map( A1 => n288, A2 => n287, ZN => Y(55));
   U177 : AOI222_X1 port map( A1 => A_shifted(55), A2 => n182, B1 => 
                           zeroSignal(55), B2 => n173, C1 => A_neg_shifted(55),
                           C2 => n162, ZN => n287);
   U178 : NAND2_X1 port map( A1 => n286, A2 => n285, ZN => Y(54));
   U179 : AOI222_X1 port map( A1 => A_shifted(54), A2 => n182, B1 => 
                           zeroSignal(54), B2 => n173, C1 => A_neg_shifted(54),
                           C2 => n162, ZN => n285);
   U180 : AOI22_X1 port map( A1 => A_neg(54), A2 => n156, B1 => A_signal(54), 
                           B2 => n147, ZN => n286);
   U181 : NAND2_X1 port map( A1 => n282, A2 => n281, ZN => Y(52));
   U182 : AOI222_X1 port map( A1 => A_shifted(52), A2 => n182, B1 => 
                           zeroSignal(52), B2 => n172, C1 => A_neg_shifted(52),
                           C2 => n162, ZN => n281);
   U183 : NAND2_X1 port map( A1 => n290, A2 => n289, ZN => Y(56));
   U184 : AOI22_X1 port map( A1 => A_neg(56), A2 => n156, B1 => A_signal(56), 
                           B2 => n147, ZN => n290);
   U185 : NAND2_X1 port map( A1 => n292, A2 => n291, ZN => Y(57));
   U186 : AOI222_X1 port map( A1 => A_shifted(57), A2 => n182, B1 => 
                           zeroSignal(57), B2 => n173, C1 => A_neg_shifted(57),
                           C2 => n161, ZN => n291);
   U187 : AOI22_X1 port map( A1 => A_neg(57), A2 => n156, B1 => A_signal(57), 
                           B2 => n147, ZN => n292);
   U188 : NAND2_X1 port map( A1 => n294, A2 => n293, ZN => Y(58));
   U189 : AOI222_X1 port map( A1 => A_shifted(58), A2 => n182, B1 => 
                           zeroSignal(58), B2 => n173, C1 => A_neg_shifted(58),
                           C2 => n161, ZN => n293);
   U190 : AOI22_X1 port map( A1 => A_neg(58), A2 => n156, B1 => A_signal(58), 
                           B2 => n147, ZN => n294);
   U191 : NAND2_X1 port map( A1 => n296, A2 => n295, ZN => Y(59));
   U192 : AOI222_X1 port map( A1 => A_shifted(59), A2 => n182, B1 => 
                           zeroSignal(59), B2 => n173, C1 => A_neg_shifted(59),
                           C2 => n161, ZN => n295);
   U193 : AOI22_X1 port map( A1 => A_neg(59), A2 => n156, B1 => A_signal(59), 
                           B2 => n147, ZN => n296);
   U194 : NAND2_X1 port map( A1 => n300, A2 => n299, ZN => Y(60));
   U195 : AOI222_X1 port map( A1 => A_shifted(60), A2 => n183, B1 => 
                           zeroSignal(60), B2 => n173, C1 => A_neg_shifted(60),
                           C2 => n161, ZN => n299);
   U196 : AOI22_X1 port map( A1 => A_neg(60), A2 => n156, B1 => A_signal(60), 
                           B2 => n147, ZN => n300);
   U197 : NAND2_X1 port map( A1 => n188, A2 => n187, ZN => Y(0));
   U198 : AOI22_X1 port map( A1 => A_neg(0), A2 => n152, B1 => A_signal(0), B2 
                           => n143, ZN => n188);
   U199 : AOI222_X1 port map( A1 => A_shifted(0), A2 => n178, B1 => 
                           zeroSignal(0), B2 => n169, C1 => A_neg_shifted(0), 
                           C2 => n166, ZN => n187);
   U200 : NAND2_X1 port map( A1 => n210, A2 => n209, ZN => Y(1));
   U201 : AOI22_X1 port map( A1 => A_neg(1), A2 => n152, B1 => A_signal(1), B2 
                           => n143, ZN => n210);
   U202 : AOI222_X1 port map( A1 => A_shifted(1), A2 => n179, B1 => 
                           zeroSignal(1), B2 => n169, C1 => A_neg_shifted(1), 
                           C2 => n165, ZN => n209);
   U203 : NAND2_X1 port map( A1 => n232, A2 => n231, ZN => Y(2));
   U204 : AOI22_X1 port map( A1 => A_neg(2), A2 => n153, B1 => A_signal(2), B2 
                           => n144, ZN => n232);
   U205 : AOI222_X1 port map( A1 => A_shifted(2), A2 => n180, B1 => 
                           zeroSignal(2), B2 => n170, C1 => A_neg_shifted(2), 
                           C2 => n164, ZN => n231);
   U206 : NAND2_X1 port map( A1 => n254, A2 => n253, ZN => Y(3));
   U207 : AOI22_X1 port map( A1 => A_neg(3), A2 => n154, B1 => A_signal(3), B2 
                           => n145, ZN => n254);
   U208 : AOI222_X1 port map( A1 => A_shifted(3), A2 => n181, B1 => 
                           zeroSignal(3), B2 => n171, C1 => A_neg_shifted(3), 
                           C2 => n163, ZN => n253);
   U209 : NAND2_X1 port map( A1 => n276, A2 => n275, ZN => Y(4));
   U210 : AOI22_X1 port map( A1 => A_neg(4), A2 => n155, B1 => A_signal(4), B2 
                           => n146, ZN => n276);
   U211 : AOI222_X1 port map( A1 => A_shifted(4), A2 => n182, B1 => 
                           zeroSignal(4), B2 => n172, C1 => A_neg_shifted(4), 
                           C2 => n162, ZN => n275);
   U212 : NAND2_X1 port map( A1 => n298, A2 => n297, ZN => Y(5));
   U213 : AOI22_X1 port map( A1 => A_neg(5), A2 => n156, B1 => A_signal(5), B2 
                           => n147, ZN => n298);
   U214 : AOI222_X1 port map( A1 => A_shifted(5), A2 => n183, B1 => 
                           zeroSignal(5), B2 => n173, C1 => A_neg_shifted(5), 
                           C2 => n161, ZN => n297);
   U215 : NAND2_X1 port map( A1 => n308, A2 => n307, ZN => Y(6));
   U216 : AOI22_X1 port map( A1 => A_neg(6), A2 => n157, B1 => A_signal(6), B2 
                           => n148, ZN => n308);
   U217 : AOI222_X1 port map( A1 => A_shifted(6), A2 => n183, B1 => 
                           zeroSignal(6), B2 => n174, C1 => A_neg_shifted(6), 
                           C2 => n161, ZN => n307);
   U218 : NAND2_X1 port map( A1 => n310, A2 => n309, ZN => Y(7));
   U219 : AOI22_X1 port map( A1 => A_neg(7), A2 => n157, B1 => A_signal(7), B2 
                           => n148, ZN => n310);
   U220 : AOI222_X1 port map( A1 => A_shifted(7), A2 => n183, B1 => 
                           zeroSignal(7), B2 => n174, C1 => A_neg_shifted(7), 
                           C2 => n161, ZN => n309);
   U221 : NAND2_X1 port map( A1 => n312, A2 => n311, ZN => Y(8));
   U222 : AOI22_X1 port map( A1 => A_neg(8), A2 => n157, B1 => A_signal(8), B2 
                           => n148, ZN => n312);
   U223 : AOI222_X1 port map( A1 => A_shifted(8), A2 => n183, B1 => 
                           zeroSignal(8), B2 => n174, C1 => A_neg_shifted(8), 
                           C2 => n161, ZN => n311);
   U224 : NAND2_X1 port map( A1 => n317, A2 => n316, ZN => Y(9));
   U225 : AOI22_X1 port map( A1 => A_neg(9), A2 => n157, B1 => A_signal(9), B2 
                           => n148, ZN => n317);
   U226 : AOI222_X1 port map( A1 => A_shifted(9), A2 => n183, B1 => 
                           zeroSignal(9), B2 => n174, C1 => A_neg_shifted(9), 
                           C2 => n161, ZN => n316);
   U227 : AOI222_X1 port map( A1 => A_shifted(11), A2 => n178, B1 => 
                           zeroSignal(11), B2 => n169, C1 => A_neg_shifted(11),
                           C2 => n166, ZN => n191);
   U228 : AOI22_X1 port map( A1 => A_neg(10), A2 => n152, B1 => A_signal(10), 
                           B2 => n143, ZN => n190);
   U229 : AOI222_X1 port map( A1 => A_shifted(17), A2 => n178, B1 => 
                           zeroSignal(17), B2 => n169, C1 => A_neg_shifted(17),
                           C2 => n165, ZN => n203);
   U230 : AOI22_X1 port map( A1 => A_neg(16), A2 => n152, B1 => A_signal(16), 
                           B2 => n143, ZN => n202);
   U231 : NAND2_X1 port map( A1 => n204, A2 => n203, ZN => Y(17));
   U232 : AOI222_X1 port map( A1 => A_shifted(16), A2 => n178, B1 => 
                           zeroSignal(16), B2 => n169, C1 => A_neg_shifted(16),
                           C2 => n165, ZN => n201);
   U233 : AOI22_X1 port map( A1 => A_neg(15), A2 => n152, B1 => A_signal(15), 
                           B2 => n143, ZN => n200);
   U234 : NAND2_X1 port map( A1 => n202, A2 => n201, ZN => Y(16));
   U235 : NAND2_X1 port map( A1 => n200, A2 => n199, ZN => Y(15));
   U236 : AOI222_X1 port map( A1 => A_shifted(14), A2 => n178, B1 => 
                           zeroSignal(14), B2 => n169, C1 => A_neg_shifted(14),
                           C2 => n165, ZN => n197);
   U237 : AOI22_X1 port map( A1 => A_neg(13), A2 => n152, B1 => A_signal(13), 
                           B2 => n143, ZN => n196);
   U238 : NAND2_X1 port map( A1 => n198, A2 => n197, ZN => Y(14));
   U239 : NAND2_X1 port map( A1 => n196, A2 => n195, ZN => Y(13));
   U240 : AOI222_X1 port map( A1 => A_shifted(56), A2 => n182, B1 => 
                           zeroSignal(56), B2 => n173, C1 => A_neg_shifted(56),
                           C2 => n162, ZN => n289);
   U241 : AOI22_X1 port map( A1 => A_neg(55), A2 => n156, B1 => A_signal(55), 
                           B2 => n147, ZN => n288);
   U242 : AOI222_X1 port map( A1 => A_shifted(53), A2 => n182, B1 => 
                           zeroSignal(53), B2 => n173, C1 => A_neg_shifted(53),
                           C2 => n162, ZN => n283);
   U243 : AOI22_X1 port map( A1 => A_neg(52), A2 => n155, B1 => A_signal(52), 
                           B2 => n146, ZN => n282);

end SYN_BEHAVIORAL_2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity MUX51_MuxNbit64_10 is

   port( zeroSignal, A_signal, A_neg, A_shifted, A_neg_shifted : in 
         std_logic_vector (63 downto 0);  Sel : in std_logic_vector (2 downto 
         0);  Y : out std_logic_vector (63 downto 0));

end MUX51_MuxNbit64_10;

architecture SYN_BEHAVIORAL_2 of MUX51_MuxNbit64_10 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, 
      n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, 
      n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, 
      n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, 
      n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, 
      n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, 
      n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, 
      n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, 
      n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, 
      n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, 
      n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, 
      n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, 
      n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, 
      n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, 
      n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, 
      n320 : std_logic;

begin
   
   U1 : AND3_X1 port map( A1 => n319, A2 => n320, A3 => Sel(2), ZN => n141);
   U2 : BUF_X1 port map( A => n141, Z => n166);
   U3 : BUF_X1 port map( A => n159, Z => n158);
   U4 : BUF_X1 port map( A => n185, Z => n184);
   U5 : BUF_X1 port map( A => n150, Z => n149);
   U6 : BUF_X1 port map( A => n141, Z => n167);
   U7 : BUF_X1 port map( A => n185, Z => n183);
   U8 : BUF_X1 port map( A => n159, Z => n157);
   U9 : BUF_X1 port map( A => n150, Z => n148);
   U10 : BUF_X1 port map( A => n176, Z => n175);
   U11 : BUF_X1 port map( A => n176, Z => n174);
   U12 : BUF_X1 port map( A => n158, Z => n151);
   U13 : BUF_X1 port map( A => n149, Z => n142);
   U14 : BUF_X1 port map( A => n184, Z => n177);
   U15 : BUF_X1 port map( A => n166, Z => n164);
   U16 : BUF_X1 port map( A => n184, Z => n178);
   U17 : BUF_X1 port map( A => n158, Z => n152);
   U18 : BUF_X1 port map( A => n149, Z => n143);
   U19 : BUF_X1 port map( A => n166, Z => n163);
   U20 : BUF_X1 port map( A => n184, Z => n179);
   U21 : BUF_X1 port map( A => n158, Z => n153);
   U22 : BUF_X1 port map( A => n149, Z => n144);
   U23 : BUF_X1 port map( A => n167, Z => n162);
   U24 : BUF_X1 port map( A => n183, Z => n180);
   U25 : BUF_X1 port map( A => n157, Z => n154);
   U26 : BUF_X1 port map( A => n148, Z => n145);
   U27 : BUF_X1 port map( A => n167, Z => n161);
   U28 : BUF_X1 port map( A => n183, Z => n181);
   U29 : BUF_X1 port map( A => n157, Z => n155);
   U30 : BUF_X1 port map( A => n148, Z => n146);
   U31 : BUF_X1 port map( A => n167, Z => n160);
   U32 : BUF_X1 port map( A => n183, Z => n182);
   U33 : BUF_X1 port map( A => n175, Z => n169);
   U34 : BUF_X1 port map( A => n175, Z => n170);
   U35 : BUF_X1 port map( A => n174, Z => n171);
   U36 : BUF_X1 port map( A => n175, Z => n168);
   U37 : BUF_X1 port map( A => n174, Z => n172);
   U38 : BUF_X1 port map( A => n166, Z => n165);
   U39 : BUF_X1 port map( A => n157, Z => n156);
   U40 : BUF_X1 port map( A => n148, Z => n147);
   U41 : BUF_X1 port map( A => n174, Z => n173);
   U42 : BUF_X1 port map( A => n314, Z => n159);
   U43 : NOR3_X1 port map( A1 => Sel(0), A2 => Sel(2), A3 => n320, ZN => n314);
   U44 : INV_X1 port map( A => Sel(1), ZN => n320);
   U45 : BUF_X1 port map( A => n313, Z => n150);
   U46 : NOR3_X1 port map( A1 => Sel(1), A2 => Sel(2), A3 => n319, ZN => n313);
   U47 : INV_X1 port map( A => Sel(0), ZN => n319);
   U48 : BUF_X1 port map( A => n316, Z => n185);
   U49 : NOR3_X1 port map( A1 => n319, A2 => Sel(2), A3 => n320, ZN => n316);
   U50 : BUF_X1 port map( A => n315, Z => n176);
   U51 : NOR2_X1 port map( A1 => n165, A2 => n186, ZN => n315);
   U52 : AOI21_X1 port map( B1 => n319, B2 => n320, A => Sel(2), ZN => n186);
   U53 : NAND2_X1 port map( A1 => n196, A2 => n195, ZN => Y(13));
   U54 : AOI22_X1 port map( A1 => A_neg(13), A2 => n151, B1 => A_signal(13), B2
                           => n142, ZN => n196);
   U55 : NAND2_X1 port map( A1 => n194, A2 => n193, ZN => Y(12));
   U56 : AOI222_X1 port map( A1 => A_shifted(12), A2 => n177, B1 => 
                           zeroSignal(12), B2 => n168, C1 => A_neg_shifted(12),
                           C2 => n165, ZN => n193);
   U57 : NAND2_X1 port map( A1 => n198, A2 => n197, ZN => Y(14));
   U58 : AOI222_X1 port map( A1 => A_shifted(14), A2 => n177, B1 => 
                           zeroSignal(14), B2 => n168, C1 => A_neg_shifted(14),
                           C2 => n164, ZN => n197);
   U59 : AOI22_X1 port map( A1 => A_neg(14), A2 => n151, B1 => A_signal(14), B2
                           => n142, ZN => n198);
   U60 : NAND2_X1 port map( A1 => n260, A2 => n259, ZN => Y(42));
   U61 : AOI222_X1 port map( A1 => A_shifted(42), A2 => n180, B1 => 
                           zeroSignal(42), B2 => n171, C1 => A_neg_shifted(42),
                           C2 => n162, ZN => n259);
   U62 : AOI22_X1 port map( A1 => A_neg(42), A2 => n154, B1 => A_signal(42), B2
                           => n145, ZN => n260);
   U63 : AOI222_X1 port map( A1 => A_shifted(15), A2 => n177, B1 => 
                           zeroSignal(15), B2 => n168, C1 => A_neg_shifted(15),
                           C2 => n164, ZN => n199);
   U64 : AOI222_X1 port map( A1 => A_shifted(16), A2 => n177, B1 => 
                           zeroSignal(16), B2 => n168, C1 => A_neg_shifted(16),
                           C2 => n164, ZN => n201);
   U65 : AOI22_X1 port map( A1 => A_neg(16), A2 => n151, B1 => A_signal(16), B2
                           => n142, ZN => n202);
   U66 : NAND2_X1 port map( A1 => n272, A2 => n271, ZN => Y(48));
   U67 : AOI222_X1 port map( A1 => A_shifted(48), A2 => n180, B1 => 
                           zeroSignal(48), B2 => n171, C1 => A_neg_shifted(48),
                           C2 => n161, ZN => n271);
   U68 : AOI22_X1 port map( A1 => A_neg(48), A2 => n154, B1 => A_signal(48), B2
                           => n145, ZN => n272);
   U69 : AOI222_X1 port map( A1 => A_shifted(17), A2 => n177, B1 => 
                           zeroSignal(17), B2 => n168, C1 => A_neg_shifted(17),
                           C2 => n164, ZN => n203);
   U70 : NAND2_X1 port map( A1 => n274, A2 => n273, ZN => Y(49));
   U71 : AOI222_X1 port map( A1 => A_shifted(49), A2 => n180, B1 => 
                           zeroSignal(49), B2 => n171, C1 => A_neg_shifted(49),
                           C2 => n161, ZN => n273);
   U72 : AOI22_X1 port map( A1 => A_neg(49), A2 => n154, B1 => A_signal(49), B2
                           => n145, ZN => n274);
   U73 : NAND2_X1 port map( A1 => n278, A2 => n277, ZN => Y(50));
   U74 : AOI22_X1 port map( A1 => A_neg(50), A2 => n154, B1 => A_signal(50), B2
                           => n145, ZN => n278);
   U75 : AOI222_X1 port map( A1 => A_shifted(50), A2 => n181, B1 => 
                           zeroSignal(50), B2 => n171, C1 => A_neg_shifted(50),
                           C2 => n161, ZN => n277);
   U76 : AOI222_X1 port map( A1 => A_shifted(18), A2 => n177, B1 => 
                           zeroSignal(18), B2 => n168, C1 => A_neg_shifted(18),
                           C2 => n164, ZN => n205);
   U77 : NAND2_X1 port map( A1 => n226, A2 => n225, ZN => Y(27));
   U78 : AOI222_X1 port map( A1 => A_shifted(27), A2 => n178, B1 => 
                           zeroSignal(27), B2 => n169, C1 => A_neg_shifted(27),
                           C2 => n163, ZN => n225);
   U79 : AOI22_X1 port map( A1 => A_neg(27), A2 => n152, B1 => A_signal(27), B2
                           => n143, ZN => n226);
   U80 : NAND2_X1 port map( A1 => n222, A2 => n221, ZN => Y(25));
   U81 : AOI222_X1 port map( A1 => A_shifted(25), A2 => n178, B1 => 
                           zeroSignal(25), B2 => n169, C1 => A_neg_shifted(25),
                           C2 => n163, ZN => n221);
   U82 : AOI22_X1 port map( A1 => A_neg(25), A2 => n152, B1 => A_signal(25), B2
                           => n143, ZN => n222);
   U83 : NAND2_X1 port map( A1 => n224, A2 => n223, ZN => Y(26));
   U84 : AOI222_X1 port map( A1 => A_shifted(26), A2 => n178, B1 => 
                           zeroSignal(26), B2 => n169, C1 => A_neg_shifted(26),
                           C2 => n163, ZN => n223);
   U85 : AOI22_X1 port map( A1 => A_neg(26), A2 => n152, B1 => A_signal(26), B2
                           => n143, ZN => n224);
   U86 : NAND2_X1 port map( A1 => n230, A2 => n229, ZN => Y(29));
   U87 : AOI222_X1 port map( A1 => A_shifted(29), A2 => n178, B1 => 
                           zeroSignal(29), B2 => n169, C1 => A_neg_shifted(29),
                           C2 => n163, ZN => n229);
   U88 : AOI22_X1 port map( A1 => A_neg(29), A2 => n152, B1 => A_signal(29), B2
                           => n143, ZN => n230);
   U89 : NAND2_X1 port map( A1 => n228, A2 => n227, ZN => Y(28));
   U90 : AOI222_X1 port map( A1 => A_shifted(28), A2 => n178, B1 => 
                           zeroSignal(28), B2 => n169, C1 => A_neg_shifted(28),
                           C2 => n163, ZN => n227);
   U91 : AOI22_X1 port map( A1 => A_neg(28), A2 => n152, B1 => A_signal(28), B2
                           => n143, ZN => n228);
   U92 : NAND2_X1 port map( A1 => n236, A2 => n235, ZN => Y(31));
   U93 : AOI222_X1 port map( A1 => A_shifted(31), A2 => n179, B1 => 
                           zeroSignal(31), B2 => n170, C1 => A_neg_shifted(31),
                           C2 => n163, ZN => n235);
   U94 : AOI22_X1 port map( A1 => A_neg(31), A2 => n153, B1 => A_signal(31), B2
                           => n144, ZN => n236);
   U95 : NAND2_X1 port map( A1 => n238, A2 => n237, ZN => Y(32));
   U96 : AOI222_X1 port map( A1 => A_shifted(32), A2 => n179, B1 => 
                           zeroSignal(32), B2 => n170, C1 => A_neg_shifted(32),
                           C2 => n163, ZN => n237);
   U97 : AOI22_X1 port map( A1 => A_neg(32), A2 => n153, B1 => A_signal(32), B2
                           => n144, ZN => n238);
   U98 : NAND2_X1 port map( A1 => n242, A2 => n241, ZN => Y(34));
   U99 : AOI222_X1 port map( A1 => A_shifted(34), A2 => n179, B1 => 
                           zeroSignal(34), B2 => n170, C1 => A_neg_shifted(34),
                           C2 => n163, ZN => n241);
   U100 : AOI22_X1 port map( A1 => A_neg(34), A2 => n153, B1 => A_signal(34), 
                           B2 => n144, ZN => n242);
   U101 : NAND2_X1 port map( A1 => n240, A2 => n239, ZN => Y(33));
   U102 : AOI222_X1 port map( A1 => A_shifted(33), A2 => n179, B1 => 
                           zeroSignal(33), B2 => n170, C1 => A_neg_shifted(33),
                           C2 => n163, ZN => n239);
   U103 : AOI22_X1 port map( A1 => A_neg(33), A2 => n153, B1 => A_signal(33), 
                           B2 => n144, ZN => n240);
   U104 : NAND2_X1 port map( A1 => n244, A2 => n243, ZN => Y(35));
   U105 : AOI222_X1 port map( A1 => A_shifted(35), A2 => n179, B1 => 
                           zeroSignal(35), B2 => n170, C1 => A_neg_shifted(35),
                           C2 => n162, ZN => n243);
   U106 : AOI22_X1 port map( A1 => A_neg(35), A2 => n153, B1 => A_signal(35), 
                           B2 => n144, ZN => n244);
   U107 : NAND2_X1 port map( A1 => n246, A2 => n245, ZN => Y(36));
   U108 : AOI222_X1 port map( A1 => A_shifted(36), A2 => n179, B1 => 
                           zeroSignal(36), B2 => n170, C1 => A_neg_shifted(36),
                           C2 => n162, ZN => n245);
   U109 : AOI22_X1 port map( A1 => A_neg(36), A2 => n153, B1 => A_signal(36), 
                           B2 => n144, ZN => n246);
   U110 : NAND2_X1 port map( A1 => n248, A2 => n247, ZN => Y(37));
   U111 : AOI222_X1 port map( A1 => A_shifted(37), A2 => n179, B1 => 
                           zeroSignal(37), B2 => n170, C1 => A_neg_shifted(37),
                           C2 => n162, ZN => n247);
   U112 : AOI22_X1 port map( A1 => A_neg(37), A2 => n153, B1 => A_signal(37), 
                           B2 => n144, ZN => n248);
   U113 : NAND2_X1 port map( A1 => n250, A2 => n249, ZN => Y(38));
   U114 : AOI222_X1 port map( A1 => A_shifted(38), A2 => n179, B1 => 
                           zeroSignal(38), B2 => n170, C1 => A_neg_shifted(38),
                           C2 => n162, ZN => n249);
   U115 : AOI22_X1 port map( A1 => A_neg(38), A2 => n153, B1 => A_signal(38), 
                           B2 => n144, ZN => n250);
   U116 : NAND2_X1 port map( A1 => n252, A2 => n251, ZN => Y(39));
   U117 : AOI222_X1 port map( A1 => A_shifted(39), A2 => n179, B1 => 
                           zeroSignal(39), B2 => n170, C1 => A_neg_shifted(39),
                           C2 => n162, ZN => n251);
   U118 : AOI22_X1 port map( A1 => A_neg(39), A2 => n153, B1 => A_signal(39), 
                           B2 => n144, ZN => n252);
   U119 : NAND2_X1 port map( A1 => n256, A2 => n255, ZN => Y(40));
   U120 : AOI222_X1 port map( A1 => A_shifted(40), A2 => n180, B1 => 
                           zeroSignal(40), B2 => n170, C1 => A_neg_shifted(40),
                           C2 => n162, ZN => n255);
   U121 : AOI22_X1 port map( A1 => A_neg(40), A2 => n153, B1 => A_signal(40), 
                           B2 => n144, ZN => n256);
   U122 : AOI22_X1 port map( A1 => A_neg(19), A2 => n151, B1 => A_signal(19), 
                           B2 => n142, ZN => n208);
   U123 : AOI222_X1 port map( A1 => A_shifted(19), A2 => n177, B1 => 
                           zeroSignal(19), B2 => n168, C1 => A_neg_shifted(19),
                           C2 => n164, ZN => n207);
   U124 : NAND2_X1 port map( A1 => n234, A2 => n233, ZN => Y(30));
   U125 : AOI22_X1 port map( A1 => A_neg(30), A2 => n152, B1 => A_signal(30), 
                           B2 => n143, ZN => n234);
   U126 : AOI222_X1 port map( A1 => A_shifted(30), A2 => n179, B1 => 
                           zeroSignal(30), B2 => n169, C1 => A_neg_shifted(30),
                           C2 => n163, ZN => n233);
   U127 : NAND2_X1 port map( A1 => n262, A2 => n261, ZN => Y(43));
   U128 : AOI222_X1 port map( A1 => A_shifted(43), A2 => n180, B1 => 
                           zeroSignal(43), B2 => n171, C1 => A_neg_shifted(43),
                           C2 => n162, ZN => n261);
   U129 : AOI22_X1 port map( A1 => A_neg(43), A2 => n154, B1 => A_signal(43), 
                           B2 => n145, ZN => n262);
   U130 : NAND2_X1 port map( A1 => n264, A2 => n263, ZN => Y(44));
   U131 : AOI222_X1 port map( A1 => A_shifted(44), A2 => n180, B1 => 
                           zeroSignal(44), B2 => n171, C1 => A_neg_shifted(44),
                           C2 => n162, ZN => n263);
   U132 : AOI22_X1 port map( A1 => A_neg(44), A2 => n154, B1 => A_signal(44), 
                           B2 => n145, ZN => n264);
   U133 : NAND2_X1 port map( A1 => n216, A2 => n215, ZN => Y(22));
   U134 : AOI222_X1 port map( A1 => A_shifted(22), A2 => n178, B1 => 
                           zeroSignal(22), B2 => n169, C1 => A_neg_shifted(22),
                           C2 => n164, ZN => n215);
   U135 : AOI22_X1 port map( A1 => A_neg(22), A2 => n152, B1 => A_signal(22), 
                           B2 => n143, ZN => n216);
   U136 : NAND2_X1 port map( A1 => n220, A2 => n219, ZN => Y(24));
   U137 : AOI222_X1 port map( A1 => A_shifted(24), A2 => n178, B1 => 
                           zeroSignal(24), B2 => n169, C1 => A_neg_shifted(24),
                           C2 => n163, ZN => n219);
   U138 : AOI22_X1 port map( A1 => A_neg(24), A2 => n152, B1 => A_signal(24), 
                           B2 => n143, ZN => n220);
   U139 : NAND2_X1 port map( A1 => n258, A2 => n257, ZN => Y(41));
   U140 : AOI22_X1 port map( A1 => A_neg(41), A2 => n153, B1 => A_signal(41), 
                           B2 => n144, ZN => n258);
   U141 : AOI222_X1 port map( A1 => A_shifted(41), A2 => n180, B1 => 
                           zeroSignal(41), B2 => n170, C1 => A_neg_shifted(41),
                           C2 => n162, ZN => n257);
   U142 : NAND2_X1 port map( A1 => n282, A2 => n281, ZN => Y(52));
   U143 : AOI222_X1 port map( A1 => A_shifted(52), A2 => n181, B1 => 
                           zeroSignal(52), B2 => n171, C1 => A_neg_shifted(52),
                           C2 => n161, ZN => n281);
   U144 : AOI22_X1 port map( A1 => A_neg(52), A2 => n154, B1 => A_signal(52), 
                           B2 => n145, ZN => n282);
   U145 : NAND2_X1 port map( A1 => n266, A2 => n265, ZN => Y(45));
   U146 : AOI222_X1 port map( A1 => A_shifted(45), A2 => n180, B1 => 
                           zeroSignal(45), B2 => n171, C1 => A_neg_shifted(45),
                           C2 => n162, ZN => n265);
   U147 : AOI22_X1 port map( A1 => A_neg(45), A2 => n154, B1 => A_signal(45), 
                           B2 => n145, ZN => n266);
   U148 : NAND2_X1 port map( A1 => n280, A2 => n279, ZN => Y(51));
   U149 : AOI22_X1 port map( A1 => A_neg(51), A2 => n154, B1 => A_signal(51), 
                           B2 => n145, ZN => n280);
   U150 : AOI222_X1 port map( A1 => A_shifted(51), A2 => n181, B1 => 
                           zeroSignal(51), B2 => n171, C1 => A_neg_shifted(51),
                           C2 => n161, ZN => n279);
   U151 : NAND2_X1 port map( A1 => n212, A2 => n211, ZN => Y(20));
   U152 : AOI22_X1 port map( A1 => A_neg(20), A2 => n152, B1 => A_signal(20), 
                           B2 => n143, ZN => n212);
   U153 : AOI222_X1 port map( A1 => A_shifted(20), A2 => n178, B1 => 
                           zeroSignal(20), B2 => n169, C1 => A_neg_shifted(20),
                           C2 => n164, ZN => n211);
   U154 : NAND2_X1 port map( A1 => n218, A2 => n217, ZN => Y(23));
   U155 : AOI22_X1 port map( A1 => A_neg(23), A2 => n152, B1 => A_signal(23), 
                           B2 => n143, ZN => n218);
   U156 : AOI222_X1 port map( A1 => A_shifted(23), A2 => n178, B1 => 
                           zeroSignal(23), B2 => n169, C1 => A_neg_shifted(23),
                           C2 => n164, ZN => n217);
   U157 : NAND2_X1 port map( A1 => n268, A2 => n267, ZN => Y(46));
   U158 : AOI222_X1 port map( A1 => A_shifted(46), A2 => n180, B1 => 
                           zeroSignal(46), B2 => n171, C1 => A_neg_shifted(46),
                           C2 => n161, ZN => n267);
   U159 : AOI22_X1 port map( A1 => A_neg(46), A2 => n154, B1 => A_signal(46), 
                           B2 => n145, ZN => n268);
   U160 : NAND2_X1 port map( A1 => n284, A2 => n283, ZN => Y(53));
   U161 : AOI22_X1 port map( A1 => A_neg(53), A2 => n155, B1 => A_signal(53), 
                           B2 => n146, ZN => n284);
   U162 : AOI222_X1 port map( A1 => A_shifted(53), A2 => n181, B1 => 
                           zeroSignal(53), B2 => n172, C1 => A_neg_shifted(53),
                           C2 => n161, ZN => n283);
   U163 : NAND2_X1 port map( A1 => n270, A2 => n269, ZN => Y(47));
   U164 : AOI222_X1 port map( A1 => A_shifted(47), A2 => n180, B1 => 
                           zeroSignal(47), B2 => n171, C1 => A_neg_shifted(47),
                           C2 => n161, ZN => n269);
   U165 : AOI22_X1 port map( A1 => A_neg(47), A2 => n154, B1 => A_signal(47), 
                           B2 => n145, ZN => n270);
   U166 : NAND2_X1 port map( A1 => n214, A2 => n213, ZN => Y(21));
   U167 : AOI22_X1 port map( A1 => A_neg(21), A2 => n152, B1 => A_signal(21), 
                           B2 => n143, ZN => n214);
   U168 : AOI222_X1 port map( A1 => A_shifted(21), A2 => n178, B1 => 
                           zeroSignal(21), B2 => n169, C1 => A_neg_shifted(21),
                           C2 => n164, ZN => n213);
   U169 : NAND2_X1 port map( A1 => n306, A2 => n305, ZN => Y(63));
   U170 : AOI222_X1 port map( A1 => A_shifted(63), A2 => n182, B1 => 
                           zeroSignal(63), B2 => n172, C1 => A_neg_shifted(63),
                           C2 => n160, ZN => n305);
   U171 : AOI22_X1 port map( A1 => A_neg(63), A2 => n155, B1 => A_signal(63), 
                           B2 => n146, ZN => n306);
   U172 : NAND2_X1 port map( A1 => n288, A2 => n287, ZN => Y(55));
   U173 : AOI22_X1 port map( A1 => A_neg(55), A2 => n155, B1 => A_signal(55), 
                           B2 => n146, ZN => n288);
   U174 : NAND2_X1 port map( A1 => n292, A2 => n291, ZN => Y(57));
   U175 : AOI222_X1 port map( A1 => A_shifted(57), A2 => n181, B1 => 
                           zeroSignal(57), B2 => n172, C1 => A_neg_shifted(57),
                           C2 => n160, ZN => n291);
   U176 : NAND2_X1 port map( A1 => n290, A2 => n289, ZN => Y(56));
   U177 : AOI222_X1 port map( A1 => A_shifted(56), A2 => n181, B1 => 
                           zeroSignal(56), B2 => n172, C1 => A_neg_shifted(56),
                           C2 => n161, ZN => n289);
   U178 : AOI22_X1 port map( A1 => A_neg(56), A2 => n155, B1 => A_signal(56), 
                           B2 => n146, ZN => n290);
   U179 : NAND2_X1 port map( A1 => n286, A2 => n285, ZN => Y(54));
   U180 : AOI222_X1 port map( A1 => A_shifted(54), A2 => n181, B1 => 
                           zeroSignal(54), B2 => n172, C1 => A_neg_shifted(54),
                           C2 => n161, ZN => n285);
   U181 : NAND2_X1 port map( A1 => n294, A2 => n293, ZN => Y(58));
   U182 : AOI22_X1 port map( A1 => A_neg(58), A2 => n155, B1 => A_signal(58), 
                           B2 => n146, ZN => n294);
   U183 : NAND2_X1 port map( A1 => n296, A2 => n295, ZN => Y(59));
   U184 : AOI222_X1 port map( A1 => A_shifted(59), A2 => n181, B1 => 
                           zeroSignal(59), B2 => n172, C1 => A_neg_shifted(59),
                           C2 => n160, ZN => n295);
   U185 : AOI22_X1 port map( A1 => A_neg(59), A2 => n155, B1 => A_signal(59), 
                           B2 => n146, ZN => n296);
   U186 : NAND2_X1 port map( A1 => n304, A2 => n303, ZN => Y(62));
   U187 : AOI222_X1 port map( A1 => A_shifted(62), A2 => n182, B1 => 
                           zeroSignal(62), B2 => n172, C1 => A_neg_shifted(62),
                           C2 => n160, ZN => n303);
   U188 : AOI22_X1 port map( A1 => A_neg(62), A2 => n155, B1 => A_signal(62), 
                           B2 => n146, ZN => n304);
   U189 : NAND2_X1 port map( A1 => n302, A2 => n301, ZN => Y(61));
   U190 : AOI222_X1 port map( A1 => A_shifted(61), A2 => n182, B1 => 
                           zeroSignal(61), B2 => n172, C1 => A_neg_shifted(61),
                           C2 => n160, ZN => n301);
   U191 : AOI22_X1 port map( A1 => A_neg(61), A2 => n155, B1 => A_signal(61), 
                           B2 => n146, ZN => n302);
   U192 : NAND2_X1 port map( A1 => n300, A2 => n299, ZN => Y(60));
   U193 : AOI222_X1 port map( A1 => A_shifted(60), A2 => n182, B1 => 
                           zeroSignal(60), B2 => n172, C1 => A_neg_shifted(60),
                           C2 => n160, ZN => n299);
   U194 : AOI22_X1 port map( A1 => A_neg(60), A2 => n155, B1 => A_signal(60), 
                           B2 => n146, ZN => n300);
   U195 : NAND2_X1 port map( A1 => n188, A2 => n187, ZN => Y(0));
   U196 : AOI22_X1 port map( A1 => A_neg(0), A2 => n151, B1 => A_signal(0), B2 
                           => n142, ZN => n188);
   U197 : AOI222_X1 port map( A1 => A_shifted(0), A2 => n177, B1 => 
                           zeroSignal(0), B2 => n168, C1 => A_neg_shifted(0), 
                           C2 => n165, ZN => n187);
   U198 : NAND2_X1 port map( A1 => n210, A2 => n209, ZN => Y(1));
   U199 : AOI22_X1 port map( A1 => A_neg(1), A2 => n151, B1 => A_signal(1), B2 
                           => n142, ZN => n210);
   U200 : AOI222_X1 port map( A1 => A_shifted(1), A2 => n178, B1 => 
                           zeroSignal(1), B2 => n168, C1 => A_neg_shifted(1), 
                           C2 => n164, ZN => n209);
   U201 : NAND2_X1 port map( A1 => n232, A2 => n231, ZN => Y(2));
   U202 : AOI22_X1 port map( A1 => A_neg(2), A2 => n152, B1 => A_signal(2), B2 
                           => n143, ZN => n232);
   U203 : AOI222_X1 port map( A1 => A_shifted(2), A2 => n179, B1 => 
                           zeroSignal(2), B2 => n169, C1 => A_neg_shifted(2), 
                           C2 => n163, ZN => n231);
   U204 : NAND2_X1 port map( A1 => n254, A2 => n253, ZN => Y(3));
   U205 : AOI22_X1 port map( A1 => A_neg(3), A2 => n153, B1 => A_signal(3), B2 
                           => n144, ZN => n254);
   U206 : AOI222_X1 port map( A1 => A_shifted(3), A2 => n180, B1 => 
                           zeroSignal(3), B2 => n170, C1 => A_neg_shifted(3), 
                           C2 => n162, ZN => n253);
   U207 : NAND2_X1 port map( A1 => n276, A2 => n275, ZN => Y(4));
   U208 : AOI22_X1 port map( A1 => A_neg(4), A2 => n154, B1 => A_signal(4), B2 
                           => n145, ZN => n276);
   U209 : AOI222_X1 port map( A1 => A_shifted(4), A2 => n181, B1 => 
                           zeroSignal(4), B2 => n171, C1 => A_neg_shifted(4), 
                           C2 => n161, ZN => n275);
   U210 : NAND2_X1 port map( A1 => n298, A2 => n297, ZN => Y(5));
   U211 : AOI22_X1 port map( A1 => A_neg(5), A2 => n155, B1 => A_signal(5), B2 
                           => n146, ZN => n298);
   U212 : AOI222_X1 port map( A1 => A_shifted(5), A2 => n182, B1 => 
                           zeroSignal(5), B2 => n172, C1 => A_neg_shifted(5), 
                           C2 => n160, ZN => n297);
   U213 : NAND2_X1 port map( A1 => n308, A2 => n307, ZN => Y(6));
   U214 : AOI22_X1 port map( A1 => A_neg(6), A2 => n156, B1 => A_signal(6), B2 
                           => n147, ZN => n308);
   U215 : AOI222_X1 port map( A1 => A_shifted(6), A2 => n182, B1 => 
                           zeroSignal(6), B2 => n173, C1 => A_neg_shifted(6), 
                           C2 => n160, ZN => n307);
   U216 : NAND2_X1 port map( A1 => n310, A2 => n309, ZN => Y(7));
   U217 : AOI22_X1 port map( A1 => A_neg(7), A2 => n156, B1 => A_signal(7), B2 
                           => n147, ZN => n310);
   U218 : AOI222_X1 port map( A1 => A_shifted(7), A2 => n182, B1 => 
                           zeroSignal(7), B2 => n173, C1 => A_neg_shifted(7), 
                           C2 => n160, ZN => n309);
   U219 : NAND2_X1 port map( A1 => n312, A2 => n311, ZN => Y(8));
   U220 : AOI22_X1 port map( A1 => A_neg(8), A2 => n156, B1 => A_signal(8), B2 
                           => n147, ZN => n312);
   U221 : AOI222_X1 port map( A1 => A_shifted(8), A2 => n182, B1 => 
                           zeroSignal(8), B2 => n173, C1 => A_neg_shifted(8), 
                           C2 => n160, ZN => n311);
   U222 : NAND2_X1 port map( A1 => n318, A2 => n317, ZN => Y(9));
   U223 : AOI22_X1 port map( A1 => A_neg(9), A2 => n156, B1 => A_signal(9), B2 
                           => n147, ZN => n318);
   U224 : AOI222_X1 port map( A1 => A_shifted(9), A2 => n182, B1 => 
                           zeroSignal(9), B2 => n173, C1 => A_neg_shifted(9), 
                           C2 => n160, ZN => n317);
   U225 : NAND2_X1 port map( A1 => n190, A2 => n189, ZN => Y(10));
   U226 : AOI22_X1 port map( A1 => A_neg(10), A2 => n151, B1 => A_signal(10), 
                           B2 => n142, ZN => n190);
   U227 : AOI222_X1 port map( A1 => A_shifted(10), A2 => n177, B1 => 
                           zeroSignal(10), B2 => n168, C1 => A_neg_shifted(10),
                           C2 => n165, ZN => n189);
   U228 : NAND2_X1 port map( A1 => n192, A2 => n191, ZN => Y(11));
   U229 : AOI22_X1 port map( A1 => A_neg(11), A2 => n151, B1 => A_signal(11), 
                           B2 => n142, ZN => n192);
   U230 : AOI222_X1 port map( A1 => A_shifted(11), A2 => n177, B1 => 
                           zeroSignal(11), B2 => n168, C1 => A_neg_shifted(11),
                           C2 => n165, ZN => n191);
   U231 : AOI222_X1 port map( A1 => A_shifted(13), A2 => n177, B1 => 
                           zeroSignal(13), B2 => n168, C1 => A_neg_shifted(13),
                           C2 => n164, ZN => n195);
   U232 : AOI22_X1 port map( A1 => A_neg(12), A2 => n151, B1 => A_signal(12), 
                           B2 => n142, ZN => n194);
   U233 : AOI22_X1 port map( A1 => A_neg(18), A2 => n151, B1 => A_signal(18), 
                           B2 => n142, ZN => n206);
   U234 : NAND2_X1 port map( A1 => n208, A2 => n207, ZN => Y(19));
   U235 : AOI22_X1 port map( A1 => A_neg(17), A2 => n151, B1 => A_signal(17), 
                           B2 => n142, ZN => n204);
   U236 : NAND2_X1 port map( A1 => n206, A2 => n205, ZN => Y(18));
   U237 : NAND2_X1 port map( A1 => n204, A2 => n203, ZN => Y(17));
   U238 : AOI22_X1 port map( A1 => A_neg(15), A2 => n151, B1 => A_signal(15), 
                           B2 => n142, ZN => n200);
   U239 : NAND2_X1 port map( A1 => n202, A2 => n201, ZN => Y(16));
   U240 : NAND2_X1 port map( A1 => n200, A2 => n199, ZN => Y(15));
   U241 : AOI222_X1 port map( A1 => A_shifted(58), A2 => n181, B1 => 
                           zeroSignal(58), B2 => n172, C1 => A_neg_shifted(58),
                           C2 => n160, ZN => n293);
   U242 : AOI22_X1 port map( A1 => A_neg(57), A2 => n155, B1 => A_signal(57), 
                           B2 => n146, ZN => n292);
   U243 : AOI222_X1 port map( A1 => A_shifted(55), A2 => n181, B1 => 
                           zeroSignal(55), B2 => n172, C1 => A_neg_shifted(55),
                           C2 => n161, ZN => n287);
   U244 : AOI22_X1 port map( A1 => A_neg(54), A2 => n155, B1 => A_signal(54), 
                           B2 => n146, ZN => n286);

end SYN_BEHAVIORAL_2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity MUX51_MuxNbit64_9 is

   port( zeroSignal, A_signal, A_neg, A_shifted, A_neg_shifted : in 
         std_logic_vector (63 downto 0);  Sel : in std_logic_vector (2 downto 
         0);  Y : out std_logic_vector (63 downto 0));

end MUX51_MuxNbit64_9;

architecture SYN_BEHAVIORAL_2 of MUX51_MuxNbit64_9 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, 
      n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, 
      n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, 
      n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, 
      n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, 
      n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, 
      n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, 
      n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, 
      n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, 
      n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, 
      n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, 
      n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, 
      n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, 
      n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, 
      n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, 
      n320 : std_logic;

begin
   
   U1 : AND3_X1 port map( A1 => n319, A2 => n320, A3 => Sel(2), ZN => n141);
   U2 : BUF_X1 port map( A => n141, Z => n166);
   U3 : BUF_X1 port map( A => n159, Z => n158);
   U4 : BUF_X1 port map( A => n185, Z => n184);
   U5 : BUF_X1 port map( A => n150, Z => n149);
   U6 : BUF_X1 port map( A => n141, Z => n167);
   U7 : BUF_X1 port map( A => n185, Z => n183);
   U8 : BUF_X1 port map( A => n159, Z => n157);
   U9 : BUF_X1 port map( A => n150, Z => n148);
   U10 : BUF_X1 port map( A => n176, Z => n175);
   U11 : BUF_X1 port map( A => n176, Z => n174);
   U12 : BUF_X1 port map( A => n158, Z => n151);
   U13 : BUF_X1 port map( A => n149, Z => n142);
   U14 : BUF_X1 port map( A => n184, Z => n177);
   U15 : BUF_X1 port map( A => n166, Z => n164);
   U16 : BUF_X1 port map( A => n184, Z => n178);
   U17 : BUF_X1 port map( A => n158, Z => n152);
   U18 : BUF_X1 port map( A => n149, Z => n143);
   U19 : BUF_X1 port map( A => n166, Z => n163);
   U20 : BUF_X1 port map( A => n184, Z => n179);
   U21 : BUF_X1 port map( A => n158, Z => n153);
   U22 : BUF_X1 port map( A => n149, Z => n144);
   U23 : BUF_X1 port map( A => n167, Z => n162);
   U24 : BUF_X1 port map( A => n183, Z => n180);
   U25 : BUF_X1 port map( A => n157, Z => n154);
   U26 : BUF_X1 port map( A => n148, Z => n145);
   U27 : BUF_X1 port map( A => n167, Z => n161);
   U28 : BUF_X1 port map( A => n183, Z => n181);
   U29 : BUF_X1 port map( A => n157, Z => n155);
   U30 : BUF_X1 port map( A => n148, Z => n146);
   U31 : BUF_X1 port map( A => n167, Z => n160);
   U32 : BUF_X1 port map( A => n183, Z => n182);
   U33 : BUF_X1 port map( A => n175, Z => n169);
   U34 : BUF_X1 port map( A => n175, Z => n170);
   U35 : BUF_X1 port map( A => n174, Z => n171);
   U36 : BUF_X1 port map( A => n175, Z => n168);
   U37 : BUF_X1 port map( A => n174, Z => n172);
   U38 : BUF_X1 port map( A => n166, Z => n165);
   U39 : BUF_X1 port map( A => n157, Z => n156);
   U40 : BUF_X1 port map( A => n148, Z => n147);
   U41 : BUF_X1 port map( A => n174, Z => n173);
   U42 : BUF_X1 port map( A => n314, Z => n159);
   U43 : NOR3_X1 port map( A1 => Sel(0), A2 => Sel(2), A3 => n320, ZN => n314);
   U44 : INV_X1 port map( A => Sel(1), ZN => n320);
   U45 : INV_X1 port map( A => Sel(0), ZN => n319);
   U46 : BUF_X1 port map( A => n313, Z => n150);
   U47 : NOR3_X1 port map( A1 => Sel(1), A2 => Sel(2), A3 => n319, ZN => n313);
   U48 : BUF_X1 port map( A => n316, Z => n185);
   U49 : NOR3_X1 port map( A1 => n319, A2 => Sel(2), A3 => n320, ZN => n316);
   U50 : BUF_X1 port map( A => n315, Z => n176);
   U51 : NOR2_X1 port map( A1 => n165, A2 => n186, ZN => n315);
   U52 : AOI21_X1 port map( B1 => n319, B2 => n320, A => Sel(2), ZN => n186);
   U53 : NAND2_X1 port map( A1 => n200, A2 => n199, ZN => Y(15));
   U54 : AOI22_X1 port map( A1 => A_neg(15), A2 => n151, B1 => A_signal(15), B2
                           => n142, ZN => n200);
   U55 : NAND2_X1 port map( A1 => n198, A2 => n197, ZN => Y(14));
   U56 : AOI222_X1 port map( A1 => A_shifted(14), A2 => n177, B1 => 
                           zeroSignal(14), B2 => n168, C1 => A_neg_shifted(14),
                           C2 => n164, ZN => n197);
   U57 : NAND2_X1 port map( A1 => n202, A2 => n201, ZN => Y(16));
   U58 : AOI222_X1 port map( A1 => A_shifted(16), A2 => n177, B1 => 
                           zeroSignal(16), B2 => n168, C1 => A_neg_shifted(16),
                           C2 => n164, ZN => n201);
   U59 : AOI22_X1 port map( A1 => A_neg(16), A2 => n151, B1 => A_signal(16), B2
                           => n142, ZN => n202);
   U60 : AOI222_X1 port map( A1 => A_shifted(17), A2 => n177, B1 => 
                           zeroSignal(17), B2 => n168, C1 => A_neg_shifted(17),
                           C2 => n164, ZN => n203);
   U61 : AOI222_X1 port map( A1 => A_shifted(18), A2 => n177, B1 => 
                           zeroSignal(18), B2 => n168, C1 => A_neg_shifted(18),
                           C2 => n164, ZN => n205);
   U62 : AOI22_X1 port map( A1 => A_neg(18), A2 => n151, B1 => A_signal(18), B2
                           => n142, ZN => n206);
   U63 : NAND2_X1 port map( A1 => n272, A2 => n271, ZN => Y(48));
   U64 : AOI222_X1 port map( A1 => A_shifted(48), A2 => n180, B1 => 
                           zeroSignal(48), B2 => n171, C1 => A_neg_shifted(48),
                           C2 => n161, ZN => n271);
   U65 : AOI22_X1 port map( A1 => A_neg(48), A2 => n154, B1 => A_signal(48), B2
                           => n145, ZN => n272);
   U66 : NAND2_X1 port map( A1 => n274, A2 => n273, ZN => Y(49));
   U67 : AOI222_X1 port map( A1 => A_shifted(49), A2 => n180, B1 => 
                           zeroSignal(49), B2 => n171, C1 => A_neg_shifted(49),
                           C2 => n161, ZN => n273);
   U68 : AOI22_X1 port map( A1 => A_neg(49), A2 => n154, B1 => A_signal(49), B2
                           => n145, ZN => n274);
   U69 : NAND2_X1 port map( A1 => n278, A2 => n277, ZN => Y(50));
   U70 : AOI222_X1 port map( A1 => A_shifted(50), A2 => n181, B1 => 
                           zeroSignal(50), B2 => n171, C1 => A_neg_shifted(50),
                           C2 => n161, ZN => n277);
   U71 : AOI22_X1 port map( A1 => A_neg(50), A2 => n154, B1 => A_signal(50), B2
                           => n145, ZN => n278);
   U72 : AOI222_X1 port map( A1 => A_shifted(19), A2 => n177, B1 => 
                           zeroSignal(19), B2 => n168, C1 => A_neg_shifted(19),
                           C2 => n164, ZN => n207);
   U73 : NAND2_X1 port map( A1 => n280, A2 => n279, ZN => Y(51));
   U74 : AOI222_X1 port map( A1 => A_shifted(51), A2 => n181, B1 => 
                           zeroSignal(51), B2 => n171, C1 => A_neg_shifted(51),
                           C2 => n161, ZN => n279);
   U75 : AOI22_X1 port map( A1 => A_neg(51), A2 => n154, B1 => A_signal(51), B2
                           => n145, ZN => n280);
   U76 : NAND2_X1 port map( A1 => n282, A2 => n281, ZN => Y(52));
   U77 : AOI22_X1 port map( A1 => A_neg(52), A2 => n154, B1 => A_signal(52), B2
                           => n145, ZN => n282);
   U78 : AOI222_X1 port map( A1 => A_shifted(52), A2 => n181, B1 => 
                           zeroSignal(52), B2 => n171, C1 => A_neg_shifted(52),
                           C2 => n161, ZN => n281);
   U79 : AOI222_X1 port map( A1 => A_shifted(20), A2 => n178, B1 => 
                           zeroSignal(20), B2 => n169, C1 => A_neg_shifted(20),
                           C2 => n164, ZN => n211);
   U80 : NAND2_X1 port map( A1 => n230, A2 => n229, ZN => Y(29));
   U81 : AOI222_X1 port map( A1 => A_shifted(29), A2 => n178, B1 => 
                           zeroSignal(29), B2 => n169, C1 => A_neg_shifted(29),
                           C2 => n163, ZN => n229);
   U82 : AOI22_X1 port map( A1 => A_neg(29), A2 => n152, B1 => A_signal(29), B2
                           => n143, ZN => n230);
   U83 : NAND2_X1 port map( A1 => n226, A2 => n225, ZN => Y(27));
   U84 : AOI222_X1 port map( A1 => A_shifted(27), A2 => n178, B1 => 
                           zeroSignal(27), B2 => n169, C1 => A_neg_shifted(27),
                           C2 => n163, ZN => n225);
   U85 : AOI22_X1 port map( A1 => A_neg(27), A2 => n152, B1 => A_signal(27), B2
                           => n143, ZN => n226);
   U86 : NAND2_X1 port map( A1 => n228, A2 => n227, ZN => Y(28));
   U87 : AOI222_X1 port map( A1 => A_shifted(28), A2 => n178, B1 => 
                           zeroSignal(28), B2 => n169, C1 => A_neg_shifted(28),
                           C2 => n163, ZN => n227);
   U88 : AOI22_X1 port map( A1 => A_neg(28), A2 => n152, B1 => A_signal(28), B2
                           => n143, ZN => n228);
   U89 : NAND2_X1 port map( A1 => n234, A2 => n233, ZN => Y(30));
   U90 : AOI222_X1 port map( A1 => A_shifted(30), A2 => n179, B1 => 
                           zeroSignal(30), B2 => n169, C1 => A_neg_shifted(30),
                           C2 => n163, ZN => n233);
   U91 : AOI22_X1 port map( A1 => A_neg(30), A2 => n152, B1 => A_signal(30), B2
                           => n143, ZN => n234);
   U92 : NAND2_X1 port map( A1 => n236, A2 => n235, ZN => Y(31));
   U93 : AOI222_X1 port map( A1 => A_shifted(31), A2 => n179, B1 => 
                           zeroSignal(31), B2 => n170, C1 => A_neg_shifted(31),
                           C2 => n163, ZN => n235);
   U94 : AOI22_X1 port map( A1 => A_neg(31), A2 => n153, B1 => A_signal(31), B2
                           => n144, ZN => n236);
   U95 : NAND2_X1 port map( A1 => n242, A2 => n241, ZN => Y(34));
   U96 : AOI222_X1 port map( A1 => A_shifted(34), A2 => n179, B1 => 
                           zeroSignal(34), B2 => n170, C1 => A_neg_shifted(34),
                           C2 => n163, ZN => n241);
   U97 : AOI22_X1 port map( A1 => A_neg(34), A2 => n153, B1 => A_signal(34), B2
                           => n144, ZN => n242);
   U98 : NAND2_X1 port map( A1 => n240, A2 => n239, ZN => Y(33));
   U99 : AOI222_X1 port map( A1 => A_shifted(33), A2 => n179, B1 => 
                           zeroSignal(33), B2 => n170, C1 => A_neg_shifted(33),
                           C2 => n163, ZN => n239);
   U100 : AOI22_X1 port map( A1 => A_neg(33), A2 => n153, B1 => A_signal(33), 
                           B2 => n144, ZN => n240);
   U101 : NAND2_X1 port map( A1 => n244, A2 => n243, ZN => Y(35));
   U102 : AOI222_X1 port map( A1 => A_shifted(35), A2 => n179, B1 => 
                           zeroSignal(35), B2 => n170, C1 => A_neg_shifted(35),
                           C2 => n162, ZN => n243);
   U103 : AOI22_X1 port map( A1 => A_neg(35), A2 => n153, B1 => A_signal(35), 
                           B2 => n144, ZN => n244);
   U104 : NAND2_X1 port map( A1 => n246, A2 => n245, ZN => Y(36));
   U105 : AOI222_X1 port map( A1 => A_shifted(36), A2 => n179, B1 => 
                           zeroSignal(36), B2 => n170, C1 => A_neg_shifted(36),
                           C2 => n162, ZN => n245);
   U106 : AOI22_X1 port map( A1 => A_neg(36), A2 => n153, B1 => A_signal(36), 
                           B2 => n144, ZN => n246);
   U107 : NAND2_X1 port map( A1 => n248, A2 => n247, ZN => Y(37));
   U108 : AOI222_X1 port map( A1 => A_shifted(37), A2 => n179, B1 => 
                           zeroSignal(37), B2 => n170, C1 => A_neg_shifted(37),
                           C2 => n162, ZN => n247);
   U109 : AOI22_X1 port map( A1 => A_neg(37), A2 => n153, B1 => A_signal(37), 
                           B2 => n144, ZN => n248);
   U110 : NAND2_X1 port map( A1 => n250, A2 => n249, ZN => Y(38));
   U111 : AOI222_X1 port map( A1 => A_shifted(38), A2 => n179, B1 => 
                           zeroSignal(38), B2 => n170, C1 => A_neg_shifted(38),
                           C2 => n162, ZN => n249);
   U112 : AOI22_X1 port map( A1 => A_neg(38), A2 => n153, B1 => A_signal(38), 
                           B2 => n144, ZN => n250);
   U113 : NAND2_X1 port map( A1 => n252, A2 => n251, ZN => Y(39));
   U114 : AOI222_X1 port map( A1 => A_shifted(39), A2 => n179, B1 => 
                           zeroSignal(39), B2 => n170, C1 => A_neg_shifted(39),
                           C2 => n162, ZN => n251);
   U115 : AOI22_X1 port map( A1 => A_neg(39), A2 => n153, B1 => A_signal(39), 
                           B2 => n144, ZN => n252);
   U116 : NAND2_X1 port map( A1 => n256, A2 => n255, ZN => Y(40));
   U117 : AOI222_X1 port map( A1 => A_shifted(40), A2 => n180, B1 => 
                           zeroSignal(40), B2 => n170, C1 => A_neg_shifted(40),
                           C2 => n162, ZN => n255);
   U118 : AOI22_X1 port map( A1 => A_neg(40), A2 => n153, B1 => A_signal(40), 
                           B2 => n144, ZN => n256);
   U119 : NAND2_X1 port map( A1 => n258, A2 => n257, ZN => Y(41));
   U120 : AOI222_X1 port map( A1 => A_shifted(41), A2 => n180, B1 => 
                           zeroSignal(41), B2 => n170, C1 => A_neg_shifted(41),
                           C2 => n162, ZN => n257);
   U121 : AOI22_X1 port map( A1 => A_neg(41), A2 => n153, B1 => A_signal(41), 
                           B2 => n144, ZN => n258);
   U122 : AOI22_X1 port map( A1 => A_neg(21), A2 => n152, B1 => A_signal(21), 
                           B2 => n143, ZN => n214);
   U123 : AOI222_X1 port map( A1 => A_shifted(21), A2 => n178, B1 => 
                           zeroSignal(21), B2 => n169, C1 => A_neg_shifted(21),
                           C2 => n164, ZN => n213);
   U124 : NAND2_X1 port map( A1 => n238, A2 => n237, ZN => Y(32));
   U125 : AOI22_X1 port map( A1 => A_neg(32), A2 => n153, B1 => A_signal(32), 
                           B2 => n144, ZN => n238);
   U126 : AOI222_X1 port map( A1 => A_shifted(32), A2 => n179, B1 => 
                           zeroSignal(32), B2 => n170, C1 => A_neg_shifted(32),
                           C2 => n163, ZN => n237);
   U127 : NAND2_X1 port map( A1 => n264, A2 => n263, ZN => Y(44));
   U128 : AOI222_X1 port map( A1 => A_shifted(44), A2 => n180, B1 => 
                           zeroSignal(44), B2 => n171, C1 => A_neg_shifted(44),
                           C2 => n162, ZN => n263);
   U129 : AOI22_X1 port map( A1 => A_neg(44), A2 => n154, B1 => A_signal(44), 
                           B2 => n145, ZN => n264);
   U130 : NAND2_X1 port map( A1 => n260, A2 => n259, ZN => Y(42));
   U131 : AOI222_X1 port map( A1 => A_shifted(42), A2 => n180, B1 => 
                           zeroSignal(42), B2 => n171, C1 => A_neg_shifted(42),
                           C2 => n162, ZN => n259);
   U132 : AOI22_X1 port map( A1 => A_neg(42), A2 => n154, B1 => A_signal(42), 
                           B2 => n145, ZN => n260);
   U133 : NAND2_X1 port map( A1 => n266, A2 => n265, ZN => Y(45));
   U134 : AOI222_X1 port map( A1 => A_shifted(45), A2 => n180, B1 => 
                           zeroSignal(45), B2 => n171, C1 => A_neg_shifted(45),
                           C2 => n162, ZN => n265);
   U135 : AOI22_X1 port map( A1 => A_neg(45), A2 => n154, B1 => A_signal(45), 
                           B2 => n145, ZN => n266);
   U136 : NAND2_X1 port map( A1 => n268, A2 => n267, ZN => Y(46));
   U137 : AOI222_X1 port map( A1 => A_shifted(46), A2 => n180, B1 => 
                           zeroSignal(46), B2 => n171, C1 => A_neg_shifted(46),
                           C2 => n161, ZN => n267);
   U138 : AOI22_X1 port map( A1 => A_neg(46), A2 => n154, B1 => A_signal(46), 
                           B2 => n145, ZN => n268);
   U139 : NAND2_X1 port map( A1 => n220, A2 => n219, ZN => Y(24));
   U140 : AOI222_X1 port map( A1 => A_shifted(24), A2 => n178, B1 => 
                           zeroSignal(24), B2 => n169, C1 => A_neg_shifted(24),
                           C2 => n163, ZN => n219);
   U141 : AOI22_X1 port map( A1 => A_neg(24), A2 => n152, B1 => A_signal(24), 
                           B2 => n143, ZN => n220);
   U142 : NAND2_X1 port map( A1 => n224, A2 => n223, ZN => Y(26));
   U143 : AOI222_X1 port map( A1 => A_shifted(26), A2 => n178, B1 => 
                           zeroSignal(26), B2 => n169, C1 => A_neg_shifted(26),
                           C2 => n163, ZN => n223);
   U144 : AOI22_X1 port map( A1 => A_neg(26), A2 => n152, B1 => A_signal(26), 
                           B2 => n143, ZN => n224);
   U145 : NAND2_X1 port map( A1 => n262, A2 => n261, ZN => Y(43));
   U146 : AOI22_X1 port map( A1 => A_neg(43), A2 => n154, B1 => A_signal(43), 
                           B2 => n145, ZN => n262);
   U147 : AOI222_X1 port map( A1 => A_shifted(43), A2 => n180, B1 => 
                           zeroSignal(43), B2 => n171, C1 => A_neg_shifted(43),
                           C2 => n162, ZN => n261);
   U148 : NAND2_X1 port map( A1 => n286, A2 => n285, ZN => Y(54));
   U149 : AOI222_X1 port map( A1 => A_shifted(54), A2 => n181, B1 => 
                           zeroSignal(54), B2 => n172, C1 => A_neg_shifted(54),
                           C2 => n161, ZN => n285);
   U150 : AOI22_X1 port map( A1 => A_neg(54), A2 => n155, B1 => A_signal(54), 
                           B2 => n146, ZN => n286);
   U151 : NAND2_X1 port map( A1 => n284, A2 => n283, ZN => Y(53));
   U152 : AOI22_X1 port map( A1 => A_neg(53), A2 => n155, B1 => A_signal(53), 
                           B2 => n146, ZN => n284);
   U153 : AOI222_X1 port map( A1 => A_shifted(53), A2 => n181, B1 => 
                           zeroSignal(53), B2 => n172, C1 => A_neg_shifted(53),
                           C2 => n161, ZN => n283);
   U154 : NAND2_X1 port map( A1 => n216, A2 => n215, ZN => Y(22));
   U155 : AOI22_X1 port map( A1 => A_neg(22), A2 => n152, B1 => A_signal(22), 
                           B2 => n143, ZN => n216);
   U156 : AOI222_X1 port map( A1 => A_shifted(22), A2 => n178, B1 => 
                           zeroSignal(22), B2 => n169, C1 => A_neg_shifted(22),
                           C2 => n164, ZN => n215);
   U157 : NAND2_X1 port map( A1 => n270, A2 => n269, ZN => Y(47));
   U158 : AOI222_X1 port map( A1 => A_shifted(47), A2 => n180, B1 => 
                           zeroSignal(47), B2 => n171, C1 => A_neg_shifted(47),
                           C2 => n161, ZN => n269);
   U159 : AOI22_X1 port map( A1 => A_neg(47), A2 => n154, B1 => A_signal(47), 
                           B2 => n145, ZN => n270);
   U160 : NAND2_X1 port map( A1 => n222, A2 => n221, ZN => Y(25));
   U161 : AOI22_X1 port map( A1 => A_neg(25), A2 => n152, B1 => A_signal(25), 
                           B2 => n143, ZN => n222);
   U162 : AOI222_X1 port map( A1 => A_shifted(25), A2 => n178, B1 => 
                           zeroSignal(25), B2 => n169, C1 => A_neg_shifted(25),
                           C2 => n163, ZN => n221);
   U163 : NAND2_X1 port map( A1 => n288, A2 => n287, ZN => Y(55));
   U164 : AOI22_X1 port map( A1 => A_neg(55), A2 => n155, B1 => A_signal(55), 
                           B2 => n146, ZN => n288);
   U165 : AOI222_X1 port map( A1 => A_shifted(55), A2 => n181, B1 => 
                           zeroSignal(55), B2 => n172, C1 => A_neg_shifted(55),
                           C2 => n161, ZN => n287);
   U166 : NAND2_X1 port map( A1 => n218, A2 => n217, ZN => Y(23));
   U167 : AOI22_X1 port map( A1 => A_neg(23), A2 => n152, B1 => A_signal(23), 
                           B2 => n143, ZN => n218);
   U168 : AOI222_X1 port map( A1 => A_shifted(23), A2 => n178, B1 => 
                           zeroSignal(23), B2 => n169, C1 => A_neg_shifted(23),
                           C2 => n164, ZN => n217);
   U169 : NAND2_X1 port map( A1 => n292, A2 => n291, ZN => Y(57));
   U170 : AOI22_X1 port map( A1 => A_neg(57), A2 => n155, B1 => A_signal(57), 
                           B2 => n146, ZN => n292);
   U171 : NAND2_X1 port map( A1 => n296, A2 => n295, ZN => Y(59));
   U172 : AOI222_X1 port map( A1 => A_shifted(59), A2 => n181, B1 => 
                           zeroSignal(59), B2 => n172, C1 => A_neg_shifted(59),
                           C2 => n160, ZN => n295);
   U173 : NAND2_X1 port map( A1 => n294, A2 => n293, ZN => Y(58));
   U174 : AOI222_X1 port map( A1 => A_shifted(58), A2 => n181, B1 => 
                           zeroSignal(58), B2 => n172, C1 => A_neg_shifted(58),
                           C2 => n160, ZN => n293);
   U175 : AOI22_X1 port map( A1 => A_neg(58), A2 => n155, B1 => A_signal(58), 
                           B2 => n146, ZN => n294);
   U176 : NAND2_X1 port map( A1 => n290, A2 => n289, ZN => Y(56));
   U177 : AOI222_X1 port map( A1 => A_shifted(56), A2 => n181, B1 => 
                           zeroSignal(56), B2 => n172, C1 => A_neg_shifted(56),
                           C2 => n161, ZN => n289);
   U178 : NAND2_X1 port map( A1 => n306, A2 => n305, ZN => Y(63));
   U179 : AOI222_X1 port map( A1 => A_shifted(63), A2 => n182, B1 => 
                           zeroSignal(63), B2 => n172, C1 => A_neg_shifted(63),
                           C2 => n160, ZN => n305);
   U180 : AOI22_X1 port map( A1 => A_neg(63), A2 => n155, B1 => A_signal(63), 
                           B2 => n146, ZN => n306);
   U181 : NAND2_X1 port map( A1 => n300, A2 => n299, ZN => Y(60));
   U182 : AOI22_X1 port map( A1 => A_neg(60), A2 => n155, B1 => A_signal(60), 
                           B2 => n146, ZN => n300);
   U183 : NAND2_X1 port map( A1 => n302, A2 => n301, ZN => Y(61));
   U184 : AOI222_X1 port map( A1 => A_shifted(61), A2 => n182, B1 => 
                           zeroSignal(61), B2 => n172, C1 => A_neg_shifted(61),
                           C2 => n160, ZN => n301);
   U185 : AOI22_X1 port map( A1 => A_neg(61), A2 => n155, B1 => A_signal(61), 
                           B2 => n146, ZN => n302);
   U186 : NAND2_X1 port map( A1 => n304, A2 => n303, ZN => Y(62));
   U187 : AOI222_X1 port map( A1 => A_shifted(62), A2 => n182, B1 => 
                           zeroSignal(62), B2 => n172, C1 => A_neg_shifted(62),
                           C2 => n160, ZN => n303);
   U188 : AOI22_X1 port map( A1 => A_neg(62), A2 => n155, B1 => A_signal(62), 
                           B2 => n146, ZN => n304);
   U189 : NAND2_X1 port map( A1 => n188, A2 => n187, ZN => Y(0));
   U190 : AOI22_X1 port map( A1 => A_neg(0), A2 => n151, B1 => A_signal(0), B2 
                           => n142, ZN => n188);
   U191 : AOI222_X1 port map( A1 => A_shifted(0), A2 => n177, B1 => 
                           zeroSignal(0), B2 => n168, C1 => A_neg_shifted(0), 
                           C2 => n165, ZN => n187);
   U192 : NAND2_X1 port map( A1 => n210, A2 => n209, ZN => Y(1));
   U193 : AOI22_X1 port map( A1 => A_neg(1), A2 => n151, B1 => A_signal(1), B2 
                           => n142, ZN => n210);
   U194 : AOI222_X1 port map( A1 => A_shifted(1), A2 => n178, B1 => 
                           zeroSignal(1), B2 => n168, C1 => A_neg_shifted(1), 
                           C2 => n164, ZN => n209);
   U195 : NAND2_X1 port map( A1 => n232, A2 => n231, ZN => Y(2));
   U196 : AOI22_X1 port map( A1 => A_neg(2), A2 => n152, B1 => A_signal(2), B2 
                           => n143, ZN => n232);
   U197 : AOI222_X1 port map( A1 => A_shifted(2), A2 => n179, B1 => 
                           zeroSignal(2), B2 => n169, C1 => A_neg_shifted(2), 
                           C2 => n163, ZN => n231);
   U198 : NAND2_X1 port map( A1 => n254, A2 => n253, ZN => Y(3));
   U199 : AOI22_X1 port map( A1 => A_neg(3), A2 => n153, B1 => A_signal(3), B2 
                           => n144, ZN => n254);
   U200 : AOI222_X1 port map( A1 => A_shifted(3), A2 => n180, B1 => 
                           zeroSignal(3), B2 => n170, C1 => A_neg_shifted(3), 
                           C2 => n162, ZN => n253);
   U201 : NAND2_X1 port map( A1 => n276, A2 => n275, ZN => Y(4));
   U202 : AOI22_X1 port map( A1 => A_neg(4), A2 => n154, B1 => A_signal(4), B2 
                           => n145, ZN => n276);
   U203 : AOI222_X1 port map( A1 => A_shifted(4), A2 => n181, B1 => 
                           zeroSignal(4), B2 => n171, C1 => A_neg_shifted(4), 
                           C2 => n161, ZN => n275);
   U204 : NAND2_X1 port map( A1 => n298, A2 => n297, ZN => Y(5));
   U205 : AOI22_X1 port map( A1 => A_neg(5), A2 => n155, B1 => A_signal(5), B2 
                           => n146, ZN => n298);
   U206 : AOI222_X1 port map( A1 => A_shifted(5), A2 => n182, B1 => 
                           zeroSignal(5), B2 => n172, C1 => A_neg_shifted(5), 
                           C2 => n160, ZN => n297);
   U207 : NAND2_X1 port map( A1 => n308, A2 => n307, ZN => Y(6));
   U208 : AOI22_X1 port map( A1 => A_neg(6), A2 => n156, B1 => A_signal(6), B2 
                           => n147, ZN => n308);
   U209 : AOI222_X1 port map( A1 => A_shifted(6), A2 => n182, B1 => 
                           zeroSignal(6), B2 => n173, C1 => A_neg_shifted(6), 
                           C2 => n160, ZN => n307);
   U210 : NAND2_X1 port map( A1 => n310, A2 => n309, ZN => Y(7));
   U211 : AOI22_X1 port map( A1 => A_neg(7), A2 => n156, B1 => A_signal(7), B2 
                           => n147, ZN => n310);
   U212 : AOI222_X1 port map( A1 => A_shifted(7), A2 => n182, B1 => 
                           zeroSignal(7), B2 => n173, C1 => A_neg_shifted(7), 
                           C2 => n160, ZN => n309);
   U213 : NAND2_X1 port map( A1 => n312, A2 => n311, ZN => Y(8));
   U214 : AOI22_X1 port map( A1 => A_neg(8), A2 => n156, B1 => A_signal(8), B2 
                           => n147, ZN => n312);
   U215 : AOI222_X1 port map( A1 => A_shifted(8), A2 => n182, B1 => 
                           zeroSignal(8), B2 => n173, C1 => A_neg_shifted(8), 
                           C2 => n160, ZN => n311);
   U216 : NAND2_X1 port map( A1 => n318, A2 => n317, ZN => Y(9));
   U217 : AOI22_X1 port map( A1 => A_neg(9), A2 => n156, B1 => A_signal(9), B2 
                           => n147, ZN => n318);
   U218 : AOI222_X1 port map( A1 => A_shifted(9), A2 => n182, B1 => 
                           zeroSignal(9), B2 => n173, C1 => A_neg_shifted(9), 
                           C2 => n160, ZN => n317);
   U219 : NAND2_X1 port map( A1 => n190, A2 => n189, ZN => Y(10));
   U220 : AOI22_X1 port map( A1 => A_neg(10), A2 => n151, B1 => A_signal(10), 
                           B2 => n142, ZN => n190);
   U221 : AOI222_X1 port map( A1 => A_shifted(10), A2 => n177, B1 => 
                           zeroSignal(10), B2 => n168, C1 => A_neg_shifted(10),
                           C2 => n165, ZN => n189);
   U222 : NAND2_X1 port map( A1 => n192, A2 => n191, ZN => Y(11));
   U223 : AOI22_X1 port map( A1 => A_neg(11), A2 => n151, B1 => A_signal(11), 
                           B2 => n142, ZN => n192);
   U224 : AOI222_X1 port map( A1 => A_shifted(11), A2 => n177, B1 => 
                           zeroSignal(11), B2 => n168, C1 => A_neg_shifted(11),
                           C2 => n165, ZN => n191);
   U225 : NAND2_X1 port map( A1 => n194, A2 => n193, ZN => Y(12));
   U226 : AOI22_X1 port map( A1 => A_neg(12), A2 => n151, B1 => A_signal(12), 
                           B2 => n142, ZN => n194);
   U227 : AOI222_X1 port map( A1 => A_shifted(12), A2 => n177, B1 => 
                           zeroSignal(12), B2 => n168, C1 => A_neg_shifted(12),
                           C2 => n165, ZN => n193);
   U228 : NAND2_X1 port map( A1 => n196, A2 => n195, ZN => Y(13));
   U229 : AOI22_X1 port map( A1 => A_neg(13), A2 => n151, B1 => A_signal(13), 
                           B2 => n142, ZN => n196);
   U230 : AOI222_X1 port map( A1 => A_shifted(13), A2 => n177, B1 => 
                           zeroSignal(13), B2 => n168, C1 => A_neg_shifted(13),
                           C2 => n164, ZN => n195);
   U231 : AOI222_X1 port map( A1 => A_shifted(15), A2 => n177, B1 => 
                           zeroSignal(15), B2 => n168, C1 => A_neg_shifted(15),
                           C2 => n164, ZN => n199);
   U232 : AOI22_X1 port map( A1 => A_neg(14), A2 => n151, B1 => A_signal(14), 
                           B2 => n142, ZN => n198);
   U233 : AOI22_X1 port map( A1 => A_neg(20), A2 => n152, B1 => A_signal(20), 
                           B2 => n143, ZN => n212);
   U234 : NAND2_X1 port map( A1 => n214, A2 => n213, ZN => Y(21));
   U235 : AOI22_X1 port map( A1 => A_neg(19), A2 => n151, B1 => A_signal(19), 
                           B2 => n142, ZN => n208);
   U236 : NAND2_X1 port map( A1 => n212, A2 => n211, ZN => Y(20));
   U237 : NAND2_X1 port map( A1 => n208, A2 => n207, ZN => Y(19));
   U238 : AOI22_X1 port map( A1 => A_neg(17), A2 => n151, B1 => A_signal(17), 
                           B2 => n142, ZN => n204);
   U239 : NAND2_X1 port map( A1 => n206, A2 => n205, ZN => Y(18));
   U240 : NAND2_X1 port map( A1 => n204, A2 => n203, ZN => Y(17));
   U241 : AOI222_X1 port map( A1 => A_shifted(60), A2 => n182, B1 => 
                           zeroSignal(60), B2 => n172, C1 => A_neg_shifted(60),
                           C2 => n160, ZN => n299);
   U242 : AOI22_X1 port map( A1 => A_neg(59), A2 => n155, B1 => A_signal(59), 
                           B2 => n146, ZN => n296);
   U243 : AOI222_X1 port map( A1 => A_shifted(57), A2 => n181, B1 => 
                           zeroSignal(57), B2 => n172, C1 => A_neg_shifted(57),
                           C2 => n160, ZN => n291);
   U244 : AOI22_X1 port map( A1 => A_neg(56), A2 => n155, B1 => A_signal(56), 
                           B2 => n146, ZN => n290);

end SYN_BEHAVIORAL_2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity MUX51_MuxNbit64_8 is

   port( zeroSignal, A_signal, A_neg, A_shifted, A_neg_shifted : in 
         std_logic_vector (63 downto 0);  Sel : in std_logic_vector (2 downto 
         0);  Y : out std_logic_vector (63 downto 0));

end MUX51_MuxNbit64_8;

architecture SYN_BEHAVIORAL_2 of MUX51_MuxNbit64_8 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, 
      n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, 
      n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, 
      n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, 
      n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, 
      n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, 
      n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, 
      n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, 
      n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, 
      n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, 
      n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, 
      n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, 
      n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, 
      n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, 
      n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, 
      n320 : std_logic;

begin
   
   U1 : AND3_X1 port map( A1 => n319, A2 => n320, A3 => Sel(2), ZN => n141);
   U2 : BUF_X1 port map( A => n141, Z => n166);
   U3 : BUF_X1 port map( A => n159, Z => n158);
   U4 : BUF_X1 port map( A => n185, Z => n184);
   U5 : BUF_X1 port map( A => n150, Z => n149);
   U6 : BUF_X1 port map( A => n141, Z => n167);
   U7 : BUF_X1 port map( A => n185, Z => n183);
   U8 : BUF_X1 port map( A => n159, Z => n157);
   U9 : BUF_X1 port map( A => n150, Z => n148);
   U10 : BUF_X1 port map( A => n176, Z => n175);
   U11 : BUF_X1 port map( A => n176, Z => n174);
   U12 : BUF_X1 port map( A => n184, Z => n177);
   U13 : BUF_X1 port map( A => n158, Z => n151);
   U14 : BUF_X1 port map( A => n149, Z => n142);
   U15 : BUF_X1 port map( A => n166, Z => n164);
   U16 : BUF_X1 port map( A => n184, Z => n178);
   U17 : BUF_X1 port map( A => n158, Z => n152);
   U18 : BUF_X1 port map( A => n149, Z => n143);
   U19 : BUF_X1 port map( A => n166, Z => n163);
   U20 : BUF_X1 port map( A => n184, Z => n179);
   U21 : BUF_X1 port map( A => n158, Z => n153);
   U22 : BUF_X1 port map( A => n149, Z => n144);
   U23 : BUF_X1 port map( A => n167, Z => n162);
   U24 : BUF_X1 port map( A => n183, Z => n180);
   U25 : BUF_X1 port map( A => n157, Z => n154);
   U26 : BUF_X1 port map( A => n148, Z => n145);
   U27 : BUF_X1 port map( A => n167, Z => n161);
   U28 : BUF_X1 port map( A => n183, Z => n181);
   U29 : BUF_X1 port map( A => n157, Z => n155);
   U30 : BUF_X1 port map( A => n148, Z => n146);
   U31 : BUF_X1 port map( A => n167, Z => n160);
   U32 : BUF_X1 port map( A => n183, Z => n182);
   U33 : BUF_X1 port map( A => n175, Z => n168);
   U34 : BUF_X1 port map( A => n175, Z => n169);
   U35 : BUF_X1 port map( A => n175, Z => n170);
   U36 : BUF_X1 port map( A => n174, Z => n171);
   U37 : BUF_X1 port map( A => n174, Z => n172);
   U38 : BUF_X1 port map( A => n166, Z => n165);
   U39 : BUF_X1 port map( A => n157, Z => n156);
   U40 : BUF_X1 port map( A => n148, Z => n147);
   U41 : BUF_X1 port map( A => n174, Z => n173);
   U42 : BUF_X1 port map( A => n316, Z => n185);
   U43 : NOR3_X1 port map( A1 => n319, A2 => Sel(2), A3 => n320, ZN => n316);
   U44 : INV_X1 port map( A => Sel(1), ZN => n320);
   U45 : BUF_X1 port map( A => n314, Z => n159);
   U46 : NOR3_X1 port map( A1 => Sel(0), A2 => Sel(2), A3 => n320, ZN => n314);
   U47 : INV_X1 port map( A => Sel(0), ZN => n319);
   U48 : BUF_X1 port map( A => n313, Z => n150);
   U49 : NOR3_X1 port map( A1 => Sel(1), A2 => Sel(2), A3 => n319, ZN => n313);
   U50 : BUF_X1 port map( A => n315, Z => n176);
   U51 : NOR2_X1 port map( A1 => n165, A2 => n186, ZN => n315);
   U52 : AOI21_X1 port map( B1 => n319, B2 => n320, A => Sel(2), ZN => n186);
   U53 : NAND2_X1 port map( A1 => n260, A2 => n259, ZN => Y(42));
   U54 : AOI222_X1 port map( A1 => A_shifted(42), A2 => n180, B1 => 
                           zeroSignal(42), B2 => n171, C1 => A_neg_shifted(42),
                           C2 => n162, ZN => n259);
   U55 : AOI22_X1 port map( A1 => A_neg(42), A2 => n154, B1 => A_signal(42), B2
                           => n145, ZN => n260);
   U56 : NAND2_X1 port map( A1 => n204, A2 => n203, ZN => Y(17));
   U57 : AOI22_X1 port map( A1 => A_neg(17), A2 => n151, B1 => A_signal(17), B2
                           => n142, ZN => n204);
   U58 : AOI222_X1 port map( A1 => A_shifted(17), A2 => n177, B1 => 
                           zeroSignal(17), B2 => n168, C1 => A_neg_shifted(17),
                           C2 => n164, ZN => n203);
   U59 : NAND2_X1 port map( A1 => n202, A2 => n201, ZN => Y(16));
   U60 : AOI222_X1 port map( A1 => A_shifted(16), A2 => n177, B1 => 
                           zeroSignal(16), B2 => n168, C1 => A_neg_shifted(16),
                           C2 => n164, ZN => n201);
   U61 : AOI22_X1 port map( A1 => A_neg(16), A2 => n151, B1 => A_signal(16), B2
                           => n142, ZN => n202);
   U62 : NAND2_X1 port map( A1 => n236, A2 => n235, ZN => Y(31));
   U63 : AOI222_X1 port map( A1 => A_shifted(31), A2 => n179, B1 => 
                           zeroSignal(31), B2 => n170, C1 => A_neg_shifted(31),
                           C2 => n163, ZN => n235);
   U64 : AOI22_X1 port map( A1 => A_neg(31), A2 => n153, B1 => A_signal(31), B2
                           => n144, ZN => n236);
   U65 : NAND2_X1 port map( A1 => n230, A2 => n229, ZN => Y(29));
   U66 : AOI222_X1 port map( A1 => A_shifted(29), A2 => n178, B1 => 
                           zeroSignal(29), B2 => n169, C1 => A_neg_shifted(29),
                           C2 => n163, ZN => n229);
   U67 : AOI22_X1 port map( A1 => A_neg(29), A2 => n152, B1 => A_signal(29), B2
                           => n143, ZN => n230);
   U68 : NAND2_X1 port map( A1 => n234, A2 => n233, ZN => Y(30));
   U69 : AOI222_X1 port map( A1 => A_shifted(30), A2 => n179, B1 => 
                           zeroSignal(30), B2 => n169, C1 => A_neg_shifted(30),
                           C2 => n163, ZN => n233);
   U70 : AOI22_X1 port map( A1 => A_neg(30), A2 => n152, B1 => A_signal(30), B2
                           => n143, ZN => n234);
   U71 : NAND2_X1 port map( A1 => n206, A2 => n205, ZN => Y(18));
   U72 : AOI22_X1 port map( A1 => A_neg(18), A2 => n151, B1 => A_signal(18), B2
                           => n142, ZN => n206);
   U73 : AOI222_X1 port map( A1 => A_shifted(18), A2 => n177, B1 => 
                           zeroSignal(18), B2 => n168, C1 => A_neg_shifted(18),
                           C2 => n164, ZN => n205);
   U74 : NAND2_X1 port map( A1 => n238, A2 => n237, ZN => Y(32));
   U75 : AOI222_X1 port map( A1 => A_shifted(32), A2 => n179, B1 => 
                           zeroSignal(32), B2 => n170, C1 => A_neg_shifted(32),
                           C2 => n163, ZN => n237);
   U76 : AOI22_X1 port map( A1 => A_neg(32), A2 => n153, B1 => A_signal(32), B2
                           => n144, ZN => n238);
   U77 : NAND2_X1 port map( A1 => n240, A2 => n239, ZN => Y(33));
   U78 : AOI222_X1 port map( A1 => A_shifted(33), A2 => n179, B1 => 
                           zeroSignal(33), B2 => n170, C1 => A_neg_shifted(33),
                           C2 => n163, ZN => n239);
   U79 : AOI22_X1 port map( A1 => A_neg(33), A2 => n153, B1 => A_signal(33), B2
                           => n144, ZN => n240);
   U80 : NAND2_X1 port map( A1 => n244, A2 => n243, ZN => Y(35));
   U81 : AOI222_X1 port map( A1 => A_shifted(35), A2 => n179, B1 => 
                           zeroSignal(35), B2 => n170, C1 => A_neg_shifted(35),
                           C2 => n162, ZN => n243);
   U82 : AOI22_X1 port map( A1 => A_neg(35), A2 => n153, B1 => A_signal(35), B2
                           => n144, ZN => n244);
   U83 : NAND2_X1 port map( A1 => n246, A2 => n245, ZN => Y(36));
   U84 : AOI222_X1 port map( A1 => A_shifted(36), A2 => n179, B1 => 
                           zeroSignal(36), B2 => n170, C1 => A_neg_shifted(36),
                           C2 => n162, ZN => n245);
   U85 : AOI22_X1 port map( A1 => A_neg(36), A2 => n153, B1 => A_signal(36), B2
                           => n144, ZN => n246);
   U86 : NAND2_X1 port map( A1 => n248, A2 => n247, ZN => Y(37));
   U87 : AOI222_X1 port map( A1 => A_shifted(37), A2 => n179, B1 => 
                           zeroSignal(37), B2 => n170, C1 => A_neg_shifted(37),
                           C2 => n162, ZN => n247);
   U88 : AOI22_X1 port map( A1 => A_neg(37), A2 => n153, B1 => A_signal(37), B2
                           => n144, ZN => n248);
   U89 : NAND2_X1 port map( A1 => n250, A2 => n249, ZN => Y(38));
   U90 : AOI222_X1 port map( A1 => A_shifted(38), A2 => n179, B1 => 
                           zeroSignal(38), B2 => n170, C1 => A_neg_shifted(38),
                           C2 => n162, ZN => n249);
   U91 : AOI22_X1 port map( A1 => A_neg(38), A2 => n153, B1 => A_signal(38), B2
                           => n144, ZN => n250);
   U92 : NAND2_X1 port map( A1 => n252, A2 => n251, ZN => Y(39));
   U93 : AOI222_X1 port map( A1 => A_shifted(39), A2 => n179, B1 => 
                           zeroSignal(39), B2 => n170, C1 => A_neg_shifted(39),
                           C2 => n162, ZN => n251);
   U94 : AOI22_X1 port map( A1 => A_neg(39), A2 => n153, B1 => A_signal(39), B2
                           => n144, ZN => n252);
   U95 : NAND2_X1 port map( A1 => n256, A2 => n255, ZN => Y(40));
   U96 : AOI222_X1 port map( A1 => A_shifted(40), A2 => n180, B1 => 
                           zeroSignal(40), B2 => n170, C1 => A_neg_shifted(40),
                           C2 => n162, ZN => n255);
   U97 : AOI22_X1 port map( A1 => A_neg(40), A2 => n153, B1 => A_signal(40), B2
                           => n144, ZN => n256);
   U98 : NAND2_X1 port map( A1 => n258, A2 => n257, ZN => Y(41));
   U99 : AOI222_X1 port map( A1 => A_shifted(41), A2 => n180, B1 => 
                           zeroSignal(41), B2 => n170, C1 => A_neg_shifted(41),
                           C2 => n162, ZN => n257);
   U100 : AOI22_X1 port map( A1 => A_neg(41), A2 => n153, B1 => A_signal(41), 
                           B2 => n144, ZN => n258);
   U101 : NAND2_X1 port map( A1 => n262, A2 => n261, ZN => Y(43));
   U102 : AOI222_X1 port map( A1 => A_shifted(43), A2 => n180, B1 => 
                           zeroSignal(43), B2 => n171, C1 => A_neg_shifted(43),
                           C2 => n162, ZN => n261);
   U103 : AOI22_X1 port map( A1 => A_neg(43), A2 => n154, B1 => A_signal(43), 
                           B2 => n145, ZN => n262);
   U104 : NAND2_X1 port map( A1 => n264, A2 => n263, ZN => Y(44));
   U105 : AOI222_X1 port map( A1 => A_shifted(44), A2 => n180, B1 => 
                           zeroSignal(44), B2 => n171, C1 => A_neg_shifted(44),
                           C2 => n162, ZN => n263);
   U106 : AOI22_X1 port map( A1 => A_neg(44), A2 => n154, B1 => A_signal(44), 
                           B2 => n145, ZN => n264);
   U107 : NAND2_X1 port map( A1 => n268, A2 => n267, ZN => Y(46));
   U108 : AOI222_X1 port map( A1 => A_shifted(46), A2 => n180, B1 => 
                           zeroSignal(46), B2 => n171, C1 => A_neg_shifted(46),
                           C2 => n161, ZN => n267);
   U109 : AOI22_X1 port map( A1 => A_neg(46), A2 => n154, B1 => A_signal(46), 
                           B2 => n145, ZN => n268);
   U110 : NAND2_X1 port map( A1 => n242, A2 => n241, ZN => Y(34));
   U111 : AOI22_X1 port map( A1 => A_neg(34), A2 => n153, B1 => A_signal(34), 
                           B2 => n144, ZN => n242);
   U112 : AOI222_X1 port map( A1 => A_shifted(34), A2 => n179, B1 => 
                           zeroSignal(34), B2 => n170, C1 => A_neg_shifted(34),
                           C2 => n163, ZN => n241);
   U113 : NAND2_X1 port map( A1 => n270, A2 => n269, ZN => Y(47));
   U114 : AOI222_X1 port map( A1 => A_shifted(47), A2 => n180, B1 => 
                           zeroSignal(47), B2 => n171, C1 => A_neg_shifted(47),
                           C2 => n161, ZN => n269);
   U115 : AOI22_X1 port map( A1 => A_neg(47), A2 => n154, B1 => A_signal(47), 
                           B2 => n145, ZN => n270);
   U116 : NAND2_X1 port map( A1 => n208, A2 => n207, ZN => Y(19));
   U117 : AOI222_X1 port map( A1 => A_shifted(19), A2 => n177, B1 => 
                           zeroSignal(19), B2 => n168, C1 => A_neg_shifted(19),
                           C2 => n164, ZN => n207);
   U118 : NAND2_X1 port map( A1 => n272, A2 => n271, ZN => Y(48));
   U119 : AOI222_X1 port map( A1 => A_shifted(48), A2 => n180, B1 => 
                           zeroSignal(48), B2 => n171, C1 => A_neg_shifted(48),
                           C2 => n161, ZN => n271);
   U120 : AOI22_X1 port map( A1 => A_neg(48), A2 => n154, B1 => A_signal(48), 
                           B2 => n145, ZN => n272);
   U121 : NAND2_X1 port map( A1 => n266, A2 => n265, ZN => Y(45));
   U122 : AOI22_X1 port map( A1 => A_neg(45), A2 => n154, B1 => A_signal(45), 
                           B2 => n145, ZN => n266);
   U123 : AOI222_X1 port map( A1 => A_shifted(45), A2 => n180, B1 => 
                           zeroSignal(45), B2 => n171, C1 => A_neg_shifted(45),
                           C2 => n162, ZN => n265);
   U124 : NAND2_X1 port map( A1 => n274, A2 => n273, ZN => Y(49));
   U125 : AOI222_X1 port map( A1 => A_shifted(49), A2 => n180, B1 => 
                           zeroSignal(49), B2 => n171, C1 => A_neg_shifted(49),
                           C2 => n161, ZN => n273);
   U126 : AOI22_X1 port map( A1 => A_neg(49), A2 => n154, B1 => A_signal(49), 
                           B2 => n145, ZN => n274);
   U127 : NAND2_X1 port map( A1 => n224, A2 => n223, ZN => Y(26));
   U128 : AOI222_X1 port map( A1 => A_shifted(26), A2 => n178, B1 => 
                           zeroSignal(26), B2 => n169, C1 => A_neg_shifted(26),
                           C2 => n163, ZN => n223);
   U129 : AOI22_X1 port map( A1 => A_neg(26), A2 => n152, B1 => A_signal(26), 
                           B2 => n143, ZN => n224);
   U130 : NAND2_X1 port map( A1 => n228, A2 => n227, ZN => Y(28));
   U131 : AOI222_X1 port map( A1 => A_shifted(28), A2 => n178, B1 => 
                           zeroSignal(28), B2 => n169, C1 => A_neg_shifted(28),
                           C2 => n163, ZN => n227);
   U132 : AOI22_X1 port map( A1 => A_neg(28), A2 => n152, B1 => A_signal(28), 
                           B2 => n143, ZN => n228);
   U133 : NAND2_X1 port map( A1 => n212, A2 => n211, ZN => Y(20));
   U134 : AOI22_X1 port map( A1 => A_neg(20), A2 => n152, B1 => A_signal(20), 
                           B2 => n143, ZN => n212);
   U135 : AOI222_X1 port map( A1 => A_shifted(20), A2 => n178, B1 => 
                           zeroSignal(20), B2 => n169, C1 => A_neg_shifted(20),
                           C2 => n164, ZN => n211);
   U136 : NAND2_X1 port map( A1 => n278, A2 => n277, ZN => Y(50));
   U137 : AOI222_X1 port map( A1 => A_shifted(50), A2 => n181, B1 => 
                           zeroSignal(50), B2 => n171, C1 => A_neg_shifted(50),
                           C2 => n161, ZN => n277);
   U138 : AOI22_X1 port map( A1 => A_neg(50), A2 => n154, B1 => A_signal(50), 
                           B2 => n145, ZN => n278);
   U139 : NAND2_X1 port map( A1 => n226, A2 => n225, ZN => Y(27));
   U140 : AOI22_X1 port map( A1 => A_neg(27), A2 => n152, B1 => A_signal(27), 
                           B2 => n143, ZN => n226);
   U141 : AOI222_X1 port map( A1 => A_shifted(27), A2 => n178, B1 => 
                           zeroSignal(27), B2 => n169, C1 => A_neg_shifted(27),
                           C2 => n163, ZN => n225);
   U142 : NAND2_X1 port map( A1 => n280, A2 => n279, ZN => Y(51));
   U143 : AOI222_X1 port map( A1 => A_shifted(51), A2 => n181, B1 => 
                           zeroSignal(51), B2 => n171, C1 => A_neg_shifted(51),
                           C2 => n161, ZN => n279);
   U144 : AOI22_X1 port map( A1 => A_neg(51), A2 => n154, B1 => A_signal(51), 
                           B2 => n145, ZN => n280);
   U145 : NAND2_X1 port map( A1 => n282, A2 => n281, ZN => Y(52));
   U146 : AOI222_X1 port map( A1 => A_shifted(52), A2 => n181, B1 => 
                           zeroSignal(52), B2 => n171, C1 => A_neg_shifted(52),
                           C2 => n161, ZN => n281);
   U147 : AOI22_X1 port map( A1 => A_neg(52), A2 => n154, B1 => A_signal(52), 
                           B2 => n145, ZN => n282);
   U148 : NAND2_X1 port map( A1 => n222, A2 => n221, ZN => Y(25));
   U149 : AOI222_X1 port map( A1 => A_shifted(25), A2 => n178, B1 => 
                           zeroSignal(25), B2 => n169, C1 => A_neg_shifted(25),
                           C2 => n163, ZN => n221);
   U150 : AOI22_X1 port map( A1 => A_neg(25), A2 => n152, B1 => A_signal(25), 
                           B2 => n143, ZN => n222);
   U151 : NAND2_X1 port map( A1 => n218, A2 => n217, ZN => Y(23));
   U152 : AOI222_X1 port map( A1 => A_shifted(23), A2 => n178, B1 => 
                           zeroSignal(23), B2 => n169, C1 => A_neg_shifted(23),
                           C2 => n164, ZN => n217);
   U153 : AOI22_X1 port map( A1 => A_neg(23), A2 => n152, B1 => A_signal(23), 
                           B2 => n143, ZN => n218);
   U154 : NAND2_X1 port map( A1 => n220, A2 => n219, ZN => Y(24));
   U155 : AOI222_X1 port map( A1 => A_shifted(24), A2 => n178, B1 => 
                           zeroSignal(24), B2 => n169, C1 => A_neg_shifted(24),
                           C2 => n163, ZN => n219);
   U156 : AOI22_X1 port map( A1 => A_neg(24), A2 => n152, B1 => A_signal(24), 
                           B2 => n143, ZN => n220);
   U157 : NAND2_X1 port map( A1 => n214, A2 => n213, ZN => Y(21));
   U158 : AOI222_X1 port map( A1 => A_shifted(21), A2 => n178, B1 => 
                           zeroSignal(21), B2 => n169, C1 => A_neg_shifted(21),
                           C2 => n164, ZN => n213);
   U159 : NAND2_X1 port map( A1 => n284, A2 => n283, ZN => Y(53));
   U160 : AOI222_X1 port map( A1 => A_shifted(53), A2 => n181, B1 => 
                           zeroSignal(53), B2 => n172, C1 => A_neg_shifted(53),
                           C2 => n161, ZN => n283);
   U161 : AOI22_X1 port map( A1 => A_neg(53), A2 => n155, B1 => A_signal(53), 
                           B2 => n146, ZN => n284);
   U162 : NAND2_X1 port map( A1 => n216, A2 => n215, ZN => Y(22));
   U163 : AOI222_X1 port map( A1 => A_shifted(22), A2 => n178, B1 => 
                           zeroSignal(22), B2 => n169, C1 => A_neg_shifted(22),
                           C2 => n164, ZN => n215);
   U164 : NAND2_X1 port map( A1 => n286, A2 => n285, ZN => Y(54));
   U165 : AOI22_X1 port map( A1 => A_neg(54), A2 => n155, B1 => A_signal(54), 
                           B2 => n146, ZN => n286);
   U166 : AOI222_X1 port map( A1 => A_shifted(54), A2 => n181, B1 => 
                           zeroSignal(54), B2 => n172, C1 => A_neg_shifted(54),
                           C2 => n161, ZN => n285);
   U167 : NAND2_X1 port map( A1 => n290, A2 => n289, ZN => Y(56));
   U168 : AOI222_X1 port map( A1 => A_shifted(56), A2 => n181, B1 => 
                           zeroSignal(56), B2 => n172, C1 => A_neg_shifted(56),
                           C2 => n161, ZN => n289);
   U169 : AOI22_X1 port map( A1 => A_neg(56), A2 => n155, B1 => A_signal(56), 
                           B2 => n146, ZN => n290);
   U170 : NAND2_X1 port map( A1 => n288, A2 => n287, ZN => Y(55));
   U171 : AOI22_X1 port map( A1 => A_neg(55), A2 => n155, B1 => A_signal(55), 
                           B2 => n146, ZN => n288);
   U172 : AOI222_X1 port map( A1 => A_shifted(55), A2 => n181, B1 => 
                           zeroSignal(55), B2 => n172, C1 => A_neg_shifted(55),
                           C2 => n161, ZN => n287);
   U173 : NAND2_X1 port map( A1 => n292, A2 => n291, ZN => Y(57));
   U174 : AOI22_X1 port map( A1 => A_neg(57), A2 => n155, B1 => A_signal(57), 
                           B2 => n146, ZN => n292);
   U175 : AOI222_X1 port map( A1 => A_shifted(57), A2 => n181, B1 => 
                           zeroSignal(57), B2 => n172, C1 => A_neg_shifted(57),
                           C2 => n160, ZN => n291);
   U176 : NAND2_X1 port map( A1 => n302, A2 => n301, ZN => Y(61));
   U177 : AOI222_X1 port map( A1 => A_shifted(61), A2 => n182, B1 => 
                           zeroSignal(61), B2 => n172, C1 => A_neg_shifted(61),
                           C2 => n160, ZN => n301);
   U178 : NAND2_X1 port map( A1 => n296, A2 => n295, ZN => Y(59));
   U179 : AOI22_X1 port map( A1 => A_neg(59), A2 => n155, B1 => A_signal(59), 
                           B2 => n146, ZN => n296);
   U180 : NAND2_X1 port map( A1 => n300, A2 => n299, ZN => Y(60));
   U181 : AOI222_X1 port map( A1 => A_shifted(60), A2 => n182, B1 => 
                           zeroSignal(60), B2 => n172, C1 => A_neg_shifted(60),
                           C2 => n160, ZN => n299);
   U182 : AOI22_X1 port map( A1 => A_neg(60), A2 => n155, B1 => A_signal(60), 
                           B2 => n146, ZN => n300);
   U183 : NAND2_X1 port map( A1 => n306, A2 => n305, ZN => Y(63));
   U184 : AOI222_X1 port map( A1 => A_shifted(63), A2 => n182, B1 => 
                           zeroSignal(63), B2 => n172, C1 => A_neg_shifted(63),
                           C2 => n160, ZN => n305);
   U185 : AOI22_X1 port map( A1 => A_neg(63), A2 => n155, B1 => A_signal(63), 
                           B2 => n146, ZN => n306);
   U186 : NAND2_X1 port map( A1 => n304, A2 => n303, ZN => Y(62));
   U187 : AOI22_X1 port map( A1 => A_neg(62), A2 => n155, B1 => A_signal(62), 
                           B2 => n146, ZN => n304);
   U188 : NAND2_X1 port map( A1 => n294, A2 => n293, ZN => Y(58));
   U189 : AOI222_X1 port map( A1 => A_shifted(58), A2 => n181, B1 => 
                           zeroSignal(58), B2 => n172, C1 => A_neg_shifted(58),
                           C2 => n160, ZN => n293);
   U190 : NAND2_X1 port map( A1 => n188, A2 => n187, ZN => Y(0));
   U191 : AOI22_X1 port map( A1 => A_neg(0), A2 => n151, B1 => A_signal(0), B2 
                           => n142, ZN => n188);
   U192 : AOI222_X1 port map( A1 => A_shifted(0), A2 => n177, B1 => 
                           zeroSignal(0), B2 => n168, C1 => A_neg_shifted(0), 
                           C2 => n165, ZN => n187);
   U193 : NAND2_X1 port map( A1 => n210, A2 => n209, ZN => Y(1));
   U194 : AOI22_X1 port map( A1 => A_neg(1), A2 => n151, B1 => A_signal(1), B2 
                           => n142, ZN => n210);
   U195 : AOI222_X1 port map( A1 => A_shifted(1), A2 => n178, B1 => 
                           zeroSignal(1), B2 => n168, C1 => A_neg_shifted(1), 
                           C2 => n164, ZN => n209);
   U196 : NAND2_X1 port map( A1 => n232, A2 => n231, ZN => Y(2));
   U197 : AOI22_X1 port map( A1 => A_neg(2), A2 => n152, B1 => A_signal(2), B2 
                           => n143, ZN => n232);
   U198 : AOI222_X1 port map( A1 => A_shifted(2), A2 => n179, B1 => 
                           zeroSignal(2), B2 => n169, C1 => A_neg_shifted(2), 
                           C2 => n163, ZN => n231);
   U199 : NAND2_X1 port map( A1 => n254, A2 => n253, ZN => Y(3));
   U200 : AOI22_X1 port map( A1 => A_neg(3), A2 => n153, B1 => A_signal(3), B2 
                           => n144, ZN => n254);
   U201 : AOI222_X1 port map( A1 => A_shifted(3), A2 => n180, B1 => 
                           zeroSignal(3), B2 => n170, C1 => A_neg_shifted(3), 
                           C2 => n162, ZN => n253);
   U202 : NAND2_X1 port map( A1 => n276, A2 => n275, ZN => Y(4));
   U203 : AOI22_X1 port map( A1 => A_neg(4), A2 => n154, B1 => A_signal(4), B2 
                           => n145, ZN => n276);
   U204 : AOI222_X1 port map( A1 => A_shifted(4), A2 => n181, B1 => 
                           zeroSignal(4), B2 => n171, C1 => A_neg_shifted(4), 
                           C2 => n161, ZN => n275);
   U205 : NAND2_X1 port map( A1 => n298, A2 => n297, ZN => Y(5));
   U206 : AOI22_X1 port map( A1 => A_neg(5), A2 => n155, B1 => A_signal(5), B2 
                           => n146, ZN => n298);
   U207 : AOI222_X1 port map( A1 => A_shifted(5), A2 => n182, B1 => 
                           zeroSignal(5), B2 => n172, C1 => A_neg_shifted(5), 
                           C2 => n160, ZN => n297);
   U208 : NAND2_X1 port map( A1 => n308, A2 => n307, ZN => Y(6));
   U209 : AOI22_X1 port map( A1 => A_neg(6), A2 => n156, B1 => A_signal(6), B2 
                           => n147, ZN => n308);
   U210 : AOI222_X1 port map( A1 => A_shifted(6), A2 => n182, B1 => 
                           zeroSignal(6), B2 => n173, C1 => A_neg_shifted(6), 
                           C2 => n160, ZN => n307);
   U211 : NAND2_X1 port map( A1 => n310, A2 => n309, ZN => Y(7));
   U212 : AOI22_X1 port map( A1 => A_neg(7), A2 => n156, B1 => A_signal(7), B2 
                           => n147, ZN => n310);
   U213 : AOI222_X1 port map( A1 => A_shifted(7), A2 => n182, B1 => 
                           zeroSignal(7), B2 => n173, C1 => A_neg_shifted(7), 
                           C2 => n160, ZN => n309);
   U214 : NAND2_X1 port map( A1 => n312, A2 => n311, ZN => Y(8));
   U215 : AOI22_X1 port map( A1 => A_neg(8), A2 => n156, B1 => A_signal(8), B2 
                           => n147, ZN => n312);
   U216 : AOI222_X1 port map( A1 => A_shifted(8), A2 => n182, B1 => 
                           zeroSignal(8), B2 => n173, C1 => A_neg_shifted(8), 
                           C2 => n160, ZN => n311);
   U217 : NAND2_X1 port map( A1 => n318, A2 => n317, ZN => Y(9));
   U218 : AOI22_X1 port map( A1 => A_neg(9), A2 => n156, B1 => A_signal(9), B2 
                           => n147, ZN => n318);
   U219 : AOI222_X1 port map( A1 => A_shifted(9), A2 => n182, B1 => 
                           zeroSignal(9), B2 => n173, C1 => A_neg_shifted(9), 
                           C2 => n160, ZN => n317);
   U220 : NAND2_X1 port map( A1 => n190, A2 => n189, ZN => Y(10));
   U221 : AOI22_X1 port map( A1 => A_neg(10), A2 => n151, B1 => A_signal(10), 
                           B2 => n142, ZN => n190);
   U222 : AOI222_X1 port map( A1 => A_shifted(10), A2 => n177, B1 => 
                           zeroSignal(10), B2 => n168, C1 => A_neg_shifted(10),
                           C2 => n165, ZN => n189);
   U223 : NAND2_X1 port map( A1 => n192, A2 => n191, ZN => Y(11));
   U224 : AOI22_X1 port map( A1 => A_neg(11), A2 => n151, B1 => A_signal(11), 
                           B2 => n142, ZN => n192);
   U225 : AOI222_X1 port map( A1 => A_shifted(11), A2 => n177, B1 => 
                           zeroSignal(11), B2 => n168, C1 => A_neg_shifted(11),
                           C2 => n165, ZN => n191);
   U226 : NAND2_X1 port map( A1 => n194, A2 => n193, ZN => Y(12));
   U227 : AOI22_X1 port map( A1 => A_neg(12), A2 => n151, B1 => A_signal(12), 
                           B2 => n142, ZN => n194);
   U228 : AOI222_X1 port map( A1 => A_shifted(12), A2 => n177, B1 => 
                           zeroSignal(12), B2 => n168, C1 => A_neg_shifted(12),
                           C2 => n165, ZN => n193);
   U229 : NAND2_X1 port map( A1 => n196, A2 => n195, ZN => Y(13));
   U230 : AOI22_X1 port map( A1 => A_neg(13), A2 => n151, B1 => A_signal(13), 
                           B2 => n142, ZN => n196);
   U231 : AOI222_X1 port map( A1 => A_shifted(13), A2 => n177, B1 => 
                           zeroSignal(13), B2 => n168, C1 => A_neg_shifted(13),
                           C2 => n164, ZN => n195);
   U232 : NAND2_X1 port map( A1 => n198, A2 => n197, ZN => Y(14));
   U233 : AOI22_X1 port map( A1 => A_neg(14), A2 => n151, B1 => A_signal(14), 
                           B2 => n142, ZN => n198);
   U234 : AOI222_X1 port map( A1 => A_shifted(14), A2 => n177, B1 => 
                           zeroSignal(14), B2 => n168, C1 => A_neg_shifted(14),
                           C2 => n164, ZN => n197);
   U235 : NAND2_X1 port map( A1 => n200, A2 => n199, ZN => Y(15));
   U236 : AOI22_X1 port map( A1 => A_neg(15), A2 => n151, B1 => A_signal(15), 
                           B2 => n142, ZN => n200);
   U237 : AOI222_X1 port map( A1 => A_shifted(15), A2 => n177, B1 => 
                           zeroSignal(15), B2 => n168, C1 => A_neg_shifted(15),
                           C2 => n164, ZN => n199);
   U238 : AOI22_X1 port map( A1 => A_neg(22), A2 => n152, B1 => A_signal(22), 
                           B2 => n143, ZN => n216);
   U239 : AOI22_X1 port map( A1 => A_neg(21), A2 => n152, B1 => A_signal(21), 
                           B2 => n143, ZN => n214);
   U240 : AOI22_X1 port map( A1 => A_neg(19), A2 => n151, B1 => A_signal(19), 
                           B2 => n142, ZN => n208);
   U241 : AOI222_X1 port map( A1 => A_shifted(62), A2 => n182, B1 => 
                           zeroSignal(62), B2 => n172, C1 => A_neg_shifted(62),
                           C2 => n160, ZN => n303);
   U242 : AOI22_X1 port map( A1 => A_neg(61), A2 => n155, B1 => A_signal(61), 
                           B2 => n146, ZN => n302);
   U243 : AOI222_X1 port map( A1 => A_shifted(59), A2 => n181, B1 => 
                           zeroSignal(59), B2 => n172, C1 => A_neg_shifted(59),
                           C2 => n160, ZN => n295);
   U244 : AOI22_X1 port map( A1 => A_neg(58), A2 => n155, B1 => A_signal(58), 
                           B2 => n146, ZN => n294);

end SYN_BEHAVIORAL_2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity MUX51_MuxNbit64_7 is

   port( zeroSignal, A_signal, A_neg, A_shifted, A_neg_shifted : in 
         std_logic_vector (63 downto 0);  Sel : in std_logic_vector (2 downto 
         0);  Y : out std_logic_vector (63 downto 0));

end MUX51_MuxNbit64_7;

architecture SYN_BEHAVIORAL_2 of MUX51_MuxNbit64_7 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, 
      n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, 
      n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, 
      n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, 
      n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, 
      n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, 
      n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, 
      n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, 
      n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, 
      n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, 
      n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, 
      n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, 
      n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, 
      n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, 
      n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, 
      n320 : std_logic;

begin
   
   U1 : AND3_X1 port map( A1 => n319, A2 => n320, A3 => Sel(2), ZN => n141);
   U2 : BUF_X1 port map( A => n141, Z => n166);
   U3 : BUF_X1 port map( A => n159, Z => n158);
   U4 : BUF_X1 port map( A => n185, Z => n184);
   U5 : BUF_X1 port map( A => n150, Z => n149);
   U6 : BUF_X1 port map( A => n141, Z => n167);
   U7 : BUF_X1 port map( A => n185, Z => n183);
   U8 : BUF_X1 port map( A => n159, Z => n157);
   U9 : BUF_X1 port map( A => n150, Z => n148);
   U10 : BUF_X1 port map( A => n176, Z => n175);
   U11 : BUF_X1 port map( A => n176, Z => n174);
   U12 : BUF_X1 port map( A => n184, Z => n177);
   U13 : BUF_X1 port map( A => n158, Z => n151);
   U14 : BUF_X1 port map( A => n149, Z => n142);
   U15 : BUF_X1 port map( A => n166, Z => n164);
   U16 : BUF_X1 port map( A => n184, Z => n178);
   U17 : BUF_X1 port map( A => n158, Z => n152);
   U18 : BUF_X1 port map( A => n149, Z => n143);
   U19 : BUF_X1 port map( A => n166, Z => n163);
   U20 : BUF_X1 port map( A => n184, Z => n179);
   U21 : BUF_X1 port map( A => n158, Z => n153);
   U22 : BUF_X1 port map( A => n149, Z => n144);
   U23 : BUF_X1 port map( A => n167, Z => n162);
   U24 : BUF_X1 port map( A => n183, Z => n180);
   U25 : BUF_X1 port map( A => n157, Z => n154);
   U26 : BUF_X1 port map( A => n148, Z => n145);
   U27 : BUF_X1 port map( A => n167, Z => n161);
   U28 : BUF_X1 port map( A => n183, Z => n181);
   U29 : BUF_X1 port map( A => n157, Z => n155);
   U30 : BUF_X1 port map( A => n148, Z => n146);
   U31 : BUF_X1 port map( A => n167, Z => n160);
   U32 : BUF_X1 port map( A => n183, Z => n182);
   U33 : BUF_X1 port map( A => n175, Z => n168);
   U34 : BUF_X1 port map( A => n175, Z => n169);
   U35 : BUF_X1 port map( A => n175, Z => n170);
   U36 : BUF_X1 port map( A => n174, Z => n171);
   U37 : BUF_X1 port map( A => n174, Z => n172);
   U38 : BUF_X1 port map( A => n166, Z => n165);
   U39 : BUF_X1 port map( A => n157, Z => n156);
   U40 : BUF_X1 port map( A => n148, Z => n147);
   U41 : BUF_X1 port map( A => n174, Z => n173);
   U42 : INV_X1 port map( A => Sel(1), ZN => n320);
   U43 : BUF_X1 port map( A => n316, Z => n185);
   U44 : NOR3_X1 port map( A1 => n319, A2 => Sel(2), A3 => n320, ZN => n316);
   U45 : BUF_X1 port map( A => n314, Z => n159);
   U46 : NOR3_X1 port map( A1 => Sel(0), A2 => Sel(2), A3 => n320, ZN => n314);
   U47 : INV_X1 port map( A => Sel(0), ZN => n319);
   U48 : BUF_X1 port map( A => n313, Z => n150);
   U49 : NOR3_X1 port map( A1 => Sel(1), A2 => Sel(2), A3 => n319, ZN => n313);
   U50 : BUF_X1 port map( A => n315, Z => n176);
   U51 : NOR2_X1 port map( A1 => n165, A2 => n186, ZN => n315);
   U52 : AOI21_X1 port map( B1 => n319, B2 => n320, A => Sel(2), ZN => n186);
   U53 : NAND2_X1 port map( A1 => n208, A2 => n207, ZN => Y(19));
   U54 : AOI22_X1 port map( A1 => A_neg(19), A2 => n151, B1 => A_signal(19), B2
                           => n142, ZN => n208);
   U55 : AOI222_X1 port map( A1 => A_shifted(19), A2 => n177, B1 => 
                           zeroSignal(19), B2 => n168, C1 => A_neg_shifted(19),
                           C2 => n164, ZN => n207);
   U56 : NAND2_X1 port map( A1 => n206, A2 => n205, ZN => Y(18));
   U57 : AOI222_X1 port map( A1 => A_shifted(18), A2 => n177, B1 => 
                           zeroSignal(18), B2 => n168, C1 => A_neg_shifted(18),
                           C2 => n164, ZN => n205);
   U58 : AOI22_X1 port map( A1 => A_neg(18), A2 => n151, B1 => A_signal(18), B2
                           => n142, ZN => n206);
   U59 : NAND2_X1 port map( A1 => n240, A2 => n239, ZN => Y(33));
   U60 : AOI222_X1 port map( A1 => A_shifted(33), A2 => n179, B1 => 
                           zeroSignal(33), B2 => n170, C1 => A_neg_shifted(33),
                           C2 => n163, ZN => n239);
   U61 : AOI22_X1 port map( A1 => A_neg(33), A2 => n153, B1 => A_signal(33), B2
                           => n144, ZN => n240);
   U62 : NAND2_X1 port map( A1 => n236, A2 => n235, ZN => Y(31));
   U63 : AOI222_X1 port map( A1 => A_shifted(31), A2 => n179, B1 => 
                           zeroSignal(31), B2 => n170, C1 => A_neg_shifted(31),
                           C2 => n163, ZN => n235);
   U64 : AOI22_X1 port map( A1 => A_neg(31), A2 => n153, B1 => A_signal(31), B2
                           => n144, ZN => n236);
   U65 : NAND2_X1 port map( A1 => n238, A2 => n237, ZN => Y(32));
   U66 : AOI222_X1 port map( A1 => A_shifted(32), A2 => n179, B1 => 
                           zeroSignal(32), B2 => n170, C1 => A_neg_shifted(32),
                           C2 => n163, ZN => n237);
   U67 : AOI22_X1 port map( A1 => A_neg(32), A2 => n153, B1 => A_signal(32), B2
                           => n144, ZN => n238);
   U68 : NAND2_X1 port map( A1 => n242, A2 => n241, ZN => Y(34));
   U69 : AOI222_X1 port map( A1 => A_shifted(34), A2 => n179, B1 => 
                           zeroSignal(34), B2 => n170, C1 => A_neg_shifted(34),
                           C2 => n163, ZN => n241);
   U70 : AOI22_X1 port map( A1 => A_neg(34), A2 => n153, B1 => A_signal(34), B2
                           => n144, ZN => n242);
   U71 : NAND2_X1 port map( A1 => n212, A2 => n211, ZN => Y(20));
   U72 : AOI22_X1 port map( A1 => A_neg(20), A2 => n152, B1 => A_signal(20), B2
                           => n143, ZN => n212);
   U73 : AOI222_X1 port map( A1 => A_shifted(20), A2 => n178, B1 => 
                           zeroSignal(20), B2 => n169, C1 => A_neg_shifted(20),
                           C2 => n164, ZN => n211);
   U74 : NAND2_X1 port map( A1 => n244, A2 => n243, ZN => Y(35));
   U75 : AOI222_X1 port map( A1 => A_shifted(35), A2 => n179, B1 => 
                           zeroSignal(35), B2 => n170, C1 => A_neg_shifted(35),
                           C2 => n162, ZN => n243);
   U76 : AOI22_X1 port map( A1 => A_neg(35), A2 => n153, B1 => A_signal(35), B2
                           => n144, ZN => n244);
   U77 : NAND2_X1 port map( A1 => n248, A2 => n247, ZN => Y(37));
   U78 : AOI222_X1 port map( A1 => A_shifted(37), A2 => n179, B1 => 
                           zeroSignal(37), B2 => n170, C1 => A_neg_shifted(37),
                           C2 => n162, ZN => n247);
   U79 : AOI22_X1 port map( A1 => A_neg(37), A2 => n153, B1 => A_signal(37), B2
                           => n144, ZN => n248);
   U80 : NAND2_X1 port map( A1 => n250, A2 => n249, ZN => Y(38));
   U81 : AOI222_X1 port map( A1 => A_shifted(38), A2 => n179, B1 => 
                           zeroSignal(38), B2 => n170, C1 => A_neg_shifted(38),
                           C2 => n162, ZN => n249);
   U82 : AOI22_X1 port map( A1 => A_neg(38), A2 => n153, B1 => A_signal(38), B2
                           => n144, ZN => n250);
   U83 : NAND2_X1 port map( A1 => n252, A2 => n251, ZN => Y(39));
   U84 : AOI222_X1 port map( A1 => A_shifted(39), A2 => n179, B1 => 
                           zeroSignal(39), B2 => n170, C1 => A_neg_shifted(39),
                           C2 => n162, ZN => n251);
   U85 : AOI22_X1 port map( A1 => A_neg(39), A2 => n153, B1 => A_signal(39), B2
                           => n144, ZN => n252);
   U86 : NAND2_X1 port map( A1 => n256, A2 => n255, ZN => Y(40));
   U87 : AOI222_X1 port map( A1 => A_shifted(40), A2 => n180, B1 => 
                           zeroSignal(40), B2 => n170, C1 => A_neg_shifted(40),
                           C2 => n162, ZN => n255);
   U88 : AOI22_X1 port map( A1 => A_neg(40), A2 => n153, B1 => A_signal(40), B2
                           => n144, ZN => n256);
   U89 : NAND2_X1 port map( A1 => n258, A2 => n257, ZN => Y(41));
   U90 : AOI222_X1 port map( A1 => A_shifted(41), A2 => n180, B1 => 
                           zeroSignal(41), B2 => n170, C1 => A_neg_shifted(41),
                           C2 => n162, ZN => n257);
   U91 : AOI22_X1 port map( A1 => A_neg(41), A2 => n153, B1 => A_signal(41), B2
                           => n144, ZN => n258);
   U92 : NAND2_X1 port map( A1 => n260, A2 => n259, ZN => Y(42));
   U93 : AOI222_X1 port map( A1 => A_shifted(42), A2 => n180, B1 => 
                           zeroSignal(42), B2 => n171, C1 => A_neg_shifted(42),
                           C2 => n162, ZN => n259);
   U94 : AOI22_X1 port map( A1 => A_neg(42), A2 => n154, B1 => A_signal(42), B2
                           => n145, ZN => n260);
   U95 : NAND2_X1 port map( A1 => n262, A2 => n261, ZN => Y(43));
   U96 : AOI222_X1 port map( A1 => A_shifted(43), A2 => n180, B1 => 
                           zeroSignal(43), B2 => n171, C1 => A_neg_shifted(43),
                           C2 => n162, ZN => n261);
   U97 : AOI22_X1 port map( A1 => A_neg(43), A2 => n154, B1 => A_signal(43), B2
                           => n145, ZN => n262);
   U98 : NAND2_X1 port map( A1 => n264, A2 => n263, ZN => Y(44));
   U99 : AOI222_X1 port map( A1 => A_shifted(44), A2 => n180, B1 => 
                           zeroSignal(44), B2 => n171, C1 => A_neg_shifted(44),
                           C2 => n162, ZN => n263);
   U100 : AOI22_X1 port map( A1 => A_neg(44), A2 => n154, B1 => A_signal(44), 
                           B2 => n145, ZN => n264);
   U101 : NAND2_X1 port map( A1 => n266, A2 => n265, ZN => Y(45));
   U102 : AOI222_X1 port map( A1 => A_shifted(45), A2 => n180, B1 => 
                           zeroSignal(45), B2 => n171, C1 => A_neg_shifted(45),
                           C2 => n162, ZN => n265);
   U103 : AOI22_X1 port map( A1 => A_neg(45), A2 => n154, B1 => A_signal(45), 
                           B2 => n145, ZN => n266);
   U104 : NAND2_X1 port map( A1 => n268, A2 => n267, ZN => Y(46));
   U105 : AOI222_X1 port map( A1 => A_shifted(46), A2 => n180, B1 => 
                           zeroSignal(46), B2 => n171, C1 => A_neg_shifted(46),
                           C2 => n161, ZN => n267);
   U106 : AOI22_X1 port map( A1 => A_neg(46), A2 => n154, B1 => A_signal(46), 
                           B2 => n145, ZN => n268);
   U107 : NAND2_X1 port map( A1 => n246, A2 => n245, ZN => Y(36));
   U108 : AOI22_X1 port map( A1 => A_neg(36), A2 => n153, B1 => A_signal(36), 
                           B2 => n144, ZN => n246);
   U109 : AOI222_X1 port map( A1 => A_shifted(36), A2 => n179, B1 => 
                           zeroSignal(36), B2 => n170, C1 => A_neg_shifted(36),
                           C2 => n162, ZN => n245);
   U110 : NAND2_X1 port map( A1 => n272, A2 => n271, ZN => Y(48));
   U111 : AOI222_X1 port map( A1 => A_shifted(48), A2 => n180, B1 => 
                           zeroSignal(48), B2 => n171, C1 => A_neg_shifted(48),
                           C2 => n161, ZN => n271);
   U112 : AOI22_X1 port map( A1 => A_neg(48), A2 => n154, B1 => A_signal(48), 
                           B2 => n145, ZN => n272);
   U113 : NAND2_X1 port map( A1 => n214, A2 => n213, ZN => Y(21));
   U114 : AOI222_X1 port map( A1 => A_shifted(21), A2 => n178, B1 => 
                           zeroSignal(21), B2 => n169, C1 => A_neg_shifted(21),
                           C2 => n164, ZN => n213);
   U115 : NAND2_X1 port map( A1 => n274, A2 => n273, ZN => Y(49));
   U116 : AOI222_X1 port map( A1 => A_shifted(49), A2 => n180, B1 => 
                           zeroSignal(49), B2 => n171, C1 => A_neg_shifted(49),
                           C2 => n161, ZN => n273);
   U117 : AOI22_X1 port map( A1 => A_neg(49), A2 => n154, B1 => A_signal(49), 
                           B2 => n145, ZN => n274);
   U118 : NAND2_X1 port map( A1 => n278, A2 => n277, ZN => Y(50));
   U119 : AOI222_X1 port map( A1 => A_shifted(50), A2 => n181, B1 => 
                           zeroSignal(50), B2 => n171, C1 => A_neg_shifted(50),
                           C2 => n161, ZN => n277);
   U120 : AOI22_X1 port map( A1 => A_neg(50), A2 => n154, B1 => A_signal(50), 
                           B2 => n145, ZN => n278);
   U121 : NAND2_X1 port map( A1 => n280, A2 => n279, ZN => Y(51));
   U122 : AOI222_X1 port map( A1 => A_shifted(51), A2 => n181, B1 => 
                           zeroSignal(51), B2 => n171, C1 => A_neg_shifted(51),
                           C2 => n161, ZN => n279);
   U123 : AOI22_X1 port map( A1 => A_neg(51), A2 => n154, B1 => A_signal(51), 
                           B2 => n145, ZN => n280);
   U124 : NAND2_X1 port map( A1 => n270, A2 => n269, ZN => Y(47));
   U125 : AOI22_X1 port map( A1 => A_neg(47), A2 => n154, B1 => A_signal(47), 
                           B2 => n145, ZN => n270);
   U126 : AOI222_X1 port map( A1 => A_shifted(47), A2 => n180, B1 => 
                           zeroSignal(47), B2 => n171, C1 => A_neg_shifted(47),
                           C2 => n161, ZN => n269);
   U127 : NAND2_X1 port map( A1 => n228, A2 => n227, ZN => Y(28));
   U128 : AOI222_X1 port map( A1 => A_shifted(28), A2 => n178, B1 => 
                           zeroSignal(28), B2 => n169, C1 => A_neg_shifted(28),
                           C2 => n163, ZN => n227);
   U129 : AOI22_X1 port map( A1 => A_neg(28), A2 => n152, B1 => A_signal(28), 
                           B2 => n143, ZN => n228);
   U130 : NAND2_X1 port map( A1 => n216, A2 => n215, ZN => Y(22));
   U131 : AOI22_X1 port map( A1 => A_neg(22), A2 => n152, B1 => A_signal(22), 
                           B2 => n143, ZN => n216);
   U132 : AOI222_X1 port map( A1 => A_shifted(22), A2 => n178, B1 => 
                           zeroSignal(22), B2 => n169, C1 => A_neg_shifted(22),
                           C2 => n164, ZN => n215);
   U133 : NAND2_X1 port map( A1 => n234, A2 => n233, ZN => Y(30));
   U134 : AOI222_X1 port map( A1 => A_shifted(30), A2 => n179, B1 => 
                           zeroSignal(30), B2 => n169, C1 => A_neg_shifted(30),
                           C2 => n163, ZN => n233);
   U135 : AOI22_X1 port map( A1 => A_neg(30), A2 => n152, B1 => A_signal(30), 
                           B2 => n143, ZN => n234);
   U136 : NAND2_X1 port map( A1 => n282, A2 => n281, ZN => Y(52));
   U137 : AOI222_X1 port map( A1 => A_shifted(52), A2 => n181, B1 => 
                           zeroSignal(52), B2 => n171, C1 => A_neg_shifted(52),
                           C2 => n161, ZN => n281);
   U138 : AOI22_X1 port map( A1 => A_neg(52), A2 => n154, B1 => A_signal(52), 
                           B2 => n145, ZN => n282);
   U139 : NAND2_X1 port map( A1 => n230, A2 => n229, ZN => Y(29));
   U140 : AOI22_X1 port map( A1 => A_neg(29), A2 => n152, B1 => A_signal(29), 
                           B2 => n143, ZN => n230);
   U141 : AOI222_X1 port map( A1 => A_shifted(29), A2 => n178, B1 => 
                           zeroSignal(29), B2 => n169, C1 => A_neg_shifted(29),
                           C2 => n163, ZN => n229);
   U142 : NAND2_X1 port map( A1 => n284, A2 => n283, ZN => Y(53));
   U143 : AOI222_X1 port map( A1 => A_shifted(53), A2 => n181, B1 => 
                           zeroSignal(53), B2 => n172, C1 => A_neg_shifted(53),
                           C2 => n161, ZN => n283);
   U144 : AOI22_X1 port map( A1 => A_neg(53), A2 => n155, B1 => A_signal(53), 
                           B2 => n146, ZN => n284);
   U145 : NAND2_X1 port map( A1 => n286, A2 => n285, ZN => Y(54));
   U146 : AOI222_X1 port map( A1 => A_shifted(54), A2 => n181, B1 => 
                           zeroSignal(54), B2 => n172, C1 => A_neg_shifted(54),
                           C2 => n161, ZN => n285);
   U147 : AOI22_X1 port map( A1 => A_neg(54), A2 => n155, B1 => A_signal(54), 
                           B2 => n146, ZN => n286);
   U148 : NAND2_X1 port map( A1 => n226, A2 => n225, ZN => Y(27));
   U149 : AOI222_X1 port map( A1 => A_shifted(27), A2 => n178, B1 => 
                           zeroSignal(27), B2 => n169, C1 => A_neg_shifted(27),
                           C2 => n163, ZN => n225);
   U150 : AOI22_X1 port map( A1 => A_neg(27), A2 => n152, B1 => A_signal(27), 
                           B2 => n143, ZN => n226);
   U151 : NAND2_X1 port map( A1 => n222, A2 => n221, ZN => Y(25));
   U152 : AOI222_X1 port map( A1 => A_shifted(25), A2 => n178, B1 => 
                           zeroSignal(25), B2 => n169, C1 => A_neg_shifted(25),
                           C2 => n163, ZN => n221);
   U153 : AOI22_X1 port map( A1 => A_neg(25), A2 => n152, B1 => A_signal(25), 
                           B2 => n143, ZN => n222);
   U154 : NAND2_X1 port map( A1 => n224, A2 => n223, ZN => Y(26));
   U155 : AOI222_X1 port map( A1 => A_shifted(26), A2 => n178, B1 => 
                           zeroSignal(26), B2 => n169, C1 => A_neg_shifted(26),
                           C2 => n163, ZN => n223);
   U156 : AOI22_X1 port map( A1 => A_neg(26), A2 => n152, B1 => A_signal(26), 
                           B2 => n143, ZN => n224);
   U157 : NAND2_X1 port map( A1 => n218, A2 => n217, ZN => Y(23));
   U158 : AOI222_X1 port map( A1 => A_shifted(23), A2 => n178, B1 => 
                           zeroSignal(23), B2 => n169, C1 => A_neg_shifted(23),
                           C2 => n164, ZN => n217);
   U159 : NAND2_X1 port map( A1 => n288, A2 => n287, ZN => Y(55));
   U160 : AOI222_X1 port map( A1 => A_shifted(55), A2 => n181, B1 => 
                           zeroSignal(55), B2 => n172, C1 => A_neg_shifted(55),
                           C2 => n161, ZN => n287);
   U161 : AOI22_X1 port map( A1 => A_neg(55), A2 => n155, B1 => A_signal(55), 
                           B2 => n146, ZN => n288);
   U162 : NAND2_X1 port map( A1 => n220, A2 => n219, ZN => Y(24));
   U163 : AOI222_X1 port map( A1 => A_shifted(24), A2 => n178, B1 => 
                           zeroSignal(24), B2 => n169, C1 => A_neg_shifted(24),
                           C2 => n163, ZN => n219);
   U164 : NAND2_X1 port map( A1 => n290, A2 => n289, ZN => Y(56));
   U165 : AOI22_X1 port map( A1 => A_neg(56), A2 => n155, B1 => A_signal(56), 
                           B2 => n146, ZN => n290);
   U166 : AOI222_X1 port map( A1 => A_shifted(56), A2 => n181, B1 => 
                           zeroSignal(56), B2 => n172, C1 => A_neg_shifted(56),
                           C2 => n161, ZN => n289);
   U167 : NAND2_X1 port map( A1 => n294, A2 => n293, ZN => Y(58));
   U168 : AOI222_X1 port map( A1 => A_shifted(58), A2 => n181, B1 => 
                           zeroSignal(58), B2 => n172, C1 => A_neg_shifted(58),
                           C2 => n160, ZN => n293);
   U169 : AOI22_X1 port map( A1 => A_neg(58), A2 => n155, B1 => A_signal(58), 
                           B2 => n146, ZN => n294);
   U170 : NAND2_X1 port map( A1 => n292, A2 => n291, ZN => Y(57));
   U171 : AOI22_X1 port map( A1 => A_neg(57), A2 => n155, B1 => A_signal(57), 
                           B2 => n146, ZN => n292);
   U172 : AOI222_X1 port map( A1 => A_shifted(57), A2 => n181, B1 => 
                           zeroSignal(57), B2 => n172, C1 => A_neg_shifted(57),
                           C2 => n160, ZN => n291);
   U173 : NAND2_X1 port map( A1 => n296, A2 => n295, ZN => Y(59));
   U174 : AOI22_X1 port map( A1 => A_neg(59), A2 => n155, B1 => A_signal(59), 
                           B2 => n146, ZN => n296);
   U175 : AOI222_X1 port map( A1 => A_shifted(59), A2 => n181, B1 => 
                           zeroSignal(59), B2 => n172, C1 => A_neg_shifted(59),
                           C2 => n160, ZN => n295);
   U176 : NAND2_X1 port map( A1 => n306, A2 => n305, ZN => Y(63));
   U177 : AOI222_X1 port map( A1 => A_shifted(63), A2 => n182, B1 => 
                           zeroSignal(63), B2 => n172, C1 => A_neg_shifted(63),
                           C2 => n160, ZN => n305);
   U178 : NAND2_X1 port map( A1 => n304, A2 => n303, ZN => Y(62));
   U179 : AOI222_X1 port map( A1 => A_shifted(62), A2 => n182, B1 => 
                           zeroSignal(62), B2 => n172, C1 => A_neg_shifted(62),
                           C2 => n160, ZN => n303);
   U180 : AOI22_X1 port map( A1 => A_neg(62), A2 => n155, B1 => A_signal(62), 
                           B2 => n146, ZN => n304);
   U181 : NAND2_X1 port map( A1 => n302, A2 => n301, ZN => Y(61));
   U182 : AOI22_X1 port map( A1 => A_neg(61), A2 => n155, B1 => A_signal(61), 
                           B2 => n146, ZN => n302);
   U183 : NAND2_X1 port map( A1 => n300, A2 => n299, ZN => Y(60));
   U184 : AOI222_X1 port map( A1 => A_shifted(60), A2 => n182, B1 => 
                           zeroSignal(60), B2 => n172, C1 => A_neg_shifted(60),
                           C2 => n160, ZN => n299);
   U185 : NAND2_X1 port map( A1 => n188, A2 => n187, ZN => Y(0));
   U186 : AOI22_X1 port map( A1 => A_neg(0), A2 => n151, B1 => A_signal(0), B2 
                           => n142, ZN => n188);
   U187 : AOI222_X1 port map( A1 => A_shifted(0), A2 => n177, B1 => 
                           zeroSignal(0), B2 => n168, C1 => A_neg_shifted(0), 
                           C2 => n165, ZN => n187);
   U188 : NAND2_X1 port map( A1 => n210, A2 => n209, ZN => Y(1));
   U189 : AOI22_X1 port map( A1 => A_neg(1), A2 => n151, B1 => A_signal(1), B2 
                           => n142, ZN => n210);
   U190 : AOI222_X1 port map( A1 => A_shifted(1), A2 => n178, B1 => 
                           zeroSignal(1), B2 => n168, C1 => A_neg_shifted(1), 
                           C2 => n164, ZN => n209);
   U191 : NAND2_X1 port map( A1 => n232, A2 => n231, ZN => Y(2));
   U192 : AOI22_X1 port map( A1 => A_neg(2), A2 => n152, B1 => A_signal(2), B2 
                           => n143, ZN => n232);
   U193 : AOI222_X1 port map( A1 => A_shifted(2), A2 => n179, B1 => 
                           zeroSignal(2), B2 => n169, C1 => A_neg_shifted(2), 
                           C2 => n163, ZN => n231);
   U194 : NAND2_X1 port map( A1 => n254, A2 => n253, ZN => Y(3));
   U195 : AOI22_X1 port map( A1 => A_neg(3), A2 => n153, B1 => A_signal(3), B2 
                           => n144, ZN => n254);
   U196 : AOI222_X1 port map( A1 => A_shifted(3), A2 => n180, B1 => 
                           zeroSignal(3), B2 => n170, C1 => A_neg_shifted(3), 
                           C2 => n162, ZN => n253);
   U197 : NAND2_X1 port map( A1 => n276, A2 => n275, ZN => Y(4));
   U198 : AOI22_X1 port map( A1 => A_neg(4), A2 => n154, B1 => A_signal(4), B2 
                           => n145, ZN => n276);
   U199 : AOI222_X1 port map( A1 => A_shifted(4), A2 => n181, B1 => 
                           zeroSignal(4), B2 => n171, C1 => A_neg_shifted(4), 
                           C2 => n161, ZN => n275);
   U200 : NAND2_X1 port map( A1 => n298, A2 => n297, ZN => Y(5));
   U201 : AOI22_X1 port map( A1 => A_neg(5), A2 => n155, B1 => A_signal(5), B2 
                           => n146, ZN => n298);
   U202 : AOI222_X1 port map( A1 => A_shifted(5), A2 => n182, B1 => 
                           zeroSignal(5), B2 => n172, C1 => A_neg_shifted(5), 
                           C2 => n160, ZN => n297);
   U203 : NAND2_X1 port map( A1 => n308, A2 => n307, ZN => Y(6));
   U204 : AOI22_X1 port map( A1 => A_neg(6), A2 => n156, B1 => A_signal(6), B2 
                           => n147, ZN => n308);
   U205 : AOI222_X1 port map( A1 => A_shifted(6), A2 => n182, B1 => 
                           zeroSignal(6), B2 => n173, C1 => A_neg_shifted(6), 
                           C2 => n160, ZN => n307);
   U206 : NAND2_X1 port map( A1 => n310, A2 => n309, ZN => Y(7));
   U207 : AOI22_X1 port map( A1 => A_neg(7), A2 => n156, B1 => A_signal(7), B2 
                           => n147, ZN => n310);
   U208 : AOI222_X1 port map( A1 => A_shifted(7), A2 => n182, B1 => 
                           zeroSignal(7), B2 => n173, C1 => A_neg_shifted(7), 
                           C2 => n160, ZN => n309);
   U209 : NAND2_X1 port map( A1 => n312, A2 => n311, ZN => Y(8));
   U210 : AOI22_X1 port map( A1 => A_neg(8), A2 => n156, B1 => A_signal(8), B2 
                           => n147, ZN => n312);
   U211 : AOI222_X1 port map( A1 => A_shifted(8), A2 => n182, B1 => 
                           zeroSignal(8), B2 => n173, C1 => A_neg_shifted(8), 
                           C2 => n160, ZN => n311);
   U212 : NAND2_X1 port map( A1 => n318, A2 => n317, ZN => Y(9));
   U213 : AOI22_X1 port map( A1 => A_neg(9), A2 => n156, B1 => A_signal(9), B2 
                           => n147, ZN => n318);
   U214 : AOI222_X1 port map( A1 => A_shifted(9), A2 => n182, B1 => 
                           zeroSignal(9), B2 => n173, C1 => A_neg_shifted(9), 
                           C2 => n160, ZN => n317);
   U215 : NAND2_X1 port map( A1 => n190, A2 => n189, ZN => Y(10));
   U216 : AOI22_X1 port map( A1 => A_neg(10), A2 => n151, B1 => A_signal(10), 
                           B2 => n142, ZN => n190);
   U217 : AOI222_X1 port map( A1 => A_shifted(10), A2 => n177, B1 => 
                           zeroSignal(10), B2 => n168, C1 => A_neg_shifted(10),
                           C2 => n165, ZN => n189);
   U218 : NAND2_X1 port map( A1 => n192, A2 => n191, ZN => Y(11));
   U219 : AOI22_X1 port map( A1 => A_neg(11), A2 => n151, B1 => A_signal(11), 
                           B2 => n142, ZN => n192);
   U220 : AOI222_X1 port map( A1 => A_shifted(11), A2 => n177, B1 => 
                           zeroSignal(11), B2 => n168, C1 => A_neg_shifted(11),
                           C2 => n165, ZN => n191);
   U221 : NAND2_X1 port map( A1 => n194, A2 => n193, ZN => Y(12));
   U222 : AOI22_X1 port map( A1 => A_neg(12), A2 => n151, B1 => A_signal(12), 
                           B2 => n142, ZN => n194);
   U223 : AOI222_X1 port map( A1 => A_shifted(12), A2 => n177, B1 => 
                           zeroSignal(12), B2 => n168, C1 => A_neg_shifted(12),
                           C2 => n165, ZN => n193);
   U224 : NAND2_X1 port map( A1 => n196, A2 => n195, ZN => Y(13));
   U225 : AOI22_X1 port map( A1 => A_neg(13), A2 => n151, B1 => A_signal(13), 
                           B2 => n142, ZN => n196);
   U226 : AOI222_X1 port map( A1 => A_shifted(13), A2 => n177, B1 => 
                           zeroSignal(13), B2 => n168, C1 => A_neg_shifted(13),
                           C2 => n164, ZN => n195);
   U227 : NAND2_X1 port map( A1 => n198, A2 => n197, ZN => Y(14));
   U228 : AOI22_X1 port map( A1 => A_neg(14), A2 => n151, B1 => A_signal(14), 
                           B2 => n142, ZN => n198);
   U229 : AOI222_X1 port map( A1 => A_shifted(14), A2 => n177, B1 => 
                           zeroSignal(14), B2 => n168, C1 => A_neg_shifted(14),
                           C2 => n164, ZN => n197);
   U230 : NAND2_X1 port map( A1 => n200, A2 => n199, ZN => Y(15));
   U231 : AOI22_X1 port map( A1 => A_neg(15), A2 => n151, B1 => A_signal(15), 
                           B2 => n142, ZN => n200);
   U232 : AOI222_X1 port map( A1 => A_shifted(15), A2 => n177, B1 => 
                           zeroSignal(15), B2 => n168, C1 => A_neg_shifted(15),
                           C2 => n164, ZN => n199);
   U233 : NAND2_X1 port map( A1 => n202, A2 => n201, ZN => Y(16));
   U234 : AOI22_X1 port map( A1 => A_neg(16), A2 => n151, B1 => A_signal(16), 
                           B2 => n142, ZN => n202);
   U235 : AOI222_X1 port map( A1 => A_shifted(16), A2 => n177, B1 => 
                           zeroSignal(16), B2 => n168, C1 => A_neg_shifted(16),
                           C2 => n164, ZN => n201);
   U236 : NAND2_X1 port map( A1 => n204, A2 => n203, ZN => Y(17));
   U237 : AOI22_X1 port map( A1 => A_neg(17), A2 => n151, B1 => A_signal(17), 
                           B2 => n142, ZN => n204);
   U238 : AOI222_X1 port map( A1 => A_shifted(17), A2 => n177, B1 => 
                           zeroSignal(17), B2 => n168, C1 => A_neg_shifted(17),
                           C2 => n164, ZN => n203);
   U239 : AOI22_X1 port map( A1 => A_neg(24), A2 => n152, B1 => A_signal(24), 
                           B2 => n143, ZN => n220);
   U240 : AOI22_X1 port map( A1 => A_neg(23), A2 => n152, B1 => A_signal(23), 
                           B2 => n143, ZN => n218);
   U241 : AOI22_X1 port map( A1 => A_neg(21), A2 => n152, B1 => A_signal(21), 
                           B2 => n143, ZN => n214);
   U242 : AOI22_X1 port map( A1 => A_neg(63), A2 => n155, B1 => A_signal(63), 
                           B2 => n146, ZN => n306);
   U243 : AOI222_X1 port map( A1 => A_shifted(61), A2 => n182, B1 => 
                           zeroSignal(61), B2 => n172, C1 => A_neg_shifted(61),
                           C2 => n160, ZN => n301);
   U244 : AOI22_X1 port map( A1 => A_neg(60), A2 => n155, B1 => A_signal(60), 
                           B2 => n146, ZN => n300);

end SYN_BEHAVIORAL_2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity MUX51_MuxNbit64_6 is

   port( zeroSignal, A_signal, A_neg, A_shifted, A_neg_shifted : in 
         std_logic_vector (63 downto 0);  Sel : in std_logic_vector (2 downto 
         0);  Y : out std_logic_vector (63 downto 0));

end MUX51_MuxNbit64_6;

architecture SYN_BEHAVIORAL_2 of MUX51_MuxNbit64_6 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, 
      n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, 
      n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, 
      n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, 
      n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, 
      n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, 
      n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, 
      n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, 
      n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, 
      n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, 
      n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, 
      n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, 
      n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, 
      n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, 
      n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, 
      n320 : std_logic;

begin
   
   U1 : AND3_X1 port map( A1 => n319, A2 => n320, A3 => Sel(2), ZN => n141);
   U2 : BUF_X1 port map( A => n141, Z => n166);
   U3 : BUF_X1 port map( A => n159, Z => n158);
   U4 : BUF_X1 port map( A => n185, Z => n184);
   U5 : BUF_X1 port map( A => n150, Z => n149);
   U6 : BUF_X1 port map( A => n141, Z => n167);
   U7 : BUF_X1 port map( A => n185, Z => n183);
   U8 : BUF_X1 port map( A => n159, Z => n157);
   U9 : BUF_X1 port map( A => n150, Z => n148);
   U10 : BUF_X1 port map( A => n176, Z => n175);
   U11 : BUF_X1 port map( A => n176, Z => n174);
   U12 : BUF_X1 port map( A => n184, Z => n178);
   U13 : BUF_X1 port map( A => n158, Z => n152);
   U14 : BUF_X1 port map( A => n149, Z => n143);
   U15 : BUF_X1 port map( A => n166, Z => n164);
   U16 : BUF_X1 port map( A => n166, Z => n163);
   U17 : BUF_X1 port map( A => n184, Z => n179);
   U18 : BUF_X1 port map( A => n158, Z => n153);
   U19 : BUF_X1 port map( A => n149, Z => n144);
   U20 : BUF_X1 port map( A => n167, Z => n162);
   U21 : BUF_X1 port map( A => n183, Z => n180);
   U22 : BUF_X1 port map( A => n157, Z => n154);
   U23 : BUF_X1 port map( A => n148, Z => n145);
   U24 : BUF_X1 port map( A => n167, Z => n161);
   U25 : BUF_X1 port map( A => n183, Z => n181);
   U26 : BUF_X1 port map( A => n157, Z => n155);
   U27 : BUF_X1 port map( A => n148, Z => n146);
   U28 : BUF_X1 port map( A => n167, Z => n160);
   U29 : BUF_X1 port map( A => n183, Z => n182);
   U30 : BUF_X1 port map( A => n158, Z => n151);
   U31 : BUF_X1 port map( A => n149, Z => n142);
   U32 : BUF_X1 port map( A => n175, Z => n168);
   U33 : BUF_X1 port map( A => n175, Z => n169);
   U34 : BUF_X1 port map( A => n175, Z => n170);
   U35 : BUF_X1 port map( A => n174, Z => n171);
   U36 : BUF_X1 port map( A => n174, Z => n172);
   U37 : BUF_X1 port map( A => n184, Z => n177);
   U38 : BUF_X1 port map( A => n166, Z => n165);
   U39 : BUF_X1 port map( A => n157, Z => n156);
   U40 : BUF_X1 port map( A => n148, Z => n147);
   U41 : BUF_X1 port map( A => n174, Z => n173);
   U42 : INV_X1 port map( A => Sel(1), ZN => n320);
   U43 : BUF_X1 port map( A => n316, Z => n185);
   U44 : NOR3_X1 port map( A1 => n319, A2 => Sel(2), A3 => n320, ZN => n316);
   U45 : BUF_X1 port map( A => n314, Z => n159);
   U46 : NOR3_X1 port map( A1 => Sel(0), A2 => Sel(2), A3 => n320, ZN => n314);
   U47 : INV_X1 port map( A => Sel(0), ZN => n319);
   U48 : BUF_X1 port map( A => n313, Z => n150);
   U49 : NOR3_X1 port map( A1 => Sel(1), A2 => Sel(2), A3 => n319, ZN => n313);
   U50 : BUF_X1 port map( A => n315, Z => n176);
   U51 : NOR2_X1 port map( A1 => n165, A2 => n186, ZN => n315);
   U52 : AOI21_X1 port map( B1 => n319, B2 => n320, A => Sel(2), ZN => n186);
   U53 : NAND2_X1 port map( A1 => n214, A2 => n213, ZN => Y(21));
   U54 : AOI22_X1 port map( A1 => A_neg(21), A2 => n152, B1 => A_signal(21), B2
                           => n143, ZN => n214);
   U55 : AOI222_X1 port map( A1 => A_shifted(21), A2 => n178, B1 => 
                           zeroSignal(21), B2 => n169, C1 => A_neg_shifted(21),
                           C2 => n164, ZN => n213);
   U56 : NAND2_X1 port map( A1 => n212, A2 => n211, ZN => Y(20));
   U57 : AOI222_X1 port map( A1 => A_shifted(20), A2 => n178, B1 => 
                           zeroSignal(20), B2 => n169, C1 => A_neg_shifted(20),
                           C2 => n164, ZN => n211);
   U58 : AOI22_X1 port map( A1 => A_neg(20), A2 => n152, B1 => A_signal(20), B2
                           => n143, ZN => n212);
   U59 : NAND2_X1 port map( A1 => n244, A2 => n243, ZN => Y(35));
   U60 : AOI222_X1 port map( A1 => A_shifted(35), A2 => n179, B1 => 
                           zeroSignal(35), B2 => n170, C1 => A_neg_shifted(35),
                           C2 => n162, ZN => n243);
   U61 : AOI22_X1 port map( A1 => A_neg(35), A2 => n153, B1 => A_signal(35), B2
                           => n144, ZN => n244);
   U62 : NAND2_X1 port map( A1 => n242, A2 => n241, ZN => Y(34));
   U63 : AOI222_X1 port map( A1 => A_shifted(34), A2 => n179, B1 => 
                           zeroSignal(34), B2 => n170, C1 => A_neg_shifted(34),
                           C2 => n163, ZN => n241);
   U64 : AOI22_X1 port map( A1 => A_neg(34), A2 => n153, B1 => A_signal(34), B2
                           => n144, ZN => n242);
   U65 : NAND2_X1 port map( A1 => n240, A2 => n239, ZN => Y(33));
   U66 : AOI222_X1 port map( A1 => A_shifted(33), A2 => n179, B1 => 
                           zeroSignal(33), B2 => n170, C1 => A_neg_shifted(33),
                           C2 => n163, ZN => n239);
   U67 : AOI22_X1 port map( A1 => A_neg(33), A2 => n153, B1 => A_signal(33), B2
                           => n144, ZN => n240);
   U68 : NAND2_X1 port map( A1 => n216, A2 => n215, ZN => Y(22));
   U69 : AOI22_X1 port map( A1 => A_neg(22), A2 => n152, B1 => A_signal(22), B2
                           => n143, ZN => n216);
   U70 : AOI222_X1 port map( A1 => A_shifted(22), A2 => n178, B1 => 
                           zeroSignal(22), B2 => n169, C1 => A_neg_shifted(22),
                           C2 => n164, ZN => n215);
   U71 : NAND2_X1 port map( A1 => n246, A2 => n245, ZN => Y(36));
   U72 : AOI222_X1 port map( A1 => A_shifted(36), A2 => n179, B1 => 
                           zeroSignal(36), B2 => n170, C1 => A_neg_shifted(36),
                           C2 => n162, ZN => n245);
   U73 : AOI22_X1 port map( A1 => A_neg(36), A2 => n153, B1 => A_signal(36), B2
                           => n144, ZN => n246);
   U74 : NAND2_X1 port map( A1 => n248, A2 => n247, ZN => Y(37));
   U75 : AOI222_X1 port map( A1 => A_shifted(37), A2 => n179, B1 => 
                           zeroSignal(37), B2 => n170, C1 => A_neg_shifted(37),
                           C2 => n162, ZN => n247);
   U76 : AOI22_X1 port map( A1 => A_neg(37), A2 => n153, B1 => A_signal(37), B2
                           => n144, ZN => n248);
   U77 : NAND2_X1 port map( A1 => n252, A2 => n251, ZN => Y(39));
   U78 : AOI222_X1 port map( A1 => A_shifted(39), A2 => n179, B1 => 
                           zeroSignal(39), B2 => n170, C1 => A_neg_shifted(39),
                           C2 => n162, ZN => n251);
   U79 : AOI22_X1 port map( A1 => A_neg(39), A2 => n153, B1 => A_signal(39), B2
                           => n144, ZN => n252);
   U80 : NAND2_X1 port map( A1 => n256, A2 => n255, ZN => Y(40));
   U81 : AOI222_X1 port map( A1 => A_shifted(40), A2 => n180, B1 => 
                           zeroSignal(40), B2 => n170, C1 => A_neg_shifted(40),
                           C2 => n162, ZN => n255);
   U82 : AOI22_X1 port map( A1 => A_neg(40), A2 => n153, B1 => A_signal(40), B2
                           => n144, ZN => n256);
   U83 : NAND2_X1 port map( A1 => n258, A2 => n257, ZN => Y(41));
   U84 : AOI222_X1 port map( A1 => A_shifted(41), A2 => n180, B1 => 
                           zeroSignal(41), B2 => n170, C1 => A_neg_shifted(41),
                           C2 => n162, ZN => n257);
   U85 : AOI22_X1 port map( A1 => A_neg(41), A2 => n153, B1 => A_signal(41), B2
                           => n144, ZN => n258);
   U86 : NAND2_X1 port map( A1 => n260, A2 => n259, ZN => Y(42));
   U87 : AOI222_X1 port map( A1 => A_shifted(42), A2 => n180, B1 => 
                           zeroSignal(42), B2 => n171, C1 => A_neg_shifted(42),
                           C2 => n162, ZN => n259);
   U88 : AOI22_X1 port map( A1 => A_neg(42), A2 => n154, B1 => A_signal(42), B2
                           => n145, ZN => n260);
   U89 : NAND2_X1 port map( A1 => n262, A2 => n261, ZN => Y(43));
   U90 : AOI222_X1 port map( A1 => A_shifted(43), A2 => n180, B1 => 
                           zeroSignal(43), B2 => n171, C1 => A_neg_shifted(43),
                           C2 => n162, ZN => n261);
   U91 : AOI22_X1 port map( A1 => A_neg(43), A2 => n154, B1 => A_signal(43), B2
                           => n145, ZN => n262);
   U92 : NAND2_X1 port map( A1 => n264, A2 => n263, ZN => Y(44));
   U93 : AOI222_X1 port map( A1 => A_shifted(44), A2 => n180, B1 => 
                           zeroSignal(44), B2 => n171, C1 => A_neg_shifted(44),
                           C2 => n162, ZN => n263);
   U94 : AOI22_X1 port map( A1 => A_neg(44), A2 => n154, B1 => A_signal(44), B2
                           => n145, ZN => n264);
   U95 : NAND2_X1 port map( A1 => n266, A2 => n265, ZN => Y(45));
   U96 : AOI222_X1 port map( A1 => A_shifted(45), A2 => n180, B1 => 
                           zeroSignal(45), B2 => n171, C1 => A_neg_shifted(45),
                           C2 => n162, ZN => n265);
   U97 : AOI22_X1 port map( A1 => A_neg(45), A2 => n154, B1 => A_signal(45), B2
                           => n145, ZN => n266);
   U98 : NAND2_X1 port map( A1 => n268, A2 => n267, ZN => Y(46));
   U99 : AOI222_X1 port map( A1 => A_shifted(46), A2 => n180, B1 => 
                           zeroSignal(46), B2 => n171, C1 => A_neg_shifted(46),
                           C2 => n161, ZN => n267);
   U100 : AOI22_X1 port map( A1 => A_neg(46), A2 => n154, B1 => A_signal(46), 
                           B2 => n145, ZN => n268);
   U101 : NAND2_X1 port map( A1 => n270, A2 => n269, ZN => Y(47));
   U102 : AOI222_X1 port map( A1 => A_shifted(47), A2 => n180, B1 => 
                           zeroSignal(47), B2 => n171, C1 => A_neg_shifted(47),
                           C2 => n161, ZN => n269);
   U103 : AOI22_X1 port map( A1 => A_neg(47), A2 => n154, B1 => A_signal(47), 
                           B2 => n145, ZN => n270);
   U104 : NAND2_X1 port map( A1 => n272, A2 => n271, ZN => Y(48));
   U105 : AOI222_X1 port map( A1 => A_shifted(48), A2 => n180, B1 => 
                           zeroSignal(48), B2 => n171, C1 => A_neg_shifted(48),
                           C2 => n161, ZN => n271);
   U106 : AOI22_X1 port map( A1 => A_neg(48), A2 => n154, B1 => A_signal(48), 
                           B2 => n145, ZN => n272);
   U107 : NAND2_X1 port map( A1 => n250, A2 => n249, ZN => Y(38));
   U108 : AOI22_X1 port map( A1 => A_neg(38), A2 => n153, B1 => A_signal(38), 
                           B2 => n144, ZN => n250);
   U109 : AOI222_X1 port map( A1 => A_shifted(38), A2 => n179, B1 => 
                           zeroSignal(38), B2 => n170, C1 => A_neg_shifted(38),
                           C2 => n162, ZN => n249);
   U110 : NAND2_X1 port map( A1 => n218, A2 => n217, ZN => Y(23));
   U111 : AOI222_X1 port map( A1 => A_shifted(23), A2 => n178, B1 => 
                           zeroSignal(23), B2 => n169, C1 => A_neg_shifted(23),
                           C2 => n164, ZN => n217);
   U112 : NAND2_X1 port map( A1 => n278, A2 => n277, ZN => Y(50));
   U113 : AOI222_X1 port map( A1 => A_shifted(50), A2 => n181, B1 => 
                           zeroSignal(50), B2 => n171, C1 => A_neg_shifted(50),
                           C2 => n161, ZN => n277);
   U114 : AOI22_X1 port map( A1 => A_neg(50), A2 => n154, B1 => A_signal(50), 
                           B2 => n145, ZN => n278);
   U115 : NAND2_X1 port map( A1 => n280, A2 => n279, ZN => Y(51));
   U116 : AOI222_X1 port map( A1 => A_shifted(51), A2 => n181, B1 => 
                           zeroSignal(51), B2 => n171, C1 => A_neg_shifted(51),
                           C2 => n161, ZN => n279);
   U117 : AOI22_X1 port map( A1 => A_neg(51), A2 => n154, B1 => A_signal(51), 
                           B2 => n145, ZN => n280);
   U118 : NAND2_X1 port map( A1 => n282, A2 => n281, ZN => Y(52));
   U119 : AOI222_X1 port map( A1 => A_shifted(52), A2 => n181, B1 => 
                           zeroSignal(52), B2 => n171, C1 => A_neg_shifted(52),
                           C2 => n161, ZN => n281);
   U120 : AOI22_X1 port map( A1 => A_neg(52), A2 => n154, B1 => A_signal(52), 
                           B2 => n145, ZN => n282);
   U121 : NAND2_X1 port map( A1 => n284, A2 => n283, ZN => Y(53));
   U122 : AOI222_X1 port map( A1 => A_shifted(53), A2 => n181, B1 => 
                           zeroSignal(53), B2 => n172, C1 => A_neg_shifted(53),
                           C2 => n161, ZN => n283);
   U123 : AOI22_X1 port map( A1 => A_neg(53), A2 => n155, B1 => A_signal(53), 
                           B2 => n146, ZN => n284);
   U124 : NAND2_X1 port map( A1 => n274, A2 => n273, ZN => Y(49));
   U125 : AOI22_X1 port map( A1 => A_neg(49), A2 => n154, B1 => A_signal(49), 
                           B2 => n145, ZN => n274);
   U126 : AOI222_X1 port map( A1 => A_shifted(49), A2 => n180, B1 => 
                           zeroSignal(49), B2 => n171, C1 => A_neg_shifted(49),
                           C2 => n161, ZN => n273);
   U127 : NAND2_X1 port map( A1 => n234, A2 => n233, ZN => Y(30));
   U128 : AOI222_X1 port map( A1 => A_shifted(30), A2 => n179, B1 => 
                           zeroSignal(30), B2 => n169, C1 => A_neg_shifted(30),
                           C2 => n163, ZN => n233);
   U129 : AOI22_X1 port map( A1 => A_neg(30), A2 => n152, B1 => A_signal(30), 
                           B2 => n143, ZN => n234);
   U130 : NAND2_X1 port map( A1 => n220, A2 => n219, ZN => Y(24));
   U131 : AOI22_X1 port map( A1 => A_neg(24), A2 => n152, B1 => A_signal(24), 
                           B2 => n143, ZN => n220);
   U132 : AOI222_X1 port map( A1 => A_shifted(24), A2 => n178, B1 => 
                           zeroSignal(24), B2 => n169, C1 => A_neg_shifted(24),
                           C2 => n163, ZN => n219);
   U133 : NAND2_X1 port map( A1 => n238, A2 => n237, ZN => Y(32));
   U134 : AOI222_X1 port map( A1 => A_shifted(32), A2 => n179, B1 => 
                           zeroSignal(32), B2 => n170, C1 => A_neg_shifted(32),
                           C2 => n163, ZN => n237);
   U135 : AOI22_X1 port map( A1 => A_neg(32), A2 => n153, B1 => A_signal(32), 
                           B2 => n144, ZN => n238);
   U136 : NAND2_X1 port map( A1 => n236, A2 => n235, ZN => Y(31));
   U137 : AOI22_X1 port map( A1 => A_neg(31), A2 => n153, B1 => A_signal(31), 
                           B2 => n144, ZN => n236);
   U138 : AOI222_X1 port map( A1 => A_shifted(31), A2 => n179, B1 => 
                           zeroSignal(31), B2 => n170, C1 => A_neg_shifted(31),
                           C2 => n163, ZN => n235);
   U139 : NAND2_X1 port map( A1 => n286, A2 => n285, ZN => Y(54));
   U140 : AOI222_X1 port map( A1 => A_shifted(54), A2 => n181, B1 => 
                           zeroSignal(54), B2 => n172, C1 => A_neg_shifted(54),
                           C2 => n161, ZN => n285);
   U141 : AOI22_X1 port map( A1 => A_neg(54), A2 => n155, B1 => A_signal(54), 
                           B2 => n146, ZN => n286);
   U142 : NAND2_X1 port map( A1 => n288, A2 => n287, ZN => Y(55));
   U143 : AOI222_X1 port map( A1 => A_shifted(55), A2 => n181, B1 => 
                           zeroSignal(55), B2 => n172, C1 => A_neg_shifted(55),
                           C2 => n161, ZN => n287);
   U144 : AOI22_X1 port map( A1 => A_neg(55), A2 => n155, B1 => A_signal(55), 
                           B2 => n146, ZN => n288);
   U145 : NAND2_X1 port map( A1 => n230, A2 => n229, ZN => Y(29));
   U146 : AOI222_X1 port map( A1 => A_shifted(29), A2 => n178, B1 => 
                           zeroSignal(29), B2 => n169, C1 => A_neg_shifted(29),
                           C2 => n163, ZN => n229);
   U147 : AOI22_X1 port map( A1 => A_neg(29), A2 => n152, B1 => A_signal(29), 
                           B2 => n143, ZN => n230);
   U148 : NAND2_X1 port map( A1 => n290, A2 => n289, ZN => Y(56));
   U149 : AOI222_X1 port map( A1 => A_shifted(56), A2 => n181, B1 => 
                           zeroSignal(56), B2 => n172, C1 => A_neg_shifted(56),
                           C2 => n161, ZN => n289);
   U150 : AOI22_X1 port map( A1 => A_neg(56), A2 => n155, B1 => A_signal(56), 
                           B2 => n146, ZN => n290);
   U151 : NAND2_X1 port map( A1 => n226, A2 => n225, ZN => Y(27));
   U152 : AOI222_X1 port map( A1 => A_shifted(27), A2 => n178, B1 => 
                           zeroSignal(27), B2 => n169, C1 => A_neg_shifted(27),
                           C2 => n163, ZN => n225);
   U153 : AOI22_X1 port map( A1 => A_neg(27), A2 => n152, B1 => A_signal(27), 
                           B2 => n143, ZN => n226);
   U154 : NAND2_X1 port map( A1 => n228, A2 => n227, ZN => Y(28));
   U155 : AOI222_X1 port map( A1 => A_shifted(28), A2 => n178, B1 => 
                           zeroSignal(28), B2 => n169, C1 => A_neg_shifted(28),
                           C2 => n163, ZN => n227);
   U156 : AOI22_X1 port map( A1 => A_neg(28), A2 => n152, B1 => A_signal(28), 
                           B2 => n143, ZN => n228);
   U157 : NAND2_X1 port map( A1 => n222, A2 => n221, ZN => Y(25));
   U158 : AOI222_X1 port map( A1 => A_shifted(25), A2 => n178, B1 => 
                           zeroSignal(25), B2 => n169, C1 => A_neg_shifted(25),
                           C2 => n163, ZN => n221);
   U159 : NAND2_X1 port map( A1 => n292, A2 => n291, ZN => Y(57));
   U160 : AOI222_X1 port map( A1 => A_shifted(57), A2 => n181, B1 => 
                           zeroSignal(57), B2 => n172, C1 => A_neg_shifted(57),
                           C2 => n160, ZN => n291);
   U161 : AOI22_X1 port map( A1 => A_neg(57), A2 => n155, B1 => A_signal(57), 
                           B2 => n146, ZN => n292);
   U162 : NAND2_X1 port map( A1 => n224, A2 => n223, ZN => Y(26));
   U163 : AOI222_X1 port map( A1 => A_shifted(26), A2 => n178, B1 => 
                           zeroSignal(26), B2 => n169, C1 => A_neg_shifted(26),
                           C2 => n163, ZN => n223);
   U164 : NAND2_X1 port map( A1 => n294, A2 => n293, ZN => Y(58));
   U165 : AOI22_X1 port map( A1 => A_neg(58), A2 => n155, B1 => A_signal(58), 
                           B2 => n146, ZN => n294);
   U166 : AOI222_X1 port map( A1 => A_shifted(58), A2 => n181, B1 => 
                           zeroSignal(58), B2 => n172, C1 => A_neg_shifted(58),
                           C2 => n160, ZN => n293);
   U167 : NAND2_X1 port map( A1 => n300, A2 => n299, ZN => Y(60));
   U168 : AOI222_X1 port map( A1 => A_shifted(60), A2 => n182, B1 => 
                           zeroSignal(60), B2 => n172, C1 => A_neg_shifted(60),
                           C2 => n160, ZN => n299);
   U169 : AOI22_X1 port map( A1 => A_neg(60), A2 => n155, B1 => A_signal(60), 
                           B2 => n146, ZN => n300);
   U170 : NAND2_X1 port map( A1 => n296, A2 => n295, ZN => Y(59));
   U171 : AOI22_X1 port map( A1 => A_neg(59), A2 => n155, B1 => A_signal(59), 
                           B2 => n146, ZN => n296);
   U172 : AOI222_X1 port map( A1 => A_shifted(59), A2 => n181, B1 => 
                           zeroSignal(59), B2 => n172, C1 => A_neg_shifted(59),
                           C2 => n160, ZN => n295);
   U173 : NAND2_X1 port map( A1 => n302, A2 => n301, ZN => Y(61));
   U174 : AOI22_X1 port map( A1 => A_neg(61), A2 => n155, B1 => A_signal(61), 
                           B2 => n146, ZN => n302);
   U175 : AOI222_X1 port map( A1 => A_shifted(61), A2 => n182, B1 => 
                           zeroSignal(61), B2 => n172, C1 => A_neg_shifted(61),
                           C2 => n160, ZN => n301);
   U176 : NAND2_X1 port map( A1 => n306, A2 => n305, ZN => Y(63));
   U177 : AOI22_X1 port map( A1 => A_neg(63), A2 => n155, B1 => A_signal(63), 
                           B2 => n146, ZN => n306);
   U178 : NAND2_X1 port map( A1 => n304, A2 => n303, ZN => Y(62));
   U179 : AOI222_X1 port map( A1 => A_shifted(62), A2 => n182, B1 => 
                           zeroSignal(62), B2 => n172, C1 => A_neg_shifted(62),
                           C2 => n160, ZN => n303);
   U180 : NAND2_X1 port map( A1 => n188, A2 => n187, ZN => Y(0));
   U181 : AOI22_X1 port map( A1 => A_neg(0), A2 => n151, B1 => A_signal(0), B2 
                           => n142, ZN => n188);
   U182 : AOI222_X1 port map( A1 => A_shifted(0), A2 => n177, B1 => 
                           zeroSignal(0), B2 => n168, C1 => A_neg_shifted(0), 
                           C2 => n165, ZN => n187);
   U183 : NAND2_X1 port map( A1 => n210, A2 => n209, ZN => Y(1));
   U184 : AOI22_X1 port map( A1 => A_neg(1), A2 => n151, B1 => A_signal(1), B2 
                           => n142, ZN => n210);
   U185 : AOI222_X1 port map( A1 => A_shifted(1), A2 => n178, B1 => 
                           zeroSignal(1), B2 => n168, C1 => A_neg_shifted(1), 
                           C2 => n164, ZN => n209);
   U186 : NAND2_X1 port map( A1 => n232, A2 => n231, ZN => Y(2));
   U187 : AOI22_X1 port map( A1 => A_neg(2), A2 => n152, B1 => A_signal(2), B2 
                           => n143, ZN => n232);
   U188 : AOI222_X1 port map( A1 => A_shifted(2), A2 => n179, B1 => 
                           zeroSignal(2), B2 => n169, C1 => A_neg_shifted(2), 
                           C2 => n163, ZN => n231);
   U189 : NAND2_X1 port map( A1 => n254, A2 => n253, ZN => Y(3));
   U190 : AOI22_X1 port map( A1 => A_neg(3), A2 => n153, B1 => A_signal(3), B2 
                           => n144, ZN => n254);
   U191 : AOI222_X1 port map( A1 => A_shifted(3), A2 => n180, B1 => 
                           zeroSignal(3), B2 => n170, C1 => A_neg_shifted(3), 
                           C2 => n162, ZN => n253);
   U192 : NAND2_X1 port map( A1 => n276, A2 => n275, ZN => Y(4));
   U193 : AOI22_X1 port map( A1 => A_neg(4), A2 => n154, B1 => A_signal(4), B2 
                           => n145, ZN => n276);
   U194 : AOI222_X1 port map( A1 => A_shifted(4), A2 => n181, B1 => 
                           zeroSignal(4), B2 => n171, C1 => A_neg_shifted(4), 
                           C2 => n161, ZN => n275);
   U195 : NAND2_X1 port map( A1 => n298, A2 => n297, ZN => Y(5));
   U196 : AOI22_X1 port map( A1 => A_neg(5), A2 => n155, B1 => A_signal(5), B2 
                           => n146, ZN => n298);
   U197 : AOI222_X1 port map( A1 => A_shifted(5), A2 => n182, B1 => 
                           zeroSignal(5), B2 => n172, C1 => A_neg_shifted(5), 
                           C2 => n160, ZN => n297);
   U198 : NAND2_X1 port map( A1 => n308, A2 => n307, ZN => Y(6));
   U199 : AOI22_X1 port map( A1 => A_neg(6), A2 => n156, B1 => A_signal(6), B2 
                           => n147, ZN => n308);
   U200 : AOI222_X1 port map( A1 => A_shifted(6), A2 => n182, B1 => 
                           zeroSignal(6), B2 => n173, C1 => A_neg_shifted(6), 
                           C2 => n160, ZN => n307);
   U201 : NAND2_X1 port map( A1 => n310, A2 => n309, ZN => Y(7));
   U202 : AOI22_X1 port map( A1 => A_neg(7), A2 => n156, B1 => A_signal(7), B2 
                           => n147, ZN => n310);
   U203 : AOI222_X1 port map( A1 => A_shifted(7), A2 => n182, B1 => 
                           zeroSignal(7), B2 => n173, C1 => A_neg_shifted(7), 
                           C2 => n160, ZN => n309);
   U204 : NAND2_X1 port map( A1 => n312, A2 => n311, ZN => Y(8));
   U205 : AOI22_X1 port map( A1 => A_neg(8), A2 => n156, B1 => A_signal(8), B2 
                           => n147, ZN => n312);
   U206 : AOI222_X1 port map( A1 => A_shifted(8), A2 => n182, B1 => 
                           zeroSignal(8), B2 => n173, C1 => A_neg_shifted(8), 
                           C2 => n160, ZN => n311);
   U207 : NAND2_X1 port map( A1 => n318, A2 => n317, ZN => Y(9));
   U208 : AOI22_X1 port map( A1 => A_neg(9), A2 => n156, B1 => A_signal(9), B2 
                           => n147, ZN => n318);
   U209 : AOI222_X1 port map( A1 => A_shifted(9), A2 => n182, B1 => 
                           zeroSignal(9), B2 => n173, C1 => A_neg_shifted(9), 
                           C2 => n160, ZN => n317);
   U210 : NAND2_X1 port map( A1 => n190, A2 => n189, ZN => Y(10));
   U211 : AOI22_X1 port map( A1 => A_neg(10), A2 => n151, B1 => A_signal(10), 
                           B2 => n142, ZN => n190);
   U212 : AOI222_X1 port map( A1 => A_shifted(10), A2 => n177, B1 => 
                           zeroSignal(10), B2 => n168, C1 => A_neg_shifted(10),
                           C2 => n165, ZN => n189);
   U213 : NAND2_X1 port map( A1 => n192, A2 => n191, ZN => Y(11));
   U214 : AOI22_X1 port map( A1 => A_neg(11), A2 => n151, B1 => A_signal(11), 
                           B2 => n142, ZN => n192);
   U215 : AOI222_X1 port map( A1 => A_shifted(11), A2 => n177, B1 => 
                           zeroSignal(11), B2 => n168, C1 => A_neg_shifted(11),
                           C2 => n165, ZN => n191);
   U216 : NAND2_X1 port map( A1 => n194, A2 => n193, ZN => Y(12));
   U217 : AOI22_X1 port map( A1 => A_neg(12), A2 => n151, B1 => A_signal(12), 
                           B2 => n142, ZN => n194);
   U218 : AOI222_X1 port map( A1 => A_shifted(12), A2 => n177, B1 => 
                           zeroSignal(12), B2 => n168, C1 => A_neg_shifted(12),
                           C2 => n165, ZN => n193);
   U219 : NAND2_X1 port map( A1 => n196, A2 => n195, ZN => Y(13));
   U220 : AOI22_X1 port map( A1 => A_neg(13), A2 => n151, B1 => A_signal(13), 
                           B2 => n142, ZN => n196);
   U221 : AOI222_X1 port map( A1 => A_shifted(13), A2 => n177, B1 => 
                           zeroSignal(13), B2 => n168, C1 => A_neg_shifted(13),
                           C2 => n164, ZN => n195);
   U222 : NAND2_X1 port map( A1 => n198, A2 => n197, ZN => Y(14));
   U223 : AOI22_X1 port map( A1 => A_neg(14), A2 => n151, B1 => A_signal(14), 
                           B2 => n142, ZN => n198);
   U224 : AOI222_X1 port map( A1 => A_shifted(14), A2 => n177, B1 => 
                           zeroSignal(14), B2 => n168, C1 => A_neg_shifted(14),
                           C2 => n164, ZN => n197);
   U225 : NAND2_X1 port map( A1 => n200, A2 => n199, ZN => Y(15));
   U226 : AOI22_X1 port map( A1 => A_neg(15), A2 => n151, B1 => A_signal(15), 
                           B2 => n142, ZN => n200);
   U227 : AOI222_X1 port map( A1 => A_shifted(15), A2 => n177, B1 => 
                           zeroSignal(15), B2 => n168, C1 => A_neg_shifted(15),
                           C2 => n164, ZN => n199);
   U228 : NAND2_X1 port map( A1 => n202, A2 => n201, ZN => Y(16));
   U229 : AOI22_X1 port map( A1 => A_neg(16), A2 => n151, B1 => A_signal(16), 
                           B2 => n142, ZN => n202);
   U230 : AOI222_X1 port map( A1 => A_shifted(16), A2 => n177, B1 => 
                           zeroSignal(16), B2 => n168, C1 => A_neg_shifted(16),
                           C2 => n164, ZN => n201);
   U231 : NAND2_X1 port map( A1 => n204, A2 => n203, ZN => Y(17));
   U232 : AOI22_X1 port map( A1 => A_neg(17), A2 => n151, B1 => A_signal(17), 
                           B2 => n142, ZN => n204);
   U233 : AOI222_X1 port map( A1 => A_shifted(17), A2 => n177, B1 => 
                           zeroSignal(17), B2 => n168, C1 => A_neg_shifted(17),
                           C2 => n164, ZN => n203);
   U234 : NAND2_X1 port map( A1 => n206, A2 => n205, ZN => Y(18));
   U235 : AOI22_X1 port map( A1 => A_neg(18), A2 => n151, B1 => A_signal(18), 
                           B2 => n142, ZN => n206);
   U236 : AOI222_X1 port map( A1 => A_shifted(18), A2 => n177, B1 => 
                           zeroSignal(18), B2 => n168, C1 => A_neg_shifted(18),
                           C2 => n164, ZN => n205);
   U237 : NAND2_X1 port map( A1 => n208, A2 => n207, ZN => Y(19));
   U238 : AOI22_X1 port map( A1 => A_neg(19), A2 => n151, B1 => A_signal(19), 
                           B2 => n142, ZN => n208);
   U239 : AOI222_X1 port map( A1 => A_shifted(19), A2 => n177, B1 => 
                           zeroSignal(19), B2 => n168, C1 => A_neg_shifted(19),
                           C2 => n164, ZN => n207);
   U240 : AOI22_X1 port map( A1 => A_neg(26), A2 => n152, B1 => A_signal(26), 
                           B2 => n143, ZN => n224);
   U241 : AOI22_X1 port map( A1 => A_neg(25), A2 => n152, B1 => A_signal(25), 
                           B2 => n143, ZN => n222);
   U242 : AOI22_X1 port map( A1 => A_neg(23), A2 => n152, B1 => A_signal(23), 
                           B2 => n143, ZN => n218);
   U243 : AOI222_X1 port map( A1 => A_shifted(63), A2 => n182, B1 => 
                           zeroSignal(63), B2 => n172, C1 => A_neg_shifted(63),
                           C2 => n160, ZN => n305);
   U244 : AOI22_X1 port map( A1 => A_neg(62), A2 => n155, B1 => A_signal(62), 
                           B2 => n146, ZN => n304);

end SYN_BEHAVIORAL_2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity MUX51_MuxNbit64_5 is

   port( zeroSignal, A_signal, A_neg, A_shifted, A_neg_shifted : in 
         std_logic_vector (63 downto 0);  Sel : in std_logic_vector (2 downto 
         0);  Y : out std_logic_vector (63 downto 0));

end MUX51_MuxNbit64_5;

architecture SYN_BEHAVIORAL_2 of MUX51_MuxNbit64_5 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, 
      n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, 
      n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, 
      n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, 
      n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, 
      n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, 
      n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, 
      n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, 
      n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, 
      n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, 
      n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, 
      n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, 
      n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, 
      n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, 
      n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, 
      n320 : std_logic;

begin
   
   U1 : AND3_X1 port map( A1 => n319, A2 => n320, A3 => Sel(2), ZN => n141);
   U2 : BUF_X1 port map( A => n141, Z => n166);
   U3 : BUF_X1 port map( A => n159, Z => n158);
   U4 : BUF_X1 port map( A => n185, Z => n184);
   U5 : BUF_X1 port map( A => n150, Z => n149);
   U6 : BUF_X1 port map( A => n141, Z => n167);
   U7 : BUF_X1 port map( A => n185, Z => n183);
   U8 : BUF_X1 port map( A => n159, Z => n157);
   U9 : BUF_X1 port map( A => n150, Z => n148);
   U10 : BUF_X1 port map( A => n176, Z => n175);
   U11 : BUF_X1 port map( A => n176, Z => n174);
   U12 : BUF_X1 port map( A => n184, Z => n178);
   U13 : BUF_X1 port map( A => n158, Z => n152);
   U14 : BUF_X1 port map( A => n149, Z => n143);
   U15 : BUF_X1 port map( A => n166, Z => n164);
   U16 : BUF_X1 port map( A => n166, Z => n163);
   U17 : BUF_X1 port map( A => n184, Z => n179);
   U18 : BUF_X1 port map( A => n158, Z => n153);
   U19 : BUF_X1 port map( A => n149, Z => n144);
   U20 : BUF_X1 port map( A => n167, Z => n162);
   U21 : BUF_X1 port map( A => n183, Z => n180);
   U22 : BUF_X1 port map( A => n157, Z => n154);
   U23 : BUF_X1 port map( A => n148, Z => n145);
   U24 : BUF_X1 port map( A => n167, Z => n161);
   U25 : BUF_X1 port map( A => n183, Z => n181);
   U26 : BUF_X1 port map( A => n157, Z => n155);
   U27 : BUF_X1 port map( A => n148, Z => n146);
   U28 : BUF_X1 port map( A => n167, Z => n160);
   U29 : BUF_X1 port map( A => n183, Z => n182);
   U30 : BUF_X1 port map( A => n158, Z => n151);
   U31 : BUF_X1 port map( A => n149, Z => n142);
   U32 : BUF_X1 port map( A => n175, Z => n168);
   U33 : BUF_X1 port map( A => n175, Z => n169);
   U34 : BUF_X1 port map( A => n175, Z => n170);
   U35 : BUF_X1 port map( A => n174, Z => n171);
   U36 : BUF_X1 port map( A => n174, Z => n172);
   U37 : BUF_X1 port map( A => n184, Z => n177);
   U38 : BUF_X1 port map( A => n166, Z => n165);
   U39 : BUF_X1 port map( A => n157, Z => n156);
   U40 : BUF_X1 port map( A => n148, Z => n147);
   U41 : BUF_X1 port map( A => n174, Z => n173);
   U42 : INV_X1 port map( A => Sel(1), ZN => n320);
   U43 : BUF_X1 port map( A => n316, Z => n185);
   U44 : NOR3_X1 port map( A1 => n319, A2 => Sel(2), A3 => n320, ZN => n316);
   U45 : BUF_X1 port map( A => n314, Z => n159);
   U46 : NOR3_X1 port map( A1 => Sel(0), A2 => Sel(2), A3 => n320, ZN => n314);
   U47 : INV_X1 port map( A => Sel(0), ZN => n319);
   U48 : BUF_X1 port map( A => n313, Z => n150);
   U49 : NOR3_X1 port map( A1 => Sel(1), A2 => Sel(2), A3 => n319, ZN => n313);
   U50 : BUF_X1 port map( A => n315, Z => n176);
   U51 : NOR2_X1 port map( A1 => n165, A2 => n186, ZN => n315);
   U52 : AOI21_X1 port map( B1 => n319, B2 => n320, A => Sel(2), ZN => n186);
   U53 : NAND2_X1 port map( A1 => n218, A2 => n217, ZN => Y(23));
   U54 : AOI22_X1 port map( A1 => A_neg(23), A2 => n152, B1 => A_signal(23), B2
                           => n143, ZN => n218);
   U55 : AOI222_X1 port map( A1 => A_shifted(23), A2 => n178, B1 => 
                           zeroSignal(23), B2 => n169, C1 => A_neg_shifted(23),
                           C2 => n164, ZN => n217);
   U56 : NAND2_X1 port map( A1 => n216, A2 => n215, ZN => Y(22));
   U57 : AOI222_X1 port map( A1 => A_shifted(22), A2 => n178, B1 => 
                           zeroSignal(22), B2 => n169, C1 => A_neg_shifted(22),
                           C2 => n164, ZN => n215);
   U58 : AOI22_X1 port map( A1 => A_neg(22), A2 => n152, B1 => A_signal(22), B2
                           => n143, ZN => n216);
   U59 : NAND2_X1 port map( A1 => n248, A2 => n247, ZN => Y(37));
   U60 : AOI222_X1 port map( A1 => A_shifted(37), A2 => n179, B1 => 
                           zeroSignal(37), B2 => n170, C1 => A_neg_shifted(37),
                           C2 => n162, ZN => n247);
   U61 : AOI22_X1 port map( A1 => A_neg(37), A2 => n153, B1 => A_signal(37), B2
                           => n144, ZN => n248);
   U62 : NAND2_X1 port map( A1 => n244, A2 => n243, ZN => Y(35));
   U63 : AOI222_X1 port map( A1 => A_shifted(35), A2 => n179, B1 => 
                           zeroSignal(35), B2 => n170, C1 => A_neg_shifted(35),
                           C2 => n162, ZN => n243);
   U64 : AOI22_X1 port map( A1 => A_neg(35), A2 => n153, B1 => A_signal(35), B2
                           => n144, ZN => n244);
   U65 : NAND2_X1 port map( A1 => n246, A2 => n245, ZN => Y(36));
   U66 : AOI222_X1 port map( A1 => A_shifted(36), A2 => n179, B1 => 
                           zeroSignal(36), B2 => n170, C1 => A_neg_shifted(36),
                           C2 => n162, ZN => n245);
   U67 : AOI22_X1 port map( A1 => A_neg(36), A2 => n153, B1 => A_signal(36), B2
                           => n144, ZN => n246);
   U68 : NAND2_X1 port map( A1 => n220, A2 => n219, ZN => Y(24));
   U69 : AOI22_X1 port map( A1 => A_neg(24), A2 => n152, B1 => A_signal(24), B2
                           => n143, ZN => n220);
   U70 : AOI222_X1 port map( A1 => A_shifted(24), A2 => n178, B1 => 
                           zeroSignal(24), B2 => n169, C1 => A_neg_shifted(24),
                           C2 => n163, ZN => n219);
   U71 : NAND2_X1 port map( A1 => n250, A2 => n249, ZN => Y(38));
   U72 : AOI222_X1 port map( A1 => A_shifted(38), A2 => n179, B1 => 
                           zeroSignal(38), B2 => n170, C1 => A_neg_shifted(38),
                           C2 => n162, ZN => n249);
   U73 : AOI22_X1 port map( A1 => A_neg(38), A2 => n153, B1 => A_signal(38), B2
                           => n144, ZN => n250);
   U74 : NAND2_X1 port map( A1 => n252, A2 => n251, ZN => Y(39));
   U75 : AOI222_X1 port map( A1 => A_shifted(39), A2 => n179, B1 => 
                           zeroSignal(39), B2 => n170, C1 => A_neg_shifted(39),
                           C2 => n162, ZN => n251);
   U76 : AOI22_X1 port map( A1 => A_neg(39), A2 => n153, B1 => A_signal(39), B2
                           => n144, ZN => n252);
   U77 : NAND2_X1 port map( A1 => n258, A2 => n257, ZN => Y(41));
   U78 : AOI222_X1 port map( A1 => A_shifted(41), A2 => n180, B1 => 
                           zeroSignal(41), B2 => n170, C1 => A_neg_shifted(41),
                           C2 => n162, ZN => n257);
   U79 : AOI22_X1 port map( A1 => A_neg(41), A2 => n153, B1 => A_signal(41), B2
                           => n144, ZN => n258);
   U80 : NAND2_X1 port map( A1 => n260, A2 => n259, ZN => Y(42));
   U81 : AOI222_X1 port map( A1 => A_shifted(42), A2 => n180, B1 => 
                           zeroSignal(42), B2 => n171, C1 => A_neg_shifted(42),
                           C2 => n162, ZN => n259);
   U82 : AOI22_X1 port map( A1 => A_neg(42), A2 => n154, B1 => A_signal(42), B2
                           => n145, ZN => n260);
   U83 : NAND2_X1 port map( A1 => n262, A2 => n261, ZN => Y(43));
   U84 : AOI222_X1 port map( A1 => A_shifted(43), A2 => n180, B1 => 
                           zeroSignal(43), B2 => n171, C1 => A_neg_shifted(43),
                           C2 => n162, ZN => n261);
   U85 : AOI22_X1 port map( A1 => A_neg(43), A2 => n154, B1 => A_signal(43), B2
                           => n145, ZN => n262);
   U86 : NAND2_X1 port map( A1 => n264, A2 => n263, ZN => Y(44));
   U87 : AOI222_X1 port map( A1 => A_shifted(44), A2 => n180, B1 => 
                           zeroSignal(44), B2 => n171, C1 => A_neg_shifted(44),
                           C2 => n162, ZN => n263);
   U88 : AOI22_X1 port map( A1 => A_neg(44), A2 => n154, B1 => A_signal(44), B2
                           => n145, ZN => n264);
   U89 : NAND2_X1 port map( A1 => n266, A2 => n265, ZN => Y(45));
   U90 : AOI222_X1 port map( A1 => A_shifted(45), A2 => n180, B1 => 
                           zeroSignal(45), B2 => n171, C1 => A_neg_shifted(45),
                           C2 => n162, ZN => n265);
   U91 : AOI22_X1 port map( A1 => A_neg(45), A2 => n154, B1 => A_signal(45), B2
                           => n145, ZN => n266);
   U92 : NAND2_X1 port map( A1 => n268, A2 => n267, ZN => Y(46));
   U93 : AOI222_X1 port map( A1 => A_shifted(46), A2 => n180, B1 => 
                           zeroSignal(46), B2 => n171, C1 => A_neg_shifted(46),
                           C2 => n161, ZN => n267);
   U94 : AOI22_X1 port map( A1 => A_neg(46), A2 => n154, B1 => A_signal(46), B2
                           => n145, ZN => n268);
   U95 : NAND2_X1 port map( A1 => n270, A2 => n269, ZN => Y(47));
   U96 : AOI222_X1 port map( A1 => A_shifted(47), A2 => n180, B1 => 
                           zeroSignal(47), B2 => n171, C1 => A_neg_shifted(47),
                           C2 => n161, ZN => n269);
   U97 : AOI22_X1 port map( A1 => A_neg(47), A2 => n154, B1 => A_signal(47), B2
                           => n145, ZN => n270);
   U98 : NAND2_X1 port map( A1 => n272, A2 => n271, ZN => Y(48));
   U99 : AOI222_X1 port map( A1 => A_shifted(48), A2 => n180, B1 => 
                           zeroSignal(48), B2 => n171, C1 => A_neg_shifted(48),
                           C2 => n161, ZN => n271);
   U100 : AOI22_X1 port map( A1 => A_neg(48), A2 => n154, B1 => A_signal(48), 
                           B2 => n145, ZN => n272);
   U101 : NAND2_X1 port map( A1 => n274, A2 => n273, ZN => Y(49));
   U102 : AOI222_X1 port map( A1 => A_shifted(49), A2 => n180, B1 => 
                           zeroSignal(49), B2 => n171, C1 => A_neg_shifted(49),
                           C2 => n161, ZN => n273);
   U103 : AOI22_X1 port map( A1 => A_neg(49), A2 => n154, B1 => A_signal(49), 
                           B2 => n145, ZN => n274);
   U104 : NAND2_X1 port map( A1 => n222, A2 => n221, ZN => Y(25));
   U105 : AOI222_X1 port map( A1 => A_shifted(25), A2 => n178, B1 => 
                           zeroSignal(25), B2 => n169, C1 => A_neg_shifted(25),
                           C2 => n163, ZN => n221);
   U106 : NAND2_X1 port map( A1 => n278, A2 => n277, ZN => Y(50));
   U107 : AOI222_X1 port map( A1 => A_shifted(50), A2 => n181, B1 => 
                           zeroSignal(50), B2 => n171, C1 => A_neg_shifted(50),
                           C2 => n161, ZN => n277);
   U108 : AOI22_X1 port map( A1 => A_neg(50), A2 => n154, B1 => A_signal(50), 
                           B2 => n145, ZN => n278);
   U109 : NAND2_X1 port map( A1 => n256, A2 => n255, ZN => Y(40));
   U110 : AOI22_X1 port map( A1 => A_neg(40), A2 => n153, B1 => A_signal(40), 
                           B2 => n144, ZN => n256);
   U111 : AOI222_X1 port map( A1 => A_shifted(40), A2 => n180, B1 => 
                           zeroSignal(40), B2 => n170, C1 => A_neg_shifted(40),
                           C2 => n162, ZN => n255);
   U112 : NAND2_X1 port map( A1 => n282, A2 => n281, ZN => Y(52));
   U113 : AOI222_X1 port map( A1 => A_shifted(52), A2 => n181, B1 => 
                           zeroSignal(52), B2 => n171, C1 => A_neg_shifted(52),
                           C2 => n161, ZN => n281);
   U114 : AOI22_X1 port map( A1 => A_neg(52), A2 => n154, B1 => A_signal(52), 
                           B2 => n145, ZN => n282);
   U115 : NAND2_X1 port map( A1 => n284, A2 => n283, ZN => Y(53));
   U116 : AOI222_X1 port map( A1 => A_shifted(53), A2 => n181, B1 => 
                           zeroSignal(53), B2 => n172, C1 => A_neg_shifted(53),
                           C2 => n161, ZN => n283);
   U117 : AOI22_X1 port map( A1 => A_neg(53), A2 => n155, B1 => A_signal(53), 
                           B2 => n146, ZN => n284);
   U118 : NAND2_X1 port map( A1 => n286, A2 => n285, ZN => Y(54));
   U119 : AOI222_X1 port map( A1 => A_shifted(54), A2 => n181, B1 => 
                           zeroSignal(54), B2 => n172, C1 => A_neg_shifted(54),
                           C2 => n161, ZN => n285);
   U120 : AOI22_X1 port map( A1 => A_neg(54), A2 => n155, B1 => A_signal(54), 
                           B2 => n146, ZN => n286);
   U121 : NAND2_X1 port map( A1 => n288, A2 => n287, ZN => Y(55));
   U122 : AOI222_X1 port map( A1 => A_shifted(55), A2 => n181, B1 => 
                           zeroSignal(55), B2 => n172, C1 => A_neg_shifted(55),
                           C2 => n161, ZN => n287);
   U123 : AOI22_X1 port map( A1 => A_neg(55), A2 => n155, B1 => A_signal(55), 
                           B2 => n146, ZN => n288);
   U124 : NAND2_X1 port map( A1 => n280, A2 => n279, ZN => Y(51));
   U125 : AOI22_X1 port map( A1 => A_neg(51), A2 => n154, B1 => A_signal(51), 
                           B2 => n145, ZN => n280);
   U126 : AOI222_X1 port map( A1 => A_shifted(51), A2 => n181, B1 => 
                           zeroSignal(51), B2 => n171, C1 => A_neg_shifted(51),
                           C2 => n161, ZN => n279);
   U127 : NAND2_X1 port map( A1 => n238, A2 => n237, ZN => Y(32));
   U128 : AOI222_X1 port map( A1 => A_shifted(32), A2 => n179, B1 => 
                           zeroSignal(32), B2 => n170, C1 => A_neg_shifted(32),
                           C2 => n163, ZN => n237);
   U129 : AOI22_X1 port map( A1 => A_neg(32), A2 => n153, B1 => A_signal(32), 
                           B2 => n144, ZN => n238);
   U130 : NAND2_X1 port map( A1 => n242, A2 => n241, ZN => Y(34));
   U131 : AOI222_X1 port map( A1 => A_shifted(34), A2 => n179, B1 => 
                           zeroSignal(34), B2 => n170, C1 => A_neg_shifted(34),
                           C2 => n163, ZN => n241);
   U132 : AOI22_X1 port map( A1 => A_neg(34), A2 => n153, B1 => A_signal(34), 
                           B2 => n144, ZN => n242);
   U133 : NAND2_X1 port map( A1 => n224, A2 => n223, ZN => Y(26));
   U134 : AOI22_X1 port map( A1 => A_neg(26), A2 => n152, B1 => A_signal(26), 
                           B2 => n143, ZN => n224);
   U135 : AOI222_X1 port map( A1 => A_shifted(26), A2 => n178, B1 => 
                           zeroSignal(26), B2 => n169, C1 => A_neg_shifted(26),
                           C2 => n163, ZN => n223);
   U136 : NAND2_X1 port map( A1 => n240, A2 => n239, ZN => Y(33));
   U137 : AOI22_X1 port map( A1 => A_neg(33), A2 => n153, B1 => A_signal(33), 
                           B2 => n144, ZN => n240);
   U138 : AOI222_X1 port map( A1 => A_shifted(33), A2 => n179, B1 => 
                           zeroSignal(33), B2 => n170, C1 => A_neg_shifted(33),
                           C2 => n163, ZN => n239);
   U139 : NAND2_X1 port map( A1 => n290, A2 => n289, ZN => Y(56));
   U140 : AOI222_X1 port map( A1 => A_shifted(56), A2 => n181, B1 => 
                           zeroSignal(56), B2 => n172, C1 => A_neg_shifted(56),
                           C2 => n161, ZN => n289);
   U141 : AOI22_X1 port map( A1 => A_neg(56), A2 => n155, B1 => A_signal(56), 
                           B2 => n146, ZN => n290);
   U142 : NAND2_X1 port map( A1 => n292, A2 => n291, ZN => Y(57));
   U143 : AOI222_X1 port map( A1 => A_shifted(57), A2 => n181, B1 => 
                           zeroSignal(57), B2 => n172, C1 => A_neg_shifted(57),
                           C2 => n160, ZN => n291);
   U144 : AOI22_X1 port map( A1 => A_neg(57), A2 => n155, B1 => A_signal(57), 
                           B2 => n146, ZN => n292);
   U145 : NAND2_X1 port map( A1 => n230, A2 => n229, ZN => Y(29));
   U146 : AOI222_X1 port map( A1 => A_shifted(29), A2 => n178, B1 => 
                           zeroSignal(29), B2 => n169, C1 => A_neg_shifted(29),
                           C2 => n163, ZN => n229);
   U147 : AOI22_X1 port map( A1 => A_neg(29), A2 => n152, B1 => A_signal(29), 
                           B2 => n143, ZN => n230);
   U148 : NAND2_X1 port map( A1 => n234, A2 => n233, ZN => Y(30));
   U149 : AOI222_X1 port map( A1 => A_shifted(30), A2 => n179, B1 => 
                           zeroSignal(30), B2 => n169, C1 => A_neg_shifted(30),
                           C2 => n163, ZN => n233);
   U150 : AOI22_X1 port map( A1 => A_neg(30), A2 => n152, B1 => A_signal(30), 
                           B2 => n143, ZN => n234);
   U151 : NAND2_X1 port map( A1 => n226, A2 => n225, ZN => Y(27));
   U152 : AOI222_X1 port map( A1 => A_shifted(27), A2 => n178, B1 => 
                           zeroSignal(27), B2 => n169, C1 => A_neg_shifted(27),
                           C2 => n163, ZN => n225);
   U153 : NAND2_X1 port map( A1 => n236, A2 => n235, ZN => Y(31));
   U154 : AOI222_X1 port map( A1 => A_shifted(31), A2 => n179, B1 => 
                           zeroSignal(31), B2 => n170, C1 => A_neg_shifted(31),
                           C2 => n163, ZN => n235);
   U155 : AOI22_X1 port map( A1 => A_neg(31), A2 => n153, B1 => A_signal(31), 
                           B2 => n144, ZN => n236);
   U156 : NAND2_X1 port map( A1 => n294, A2 => n293, ZN => Y(58));
   U157 : AOI222_X1 port map( A1 => A_shifted(58), A2 => n181, B1 => 
                           zeroSignal(58), B2 => n172, C1 => A_neg_shifted(58),
                           C2 => n160, ZN => n293);
   U158 : AOI22_X1 port map( A1 => A_neg(58), A2 => n155, B1 => A_signal(58), 
                           B2 => n146, ZN => n294);
   U159 : NAND2_X1 port map( A1 => n296, A2 => n295, ZN => Y(59));
   U160 : AOI222_X1 port map( A1 => A_shifted(59), A2 => n181, B1 => 
                           zeroSignal(59), B2 => n172, C1 => A_neg_shifted(59),
                           C2 => n160, ZN => n295);
   U161 : AOI22_X1 port map( A1 => A_neg(59), A2 => n155, B1 => A_signal(59), 
                           B2 => n146, ZN => n296);
   U162 : NAND2_X1 port map( A1 => n228, A2 => n227, ZN => Y(28));
   U163 : AOI222_X1 port map( A1 => A_shifted(28), A2 => n178, B1 => 
                           zeroSignal(28), B2 => n169, C1 => A_neg_shifted(28),
                           C2 => n163, ZN => n227);
   U164 : NAND2_X1 port map( A1 => n300, A2 => n299, ZN => Y(60));
   U165 : AOI22_X1 port map( A1 => A_neg(60), A2 => n155, B1 => A_signal(60), 
                           B2 => n146, ZN => n300);
   U166 : AOI222_X1 port map( A1 => A_shifted(60), A2 => n182, B1 => 
                           zeroSignal(60), B2 => n172, C1 => A_neg_shifted(60),
                           C2 => n160, ZN => n299);
   U167 : NAND2_X1 port map( A1 => n304, A2 => n303, ZN => Y(62));
   U168 : AOI222_X1 port map( A1 => A_shifted(62), A2 => n182, B1 => 
                           zeroSignal(62), B2 => n172, C1 => A_neg_shifted(62),
                           C2 => n160, ZN => n303);
   U169 : AOI22_X1 port map( A1 => A_neg(62), A2 => n155, B1 => A_signal(62), 
                           B2 => n146, ZN => n304);
   U170 : NAND2_X1 port map( A1 => n302, A2 => n301, ZN => Y(61));
   U171 : AOI22_X1 port map( A1 => A_neg(61), A2 => n155, B1 => A_signal(61), 
                           B2 => n146, ZN => n302);
   U172 : AOI222_X1 port map( A1 => A_shifted(61), A2 => n182, B1 => 
                           zeroSignal(61), B2 => n172, C1 => A_neg_shifted(61),
                           C2 => n160, ZN => n301);
   U173 : NAND2_X1 port map( A1 => n306, A2 => n305, ZN => Y(63));
   U174 : AOI22_X1 port map( A1 => A_neg(63), A2 => n155, B1 => A_signal(63), 
                           B2 => n146, ZN => n306);
   U175 : AOI222_X1 port map( A1 => A_shifted(63), A2 => n182, B1 => 
                           zeroSignal(63), B2 => n172, C1 => A_neg_shifted(63),
                           C2 => n160, ZN => n305);
   U176 : NAND2_X1 port map( A1 => n188, A2 => n187, ZN => Y(0));
   U177 : AOI22_X1 port map( A1 => A_neg(0), A2 => n151, B1 => A_signal(0), B2 
                           => n142, ZN => n188);
   U178 : AOI222_X1 port map( A1 => A_shifted(0), A2 => n177, B1 => 
                           zeroSignal(0), B2 => n168, C1 => A_neg_shifted(0), 
                           C2 => n165, ZN => n187);
   U179 : NAND2_X1 port map( A1 => n210, A2 => n209, ZN => Y(1));
   U180 : AOI22_X1 port map( A1 => A_neg(1), A2 => n151, B1 => A_signal(1), B2 
                           => n142, ZN => n210);
   U181 : AOI222_X1 port map( A1 => A_shifted(1), A2 => n178, B1 => 
                           zeroSignal(1), B2 => n168, C1 => A_neg_shifted(1), 
                           C2 => n164, ZN => n209);
   U182 : NAND2_X1 port map( A1 => n232, A2 => n231, ZN => Y(2));
   U183 : AOI22_X1 port map( A1 => A_neg(2), A2 => n152, B1 => A_signal(2), B2 
                           => n143, ZN => n232);
   U184 : AOI222_X1 port map( A1 => A_shifted(2), A2 => n179, B1 => 
                           zeroSignal(2), B2 => n169, C1 => A_neg_shifted(2), 
                           C2 => n163, ZN => n231);
   U185 : NAND2_X1 port map( A1 => n254, A2 => n253, ZN => Y(3));
   U186 : AOI22_X1 port map( A1 => A_neg(3), A2 => n153, B1 => A_signal(3), B2 
                           => n144, ZN => n254);
   U187 : AOI222_X1 port map( A1 => A_shifted(3), A2 => n180, B1 => 
                           zeroSignal(3), B2 => n170, C1 => A_neg_shifted(3), 
                           C2 => n162, ZN => n253);
   U188 : NAND2_X1 port map( A1 => n276, A2 => n275, ZN => Y(4));
   U189 : AOI22_X1 port map( A1 => A_neg(4), A2 => n154, B1 => A_signal(4), B2 
                           => n145, ZN => n276);
   U190 : AOI222_X1 port map( A1 => A_shifted(4), A2 => n181, B1 => 
                           zeroSignal(4), B2 => n171, C1 => A_neg_shifted(4), 
                           C2 => n161, ZN => n275);
   U191 : NAND2_X1 port map( A1 => n298, A2 => n297, ZN => Y(5));
   U192 : AOI22_X1 port map( A1 => A_neg(5), A2 => n155, B1 => A_signal(5), B2 
                           => n146, ZN => n298);
   U193 : AOI222_X1 port map( A1 => A_shifted(5), A2 => n182, B1 => 
                           zeroSignal(5), B2 => n172, C1 => A_neg_shifted(5), 
                           C2 => n160, ZN => n297);
   U194 : NAND2_X1 port map( A1 => n308, A2 => n307, ZN => Y(6));
   U195 : AOI22_X1 port map( A1 => A_neg(6), A2 => n156, B1 => A_signal(6), B2 
                           => n147, ZN => n308);
   U196 : AOI222_X1 port map( A1 => A_shifted(6), A2 => n182, B1 => 
                           zeroSignal(6), B2 => n173, C1 => A_neg_shifted(6), 
                           C2 => n160, ZN => n307);
   U197 : NAND2_X1 port map( A1 => n310, A2 => n309, ZN => Y(7));
   U198 : AOI22_X1 port map( A1 => A_neg(7), A2 => n156, B1 => A_signal(7), B2 
                           => n147, ZN => n310);
   U199 : AOI222_X1 port map( A1 => A_shifted(7), A2 => n182, B1 => 
                           zeroSignal(7), B2 => n173, C1 => A_neg_shifted(7), 
                           C2 => n160, ZN => n309);
   U200 : NAND2_X1 port map( A1 => n312, A2 => n311, ZN => Y(8));
   U201 : AOI22_X1 port map( A1 => A_neg(8), A2 => n156, B1 => A_signal(8), B2 
                           => n147, ZN => n312);
   U202 : AOI222_X1 port map( A1 => A_shifted(8), A2 => n182, B1 => 
                           zeroSignal(8), B2 => n173, C1 => A_neg_shifted(8), 
                           C2 => n160, ZN => n311);
   U203 : NAND2_X1 port map( A1 => n318, A2 => n317, ZN => Y(9));
   U204 : AOI22_X1 port map( A1 => A_neg(9), A2 => n156, B1 => A_signal(9), B2 
                           => n147, ZN => n318);
   U205 : AOI222_X1 port map( A1 => A_shifted(9), A2 => n182, B1 => 
                           zeroSignal(9), B2 => n173, C1 => A_neg_shifted(9), 
                           C2 => n160, ZN => n317);
   U206 : NAND2_X1 port map( A1 => n190, A2 => n189, ZN => Y(10));
   U207 : AOI22_X1 port map( A1 => A_neg(10), A2 => n151, B1 => A_signal(10), 
                           B2 => n142, ZN => n190);
   U208 : AOI222_X1 port map( A1 => A_shifted(10), A2 => n177, B1 => 
                           zeroSignal(10), B2 => n168, C1 => A_neg_shifted(10),
                           C2 => n165, ZN => n189);
   U209 : NAND2_X1 port map( A1 => n192, A2 => n191, ZN => Y(11));
   U210 : AOI22_X1 port map( A1 => A_neg(11), A2 => n151, B1 => A_signal(11), 
                           B2 => n142, ZN => n192);
   U211 : AOI222_X1 port map( A1 => A_shifted(11), A2 => n177, B1 => 
                           zeroSignal(11), B2 => n168, C1 => A_neg_shifted(11),
                           C2 => n165, ZN => n191);
   U212 : NAND2_X1 port map( A1 => n194, A2 => n193, ZN => Y(12));
   U213 : AOI22_X1 port map( A1 => A_neg(12), A2 => n151, B1 => A_signal(12), 
                           B2 => n142, ZN => n194);
   U214 : AOI222_X1 port map( A1 => A_shifted(12), A2 => n177, B1 => 
                           zeroSignal(12), B2 => n168, C1 => A_neg_shifted(12),
                           C2 => n165, ZN => n193);
   U215 : NAND2_X1 port map( A1 => n196, A2 => n195, ZN => Y(13));
   U216 : AOI22_X1 port map( A1 => A_neg(13), A2 => n151, B1 => A_signal(13), 
                           B2 => n142, ZN => n196);
   U217 : AOI222_X1 port map( A1 => A_shifted(13), A2 => n177, B1 => 
                           zeroSignal(13), B2 => n168, C1 => A_neg_shifted(13),
                           C2 => n164, ZN => n195);
   U218 : NAND2_X1 port map( A1 => n198, A2 => n197, ZN => Y(14));
   U219 : AOI22_X1 port map( A1 => A_neg(14), A2 => n151, B1 => A_signal(14), 
                           B2 => n142, ZN => n198);
   U220 : AOI222_X1 port map( A1 => A_shifted(14), A2 => n177, B1 => 
                           zeroSignal(14), B2 => n168, C1 => A_neg_shifted(14),
                           C2 => n164, ZN => n197);
   U221 : NAND2_X1 port map( A1 => n200, A2 => n199, ZN => Y(15));
   U222 : AOI22_X1 port map( A1 => A_neg(15), A2 => n151, B1 => A_signal(15), 
                           B2 => n142, ZN => n200);
   U223 : AOI222_X1 port map( A1 => A_shifted(15), A2 => n177, B1 => 
                           zeroSignal(15), B2 => n168, C1 => A_neg_shifted(15),
                           C2 => n164, ZN => n199);
   U224 : NAND2_X1 port map( A1 => n202, A2 => n201, ZN => Y(16));
   U225 : AOI22_X1 port map( A1 => A_neg(16), A2 => n151, B1 => A_signal(16), 
                           B2 => n142, ZN => n202);
   U226 : AOI222_X1 port map( A1 => A_shifted(16), A2 => n177, B1 => 
                           zeroSignal(16), B2 => n168, C1 => A_neg_shifted(16),
                           C2 => n164, ZN => n201);
   U227 : NAND2_X1 port map( A1 => n204, A2 => n203, ZN => Y(17));
   U228 : AOI22_X1 port map( A1 => A_neg(17), A2 => n151, B1 => A_signal(17), 
                           B2 => n142, ZN => n204);
   U229 : AOI222_X1 port map( A1 => A_shifted(17), A2 => n177, B1 => 
                           zeroSignal(17), B2 => n168, C1 => A_neg_shifted(17),
                           C2 => n164, ZN => n203);
   U230 : NAND2_X1 port map( A1 => n206, A2 => n205, ZN => Y(18));
   U231 : AOI22_X1 port map( A1 => A_neg(18), A2 => n151, B1 => A_signal(18), 
                           B2 => n142, ZN => n206);
   U232 : AOI222_X1 port map( A1 => A_shifted(18), A2 => n177, B1 => 
                           zeroSignal(18), B2 => n168, C1 => A_neg_shifted(18),
                           C2 => n164, ZN => n205);
   U233 : NAND2_X1 port map( A1 => n208, A2 => n207, ZN => Y(19));
   U234 : AOI22_X1 port map( A1 => A_neg(19), A2 => n151, B1 => A_signal(19), 
                           B2 => n142, ZN => n208);
   U235 : AOI222_X1 port map( A1 => A_shifted(19), A2 => n177, B1 => 
                           zeroSignal(19), B2 => n168, C1 => A_neg_shifted(19),
                           C2 => n164, ZN => n207);
   U236 : NAND2_X1 port map( A1 => n212, A2 => n211, ZN => Y(20));
   U237 : AOI22_X1 port map( A1 => A_neg(20), A2 => n152, B1 => A_signal(20), 
                           B2 => n143, ZN => n212);
   U238 : AOI222_X1 port map( A1 => A_shifted(20), A2 => n178, B1 => 
                           zeroSignal(20), B2 => n169, C1 => A_neg_shifted(20),
                           C2 => n164, ZN => n211);
   U239 : NAND2_X1 port map( A1 => n214, A2 => n213, ZN => Y(21));
   U240 : AOI22_X1 port map( A1 => A_neg(21), A2 => n152, B1 => A_signal(21), 
                           B2 => n143, ZN => n214);
   U241 : AOI222_X1 port map( A1 => A_shifted(21), A2 => n178, B1 => 
                           zeroSignal(21), B2 => n169, C1 => A_neg_shifted(21),
                           C2 => n164, ZN => n213);
   U242 : AOI22_X1 port map( A1 => A_neg(28), A2 => n152, B1 => A_signal(28), 
                           B2 => n143, ZN => n228);
   U243 : AOI22_X1 port map( A1 => A_neg(27), A2 => n152, B1 => A_signal(27), 
                           B2 => n143, ZN => n226);
   U244 : AOI22_X1 port map( A1 => A_neg(25), A2 => n152, B1 => A_signal(25), 
                           B2 => n143, ZN => n222);

end SYN_BEHAVIORAL_2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity MUX51_MuxNbit64_4 is

   port( zeroSignal, A_signal, A_neg, A_shifted, A_neg_shifted : in 
         std_logic_vector (63 downto 0);  Sel : in std_logic_vector (2 downto 
         0);  Y : out std_logic_vector (63 downto 0));

end MUX51_MuxNbit64_4;

architecture SYN_BEHAVIORAL_2 of MUX51_MuxNbit64_4 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, 
      n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, 
      n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, 
      n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, 
      n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, 
      n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, 
      n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, 
      n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, 
      n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, 
      n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, 
      n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, 
      n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, 
      n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, 
      n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, 
      n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, 
      n320 : std_logic;

begin
   
   U1 : AND3_X1 port map( A1 => n319, A2 => n320, A3 => Sel(2), ZN => n141);
   U2 : BUF_X1 port map( A => n141, Z => n166);
   U3 : BUF_X1 port map( A => n159, Z => n158);
   U4 : BUF_X1 port map( A => n185, Z => n184);
   U5 : BUF_X1 port map( A => n150, Z => n149);
   U6 : BUF_X1 port map( A => n141, Z => n167);
   U7 : BUF_X1 port map( A => n185, Z => n183);
   U8 : BUF_X1 port map( A => n159, Z => n157);
   U9 : BUF_X1 port map( A => n150, Z => n148);
   U10 : BUF_X1 port map( A => n176, Z => n175);
   U11 : BUF_X1 port map( A => n176, Z => n174);
   U12 : BUF_X1 port map( A => n184, Z => n178);
   U13 : BUF_X1 port map( A => n158, Z => n152);
   U14 : BUF_X1 port map( A => n149, Z => n143);
   U15 : BUF_X1 port map( A => n166, Z => n163);
   U16 : BUF_X1 port map( A => n184, Z => n179);
   U17 : BUF_X1 port map( A => n158, Z => n153);
   U18 : BUF_X1 port map( A => n149, Z => n144);
   U19 : BUF_X1 port map( A => n167, Z => n162);
   U20 : BUF_X1 port map( A => n183, Z => n180);
   U21 : BUF_X1 port map( A => n157, Z => n154);
   U22 : BUF_X1 port map( A => n148, Z => n145);
   U23 : BUF_X1 port map( A => n167, Z => n161);
   U24 : BUF_X1 port map( A => n183, Z => n181);
   U25 : BUF_X1 port map( A => n157, Z => n155);
   U26 : BUF_X1 port map( A => n148, Z => n146);
   U27 : BUF_X1 port map( A => n167, Z => n160);
   U28 : BUF_X1 port map( A => n183, Z => n182);
   U29 : BUF_X1 port map( A => n158, Z => n151);
   U30 : BUF_X1 port map( A => n149, Z => n142);
   U31 : BUF_X1 port map( A => n175, Z => n168);
   U32 : BUF_X1 port map( A => n175, Z => n169);
   U33 : BUF_X1 port map( A => n175, Z => n170);
   U34 : BUF_X1 port map( A => n174, Z => n171);
   U35 : BUF_X1 port map( A => n174, Z => n172);
   U36 : BUF_X1 port map( A => n166, Z => n164);
   U37 : BUF_X1 port map( A => n184, Z => n177);
   U38 : BUF_X1 port map( A => n166, Z => n165);
   U39 : BUF_X1 port map( A => n157, Z => n156);
   U40 : BUF_X1 port map( A => n148, Z => n147);
   U41 : BUF_X1 port map( A => n174, Z => n173);
   U42 : INV_X1 port map( A => Sel(1), ZN => n320);
   U43 : BUF_X1 port map( A => n316, Z => n185);
   U44 : NOR3_X1 port map( A1 => n319, A2 => Sel(2), A3 => n320, ZN => n316);
   U45 : BUF_X1 port map( A => n314, Z => n159);
   U46 : NOR3_X1 port map( A1 => Sel(0), A2 => Sel(2), A3 => n320, ZN => n314);
   U47 : INV_X1 port map( A => Sel(0), ZN => n319);
   U48 : BUF_X1 port map( A => n313, Z => n150);
   U49 : NOR3_X1 port map( A1 => Sel(1), A2 => Sel(2), A3 => n319, ZN => n313);
   U50 : BUF_X1 port map( A => n315, Z => n176);
   U51 : NOR2_X1 port map( A1 => n165, A2 => n186, ZN => n315);
   U52 : AOI21_X1 port map( B1 => n319, B2 => n320, A => Sel(2), ZN => n186);
   U53 : NAND2_X1 port map( A1 => n222, A2 => n221, ZN => Y(25));
   U54 : AOI22_X1 port map( A1 => A_neg(25), A2 => n152, B1 => A_signal(25), B2
                           => n143, ZN => n222);
   U55 : AOI222_X1 port map( A1 => A_shifted(25), A2 => n178, B1 => 
                           zeroSignal(25), B2 => n169, C1 => A_neg_shifted(25),
                           C2 => n163, ZN => n221);
   U56 : NAND2_X1 port map( A1 => n220, A2 => n219, ZN => Y(24));
   U57 : AOI222_X1 port map( A1 => A_shifted(24), A2 => n178, B1 => 
                           zeroSignal(24), B2 => n169, C1 => A_neg_shifted(24),
                           C2 => n163, ZN => n219);
   U58 : AOI22_X1 port map( A1 => A_neg(24), A2 => n152, B1 => A_signal(24), B2
                           => n143, ZN => n220);
   U59 : NAND2_X1 port map( A1 => n252, A2 => n251, ZN => Y(39));
   U60 : AOI222_X1 port map( A1 => A_shifted(39), A2 => n179, B1 => 
                           zeroSignal(39), B2 => n170, C1 => A_neg_shifted(39),
                           C2 => n162, ZN => n251);
   U61 : AOI22_X1 port map( A1 => A_neg(39), A2 => n153, B1 => A_signal(39), B2
                           => n144, ZN => n252);
   U62 : NAND2_X1 port map( A1 => n248, A2 => n247, ZN => Y(37));
   U63 : AOI222_X1 port map( A1 => A_shifted(37), A2 => n179, B1 => 
                           zeroSignal(37), B2 => n170, C1 => A_neg_shifted(37),
                           C2 => n162, ZN => n247);
   U64 : AOI22_X1 port map( A1 => A_neg(37), A2 => n153, B1 => A_signal(37), B2
                           => n144, ZN => n248);
   U65 : NAND2_X1 port map( A1 => n224, A2 => n223, ZN => Y(26));
   U66 : AOI22_X1 port map( A1 => A_neg(26), A2 => n152, B1 => A_signal(26), B2
                           => n143, ZN => n224);
   U67 : AOI222_X1 port map( A1 => A_shifted(26), A2 => n178, B1 => 
                           zeroSignal(26), B2 => n169, C1 => A_neg_shifted(26),
                           C2 => n163, ZN => n223);
   U68 : NAND2_X1 port map( A1 => n250, A2 => n249, ZN => Y(38));
   U69 : AOI222_X1 port map( A1 => A_shifted(38), A2 => n179, B1 => 
                           zeroSignal(38), B2 => n170, C1 => A_neg_shifted(38),
                           C2 => n162, ZN => n249);
   U70 : AOI22_X1 port map( A1 => A_neg(38), A2 => n153, B1 => A_signal(38), B2
                           => n144, ZN => n250);
   U71 : NAND2_X1 port map( A1 => n256, A2 => n255, ZN => Y(40));
   U72 : AOI222_X1 port map( A1 => A_shifted(40), A2 => n180, B1 => 
                           zeroSignal(40), B2 => n170, C1 => A_neg_shifted(40),
                           C2 => n162, ZN => n255);
   U73 : AOI22_X1 port map( A1 => A_neg(40), A2 => n153, B1 => A_signal(40), B2
                           => n144, ZN => n256);
   U74 : NAND2_X1 port map( A1 => n258, A2 => n257, ZN => Y(41));
   U75 : AOI222_X1 port map( A1 => A_shifted(41), A2 => n180, B1 => 
                           zeroSignal(41), B2 => n170, C1 => A_neg_shifted(41),
                           C2 => n162, ZN => n257);
   U76 : AOI22_X1 port map( A1 => A_neg(41), A2 => n153, B1 => A_signal(41), B2
                           => n144, ZN => n258);
   U77 : NAND2_X1 port map( A1 => n262, A2 => n261, ZN => Y(43));
   U78 : AOI222_X1 port map( A1 => A_shifted(43), A2 => n180, B1 => 
                           zeroSignal(43), B2 => n171, C1 => A_neg_shifted(43),
                           C2 => n162, ZN => n261);
   U79 : AOI22_X1 port map( A1 => A_neg(43), A2 => n154, B1 => A_signal(43), B2
                           => n145, ZN => n262);
   U80 : NAND2_X1 port map( A1 => n264, A2 => n263, ZN => Y(44));
   U81 : AOI222_X1 port map( A1 => A_shifted(44), A2 => n180, B1 => 
                           zeroSignal(44), B2 => n171, C1 => A_neg_shifted(44),
                           C2 => n162, ZN => n263);
   U82 : AOI22_X1 port map( A1 => A_neg(44), A2 => n154, B1 => A_signal(44), B2
                           => n145, ZN => n264);
   U83 : NAND2_X1 port map( A1 => n266, A2 => n265, ZN => Y(45));
   U84 : AOI222_X1 port map( A1 => A_shifted(45), A2 => n180, B1 => 
                           zeroSignal(45), B2 => n171, C1 => A_neg_shifted(45),
                           C2 => n162, ZN => n265);
   U85 : AOI22_X1 port map( A1 => A_neg(45), A2 => n154, B1 => A_signal(45), B2
                           => n145, ZN => n266);
   U86 : NAND2_X1 port map( A1 => n268, A2 => n267, ZN => Y(46));
   U87 : AOI222_X1 port map( A1 => A_shifted(46), A2 => n180, B1 => 
                           zeroSignal(46), B2 => n171, C1 => A_neg_shifted(46),
                           C2 => n161, ZN => n267);
   U88 : AOI22_X1 port map( A1 => A_neg(46), A2 => n154, B1 => A_signal(46), B2
                           => n145, ZN => n268);
   U89 : NAND2_X1 port map( A1 => n270, A2 => n269, ZN => Y(47));
   U90 : AOI222_X1 port map( A1 => A_shifted(47), A2 => n180, B1 => 
                           zeroSignal(47), B2 => n171, C1 => A_neg_shifted(47),
                           C2 => n161, ZN => n269);
   U91 : AOI22_X1 port map( A1 => A_neg(47), A2 => n154, B1 => A_signal(47), B2
                           => n145, ZN => n270);
   U92 : NAND2_X1 port map( A1 => n272, A2 => n271, ZN => Y(48));
   U93 : AOI222_X1 port map( A1 => A_shifted(48), A2 => n180, B1 => 
                           zeroSignal(48), B2 => n171, C1 => A_neg_shifted(48),
                           C2 => n161, ZN => n271);
   U94 : AOI22_X1 port map( A1 => A_neg(48), A2 => n154, B1 => A_signal(48), B2
                           => n145, ZN => n272);
   U95 : NAND2_X1 port map( A1 => n274, A2 => n273, ZN => Y(49));
   U96 : AOI222_X1 port map( A1 => A_shifted(49), A2 => n180, B1 => 
                           zeroSignal(49), B2 => n171, C1 => A_neg_shifted(49),
                           C2 => n161, ZN => n273);
   U97 : AOI22_X1 port map( A1 => A_neg(49), A2 => n154, B1 => A_signal(49), B2
                           => n145, ZN => n274);
   U98 : NAND2_X1 port map( A1 => n278, A2 => n277, ZN => Y(50));
   U99 : AOI222_X1 port map( A1 => A_shifted(50), A2 => n181, B1 => 
                           zeroSignal(50), B2 => n171, C1 => A_neg_shifted(50),
                           C2 => n161, ZN => n277);
   U100 : AOI22_X1 port map( A1 => A_neg(50), A2 => n154, B1 => A_signal(50), 
                           B2 => n145, ZN => n278);
   U101 : NAND2_X1 port map( A1 => n226, A2 => n225, ZN => Y(27));
   U102 : AOI222_X1 port map( A1 => A_shifted(27), A2 => n178, B1 => 
                           zeroSignal(27), B2 => n169, C1 => A_neg_shifted(27),
                           C2 => n163, ZN => n225);
   U103 : NAND2_X1 port map( A1 => n280, A2 => n279, ZN => Y(51));
   U104 : AOI222_X1 port map( A1 => A_shifted(51), A2 => n181, B1 => 
                           zeroSignal(51), B2 => n171, C1 => A_neg_shifted(51),
                           C2 => n161, ZN => n279);
   U105 : AOI22_X1 port map( A1 => A_neg(51), A2 => n154, B1 => A_signal(51), 
                           B2 => n145, ZN => n280);
   U106 : NAND2_X1 port map( A1 => n282, A2 => n281, ZN => Y(52));
   U107 : AOI222_X1 port map( A1 => A_shifted(52), A2 => n181, B1 => 
                           zeroSignal(52), B2 => n171, C1 => A_neg_shifted(52),
                           C2 => n161, ZN => n281);
   U108 : AOI22_X1 port map( A1 => A_neg(52), A2 => n154, B1 => A_signal(52), 
                           B2 => n145, ZN => n282);
   U109 : NAND2_X1 port map( A1 => n260, A2 => n259, ZN => Y(42));
   U110 : AOI22_X1 port map( A1 => A_neg(42), A2 => n154, B1 => A_signal(42), 
                           B2 => n145, ZN => n260);
   U111 : AOI222_X1 port map( A1 => A_shifted(42), A2 => n180, B1 => 
                           zeroSignal(42), B2 => n171, C1 => A_neg_shifted(42),
                           C2 => n162, ZN => n259);
   U112 : NAND2_X1 port map( A1 => n286, A2 => n285, ZN => Y(54));
   U113 : AOI222_X1 port map( A1 => A_shifted(54), A2 => n181, B1 => 
                           zeroSignal(54), B2 => n172, C1 => A_neg_shifted(54),
                           C2 => n161, ZN => n285);
   U114 : AOI22_X1 port map( A1 => A_neg(54), A2 => n155, B1 => A_signal(54), 
                           B2 => n146, ZN => n286);
   U115 : NAND2_X1 port map( A1 => n288, A2 => n287, ZN => Y(55));
   U116 : AOI222_X1 port map( A1 => A_shifted(55), A2 => n181, B1 => 
                           zeroSignal(55), B2 => n172, C1 => A_neg_shifted(55),
                           C2 => n161, ZN => n287);
   U117 : AOI22_X1 port map( A1 => A_neg(55), A2 => n155, B1 => A_signal(55), 
                           B2 => n146, ZN => n288);
   U118 : NAND2_X1 port map( A1 => n290, A2 => n289, ZN => Y(56));
   U119 : AOI222_X1 port map( A1 => A_shifted(56), A2 => n181, B1 => 
                           zeroSignal(56), B2 => n172, C1 => A_neg_shifted(56),
                           C2 => n161, ZN => n289);
   U120 : AOI22_X1 port map( A1 => A_neg(56), A2 => n155, B1 => A_signal(56), 
                           B2 => n146, ZN => n290);
   U121 : NAND2_X1 port map( A1 => n242, A2 => n241, ZN => Y(34));
   U122 : AOI222_X1 port map( A1 => A_shifted(34), A2 => n179, B1 => 
                           zeroSignal(34), B2 => n170, C1 => A_neg_shifted(34),
                           C2 => n163, ZN => n241);
   U123 : AOI22_X1 port map( A1 => A_neg(34), A2 => n153, B1 => A_signal(34), 
                           B2 => n144, ZN => n242);
   U124 : NAND2_X1 port map( A1 => n292, A2 => n291, ZN => Y(57));
   U125 : AOI222_X1 port map( A1 => A_shifted(57), A2 => n181, B1 => 
                           zeroSignal(57), B2 => n172, C1 => A_neg_shifted(57),
                           C2 => n160, ZN => n291);
   U126 : AOI22_X1 port map( A1 => A_neg(57), A2 => n155, B1 => A_signal(57), 
                           B2 => n146, ZN => n292);
   U127 : NAND2_X1 port map( A1 => n284, A2 => n283, ZN => Y(53));
   U128 : AOI22_X1 port map( A1 => A_neg(53), A2 => n155, B1 => A_signal(53), 
                           B2 => n146, ZN => n284);
   U129 : AOI222_X1 port map( A1 => A_shifted(53), A2 => n181, B1 => 
                           zeroSignal(53), B2 => n172, C1 => A_neg_shifted(53),
                           C2 => n161, ZN => n283);
   U130 : NAND2_X1 port map( A1 => n228, A2 => n227, ZN => Y(28));
   U131 : AOI22_X1 port map( A1 => A_neg(28), A2 => n152, B1 => A_signal(28), 
                           B2 => n143, ZN => n228);
   U132 : AOI222_X1 port map( A1 => A_shifted(28), A2 => n178, B1 => 
                           zeroSignal(28), B2 => n169, C1 => A_neg_shifted(28),
                           C2 => n163, ZN => n227);
   U133 : NAND2_X1 port map( A1 => n246, A2 => n245, ZN => Y(36));
   U134 : AOI222_X1 port map( A1 => A_shifted(36), A2 => n179, B1 => 
                           zeroSignal(36), B2 => n170, C1 => A_neg_shifted(36),
                           C2 => n162, ZN => n245);
   U135 : AOI22_X1 port map( A1 => A_neg(36), A2 => n153, B1 => A_signal(36), 
                           B2 => n144, ZN => n246);
   U136 : NAND2_X1 port map( A1 => n244, A2 => n243, ZN => Y(35));
   U137 : AOI22_X1 port map( A1 => A_neg(35), A2 => n153, B1 => A_signal(35), 
                           B2 => n144, ZN => n244);
   U138 : AOI222_X1 port map( A1 => A_shifted(35), A2 => n179, B1 => 
                           zeroSignal(35), B2 => n170, C1 => A_neg_shifted(35),
                           C2 => n162, ZN => n243);
   U139 : NAND2_X1 port map( A1 => n294, A2 => n293, ZN => Y(58));
   U140 : AOI222_X1 port map( A1 => A_shifted(58), A2 => n181, B1 => 
                           zeroSignal(58), B2 => n172, C1 => A_neg_shifted(58),
                           C2 => n160, ZN => n293);
   U141 : AOI22_X1 port map( A1 => A_neg(58), A2 => n155, B1 => A_signal(58), 
                           B2 => n146, ZN => n294);
   U142 : NAND2_X1 port map( A1 => n296, A2 => n295, ZN => Y(59));
   U143 : AOI222_X1 port map( A1 => A_shifted(59), A2 => n181, B1 => 
                           zeroSignal(59), B2 => n172, C1 => A_neg_shifted(59),
                           C2 => n160, ZN => n295);
   U144 : AOI22_X1 port map( A1 => A_neg(59), A2 => n155, B1 => A_signal(59), 
                           B2 => n146, ZN => n296);
   U145 : NAND2_X1 port map( A1 => n230, A2 => n229, ZN => Y(29));
   U146 : AOI222_X1 port map( A1 => A_shifted(29), A2 => n178, B1 => 
                           zeroSignal(29), B2 => n169, C1 => A_neg_shifted(29),
                           C2 => n163, ZN => n229);
   U147 : NAND2_X1 port map( A1 => n236, A2 => n235, ZN => Y(31));
   U148 : AOI222_X1 port map( A1 => A_shifted(31), A2 => n179, B1 => 
                           zeroSignal(31), B2 => n170, C1 => A_neg_shifted(31),
                           C2 => n163, ZN => n235);
   U149 : AOI22_X1 port map( A1 => A_neg(31), A2 => n153, B1 => A_signal(31), 
                           B2 => n144, ZN => n236);
   U150 : NAND2_X1 port map( A1 => n238, A2 => n237, ZN => Y(32));
   U151 : AOI222_X1 port map( A1 => A_shifted(32), A2 => n179, B1 => 
                           zeroSignal(32), B2 => n170, C1 => A_neg_shifted(32),
                           C2 => n163, ZN => n237);
   U152 : AOI22_X1 port map( A1 => A_neg(32), A2 => n153, B1 => A_signal(32), 
                           B2 => n144, ZN => n238);
   U153 : NAND2_X1 port map( A1 => n240, A2 => n239, ZN => Y(33));
   U154 : AOI222_X1 port map( A1 => A_shifted(33), A2 => n179, B1 => 
                           zeroSignal(33), B2 => n170, C1 => A_neg_shifted(33),
                           C2 => n163, ZN => n239);
   U155 : AOI22_X1 port map( A1 => A_neg(33), A2 => n153, B1 => A_signal(33), 
                           B2 => n144, ZN => n240);
   U156 : NAND2_X1 port map( A1 => n300, A2 => n299, ZN => Y(60));
   U157 : AOI222_X1 port map( A1 => A_shifted(60), A2 => n182, B1 => 
                           zeroSignal(60), B2 => n172, C1 => A_neg_shifted(60),
                           C2 => n160, ZN => n299);
   U158 : AOI22_X1 port map( A1 => A_neg(60), A2 => n155, B1 => A_signal(60), 
                           B2 => n146, ZN => n300);
   U159 : NAND2_X1 port map( A1 => n302, A2 => n301, ZN => Y(61));
   U160 : AOI222_X1 port map( A1 => A_shifted(61), A2 => n182, B1 => 
                           zeroSignal(61), B2 => n172, C1 => A_neg_shifted(61),
                           C2 => n160, ZN => n301);
   U161 : AOI22_X1 port map( A1 => A_neg(61), A2 => n155, B1 => A_signal(61), 
                           B2 => n146, ZN => n302);
   U162 : NAND2_X1 port map( A1 => n234, A2 => n233, ZN => Y(30));
   U163 : AOI222_X1 port map( A1 => A_shifted(30), A2 => n179, B1 => 
                           zeroSignal(30), B2 => n169, C1 => A_neg_shifted(30),
                           C2 => n163, ZN => n233);
   U164 : NAND2_X1 port map( A1 => n304, A2 => n303, ZN => Y(62));
   U165 : AOI22_X1 port map( A1 => A_neg(62), A2 => n155, B1 => A_signal(62), 
                           B2 => n146, ZN => n304);
   U166 : AOI222_X1 port map( A1 => A_shifted(62), A2 => n182, B1 => 
                           zeroSignal(62), B2 => n172, C1 => A_neg_shifted(62),
                           C2 => n160, ZN => n303);
   U167 : NAND2_X1 port map( A1 => n306, A2 => n305, ZN => Y(63));
   U168 : AOI22_X1 port map( A1 => A_neg(63), A2 => n155, B1 => A_signal(63), 
                           B2 => n146, ZN => n306);
   U169 : AOI222_X1 port map( A1 => A_shifted(63), A2 => n182, B1 => 
                           zeroSignal(63), B2 => n172, C1 => A_neg_shifted(63),
                           C2 => n160, ZN => n305);
   U170 : NAND2_X1 port map( A1 => n188, A2 => n187, ZN => Y(0));
   U171 : AOI22_X1 port map( A1 => A_neg(0), A2 => n151, B1 => A_signal(0), B2 
                           => n142, ZN => n188);
   U172 : AOI222_X1 port map( A1 => A_shifted(0), A2 => n177, B1 => 
                           zeroSignal(0), B2 => n168, C1 => A_neg_shifted(0), 
                           C2 => n165, ZN => n187);
   U173 : NAND2_X1 port map( A1 => n210, A2 => n209, ZN => Y(1));
   U174 : AOI22_X1 port map( A1 => A_neg(1), A2 => n151, B1 => A_signal(1), B2 
                           => n142, ZN => n210);
   U175 : AOI222_X1 port map( A1 => A_shifted(1), A2 => n178, B1 => 
                           zeroSignal(1), B2 => n168, C1 => A_neg_shifted(1), 
                           C2 => n164, ZN => n209);
   U176 : NAND2_X1 port map( A1 => n232, A2 => n231, ZN => Y(2));
   U177 : AOI22_X1 port map( A1 => A_neg(2), A2 => n152, B1 => A_signal(2), B2 
                           => n143, ZN => n232);
   U178 : AOI222_X1 port map( A1 => A_shifted(2), A2 => n179, B1 => 
                           zeroSignal(2), B2 => n169, C1 => A_neg_shifted(2), 
                           C2 => n163, ZN => n231);
   U179 : NAND2_X1 port map( A1 => n254, A2 => n253, ZN => Y(3));
   U180 : AOI22_X1 port map( A1 => A_neg(3), A2 => n153, B1 => A_signal(3), B2 
                           => n144, ZN => n254);
   U181 : AOI222_X1 port map( A1 => A_shifted(3), A2 => n180, B1 => 
                           zeroSignal(3), B2 => n170, C1 => A_neg_shifted(3), 
                           C2 => n162, ZN => n253);
   U182 : NAND2_X1 port map( A1 => n276, A2 => n275, ZN => Y(4));
   U183 : AOI22_X1 port map( A1 => A_neg(4), A2 => n154, B1 => A_signal(4), B2 
                           => n145, ZN => n276);
   U184 : AOI222_X1 port map( A1 => A_shifted(4), A2 => n181, B1 => 
                           zeroSignal(4), B2 => n171, C1 => A_neg_shifted(4), 
                           C2 => n161, ZN => n275);
   U185 : NAND2_X1 port map( A1 => n298, A2 => n297, ZN => Y(5));
   U186 : AOI22_X1 port map( A1 => A_neg(5), A2 => n155, B1 => A_signal(5), B2 
                           => n146, ZN => n298);
   U187 : AOI222_X1 port map( A1 => A_shifted(5), A2 => n182, B1 => 
                           zeroSignal(5), B2 => n172, C1 => A_neg_shifted(5), 
                           C2 => n160, ZN => n297);
   U188 : NAND2_X1 port map( A1 => n308, A2 => n307, ZN => Y(6));
   U189 : AOI22_X1 port map( A1 => A_neg(6), A2 => n156, B1 => A_signal(6), B2 
                           => n147, ZN => n308);
   U190 : AOI222_X1 port map( A1 => A_shifted(6), A2 => n182, B1 => 
                           zeroSignal(6), B2 => n173, C1 => A_neg_shifted(6), 
                           C2 => n160, ZN => n307);
   U191 : NAND2_X1 port map( A1 => n310, A2 => n309, ZN => Y(7));
   U192 : AOI22_X1 port map( A1 => A_neg(7), A2 => n156, B1 => A_signal(7), B2 
                           => n147, ZN => n310);
   U193 : AOI222_X1 port map( A1 => A_shifted(7), A2 => n182, B1 => 
                           zeroSignal(7), B2 => n173, C1 => A_neg_shifted(7), 
                           C2 => n160, ZN => n309);
   U194 : NAND2_X1 port map( A1 => n312, A2 => n311, ZN => Y(8));
   U195 : AOI22_X1 port map( A1 => A_neg(8), A2 => n156, B1 => A_signal(8), B2 
                           => n147, ZN => n312);
   U196 : AOI222_X1 port map( A1 => A_shifted(8), A2 => n182, B1 => 
                           zeroSignal(8), B2 => n173, C1 => A_neg_shifted(8), 
                           C2 => n160, ZN => n311);
   U197 : NAND2_X1 port map( A1 => n318, A2 => n317, ZN => Y(9));
   U198 : AOI22_X1 port map( A1 => A_neg(9), A2 => n156, B1 => A_signal(9), B2 
                           => n147, ZN => n318);
   U199 : AOI222_X1 port map( A1 => A_shifted(9), A2 => n182, B1 => 
                           zeroSignal(9), B2 => n173, C1 => A_neg_shifted(9), 
                           C2 => n160, ZN => n317);
   U200 : NAND2_X1 port map( A1 => n190, A2 => n189, ZN => Y(10));
   U201 : AOI22_X1 port map( A1 => A_neg(10), A2 => n151, B1 => A_signal(10), 
                           B2 => n142, ZN => n190);
   U202 : AOI222_X1 port map( A1 => A_shifted(10), A2 => n177, B1 => 
                           zeroSignal(10), B2 => n168, C1 => A_neg_shifted(10),
                           C2 => n165, ZN => n189);
   U203 : NAND2_X1 port map( A1 => n192, A2 => n191, ZN => Y(11));
   U204 : AOI22_X1 port map( A1 => A_neg(11), A2 => n151, B1 => A_signal(11), 
                           B2 => n142, ZN => n192);
   U205 : AOI222_X1 port map( A1 => A_shifted(11), A2 => n177, B1 => 
                           zeroSignal(11), B2 => n168, C1 => A_neg_shifted(11),
                           C2 => n165, ZN => n191);
   U206 : NAND2_X1 port map( A1 => n194, A2 => n193, ZN => Y(12));
   U207 : AOI22_X1 port map( A1 => A_neg(12), A2 => n151, B1 => A_signal(12), 
                           B2 => n142, ZN => n194);
   U208 : AOI222_X1 port map( A1 => A_shifted(12), A2 => n177, B1 => 
                           zeroSignal(12), B2 => n168, C1 => A_neg_shifted(12),
                           C2 => n165, ZN => n193);
   U209 : NAND2_X1 port map( A1 => n196, A2 => n195, ZN => Y(13));
   U210 : AOI22_X1 port map( A1 => A_neg(13), A2 => n151, B1 => A_signal(13), 
                           B2 => n142, ZN => n196);
   U211 : AOI222_X1 port map( A1 => A_shifted(13), A2 => n177, B1 => 
                           zeroSignal(13), B2 => n168, C1 => A_neg_shifted(13),
                           C2 => n164, ZN => n195);
   U212 : NAND2_X1 port map( A1 => n198, A2 => n197, ZN => Y(14));
   U213 : AOI22_X1 port map( A1 => A_neg(14), A2 => n151, B1 => A_signal(14), 
                           B2 => n142, ZN => n198);
   U214 : AOI222_X1 port map( A1 => A_shifted(14), A2 => n177, B1 => 
                           zeroSignal(14), B2 => n168, C1 => A_neg_shifted(14),
                           C2 => n164, ZN => n197);
   U215 : NAND2_X1 port map( A1 => n200, A2 => n199, ZN => Y(15));
   U216 : AOI22_X1 port map( A1 => A_neg(15), A2 => n151, B1 => A_signal(15), 
                           B2 => n142, ZN => n200);
   U217 : AOI222_X1 port map( A1 => A_shifted(15), A2 => n177, B1 => 
                           zeroSignal(15), B2 => n168, C1 => A_neg_shifted(15),
                           C2 => n164, ZN => n199);
   U218 : NAND2_X1 port map( A1 => n202, A2 => n201, ZN => Y(16));
   U219 : AOI22_X1 port map( A1 => A_neg(16), A2 => n151, B1 => A_signal(16), 
                           B2 => n142, ZN => n202);
   U220 : AOI222_X1 port map( A1 => A_shifted(16), A2 => n177, B1 => 
                           zeroSignal(16), B2 => n168, C1 => A_neg_shifted(16),
                           C2 => n164, ZN => n201);
   U221 : NAND2_X1 port map( A1 => n204, A2 => n203, ZN => Y(17));
   U222 : AOI22_X1 port map( A1 => A_neg(17), A2 => n151, B1 => A_signal(17), 
                           B2 => n142, ZN => n204);
   U223 : AOI222_X1 port map( A1 => A_shifted(17), A2 => n177, B1 => 
                           zeroSignal(17), B2 => n168, C1 => A_neg_shifted(17),
                           C2 => n164, ZN => n203);
   U224 : NAND2_X1 port map( A1 => n206, A2 => n205, ZN => Y(18));
   U225 : AOI22_X1 port map( A1 => A_neg(18), A2 => n151, B1 => A_signal(18), 
                           B2 => n142, ZN => n206);
   U226 : AOI222_X1 port map( A1 => A_shifted(18), A2 => n177, B1 => 
                           zeroSignal(18), B2 => n168, C1 => A_neg_shifted(18),
                           C2 => n164, ZN => n205);
   U227 : NAND2_X1 port map( A1 => n208, A2 => n207, ZN => Y(19));
   U228 : AOI22_X1 port map( A1 => A_neg(19), A2 => n151, B1 => A_signal(19), 
                           B2 => n142, ZN => n208);
   U229 : AOI222_X1 port map( A1 => A_shifted(19), A2 => n177, B1 => 
                           zeroSignal(19), B2 => n168, C1 => A_neg_shifted(19),
                           C2 => n164, ZN => n207);
   U230 : NAND2_X1 port map( A1 => n212, A2 => n211, ZN => Y(20));
   U231 : AOI22_X1 port map( A1 => A_neg(20), A2 => n152, B1 => A_signal(20), 
                           B2 => n143, ZN => n212);
   U232 : AOI222_X1 port map( A1 => A_shifted(20), A2 => n178, B1 => 
                           zeroSignal(20), B2 => n169, C1 => A_neg_shifted(20),
                           C2 => n164, ZN => n211);
   U233 : NAND2_X1 port map( A1 => n214, A2 => n213, ZN => Y(21));
   U234 : AOI22_X1 port map( A1 => A_neg(21), A2 => n152, B1 => A_signal(21), 
                           B2 => n143, ZN => n214);
   U235 : AOI222_X1 port map( A1 => A_shifted(21), A2 => n178, B1 => 
                           zeroSignal(21), B2 => n169, C1 => A_neg_shifted(21),
                           C2 => n164, ZN => n213);
   U236 : NAND2_X1 port map( A1 => n216, A2 => n215, ZN => Y(22));
   U237 : AOI22_X1 port map( A1 => A_neg(22), A2 => n152, B1 => A_signal(22), 
                           B2 => n143, ZN => n216);
   U238 : AOI222_X1 port map( A1 => A_shifted(22), A2 => n178, B1 => 
                           zeroSignal(22), B2 => n169, C1 => A_neg_shifted(22),
                           C2 => n164, ZN => n215);
   U239 : NAND2_X1 port map( A1 => n218, A2 => n217, ZN => Y(23));
   U240 : AOI22_X1 port map( A1 => A_neg(23), A2 => n152, B1 => A_signal(23), 
                           B2 => n143, ZN => n218);
   U241 : AOI222_X1 port map( A1 => A_shifted(23), A2 => n178, B1 => 
                           zeroSignal(23), B2 => n169, C1 => A_neg_shifted(23),
                           C2 => n164, ZN => n217);
   U242 : AOI22_X1 port map( A1 => A_neg(30), A2 => n152, B1 => A_signal(30), 
                           B2 => n143, ZN => n234);
   U243 : AOI22_X1 port map( A1 => A_neg(29), A2 => n152, B1 => A_signal(29), 
                           B2 => n143, ZN => n230);
   U244 : AOI22_X1 port map( A1 => A_neg(27), A2 => n152, B1 => A_signal(27), 
                           B2 => n143, ZN => n226);

end SYN_BEHAVIORAL_2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity MUX51_MuxNbit64_3 is

   port( zeroSignal, A_signal, A_neg, A_shifted, A_neg_shifted : in 
         std_logic_vector (63 downto 0);  Sel : in std_logic_vector (2 downto 
         0);  Y : out std_logic_vector (63 downto 0));

end MUX51_MuxNbit64_3;

architecture SYN_BEHAVIORAL_2 of MUX51_MuxNbit64_3 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, 
      n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, 
      n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, 
      n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, 
      n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, 
      n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, 
      n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, 
      n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, 
      n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, 
      n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, 
      n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, 
      n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, 
      n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, 
      n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, 
      n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, 
      n320 : std_logic;

begin
   
   U1 : AND3_X1 port map( A1 => n319, A2 => n320, A3 => Sel(2), ZN => n141);
   U2 : BUF_X1 port map( A => n141, Z => n166);
   U3 : BUF_X1 port map( A => n159, Z => n158);
   U4 : BUF_X1 port map( A => n185, Z => n184);
   U5 : BUF_X1 port map( A => n150, Z => n149);
   U6 : BUF_X1 port map( A => n141, Z => n167);
   U7 : BUF_X1 port map( A => n185, Z => n183);
   U8 : BUF_X1 port map( A => n159, Z => n157);
   U9 : BUF_X1 port map( A => n150, Z => n148);
   U10 : BUF_X1 port map( A => n176, Z => n175);
   U11 : BUF_X1 port map( A => n176, Z => n174);
   U12 : BUF_X1 port map( A => n184, Z => n178);
   U13 : BUF_X1 port map( A => n158, Z => n152);
   U14 : BUF_X1 port map( A => n149, Z => n143);
   U15 : BUF_X1 port map( A => n166, Z => n163);
   U16 : BUF_X1 port map( A => n184, Z => n179);
   U17 : BUF_X1 port map( A => n158, Z => n153);
   U18 : BUF_X1 port map( A => n149, Z => n144);
   U19 : BUF_X1 port map( A => n167, Z => n162);
   U20 : BUF_X1 port map( A => n183, Z => n180);
   U21 : BUF_X1 port map( A => n157, Z => n154);
   U22 : BUF_X1 port map( A => n148, Z => n145);
   U23 : BUF_X1 port map( A => n167, Z => n161);
   U24 : BUF_X1 port map( A => n183, Z => n181);
   U25 : BUF_X1 port map( A => n157, Z => n155);
   U26 : BUF_X1 port map( A => n148, Z => n146);
   U27 : BUF_X1 port map( A => n167, Z => n160);
   U28 : BUF_X1 port map( A => n183, Z => n182);
   U29 : BUF_X1 port map( A => n158, Z => n151);
   U30 : BUF_X1 port map( A => n149, Z => n142);
   U31 : BUF_X1 port map( A => n175, Z => n168);
   U32 : BUF_X1 port map( A => n175, Z => n169);
   U33 : BUF_X1 port map( A => n175, Z => n170);
   U34 : BUF_X1 port map( A => n174, Z => n171);
   U35 : BUF_X1 port map( A => n174, Z => n172);
   U36 : BUF_X1 port map( A => n166, Z => n164);
   U37 : BUF_X1 port map( A => n184, Z => n177);
   U38 : BUF_X1 port map( A => n166, Z => n165);
   U39 : BUF_X1 port map( A => n157, Z => n156);
   U40 : BUF_X1 port map( A => n148, Z => n147);
   U41 : BUF_X1 port map( A => n174, Z => n173);
   U42 : INV_X1 port map( A => Sel(1), ZN => n320);
   U43 : BUF_X1 port map( A => n316, Z => n185);
   U44 : NOR3_X1 port map( A1 => n319, A2 => Sel(2), A3 => n320, ZN => n316);
   U45 : BUF_X1 port map( A => n314, Z => n159);
   U46 : NOR3_X1 port map( A1 => Sel(0), A2 => Sel(2), A3 => n320, ZN => n314);
   U47 : INV_X1 port map( A => Sel(0), ZN => n319);
   U48 : BUF_X1 port map( A => n313, Z => n150);
   U49 : NOR3_X1 port map( A1 => Sel(1), A2 => Sel(2), A3 => n319, ZN => n313);
   U50 : BUF_X1 port map( A => n315, Z => n176);
   U51 : NOR2_X1 port map( A1 => n165, A2 => n186, ZN => n315);
   U52 : AOI21_X1 port map( B1 => n319, B2 => n320, A => Sel(2), ZN => n186);
   U53 : NAND2_X1 port map( A1 => n260, A2 => n259, ZN => Y(42));
   U54 : AOI222_X1 port map( A1 => A_shifted(42), A2 => n180, B1 => 
                           zeroSignal(42), B2 => n171, C1 => A_neg_shifted(42),
                           C2 => n162, ZN => n259);
   U55 : AOI22_X1 port map( A1 => A_neg(42), A2 => n154, B1 => A_signal(42), B2
                           => n145, ZN => n260);
   U56 : NAND2_X1 port map( A1 => n226, A2 => n225, ZN => Y(27));
   U57 : AOI22_X1 port map( A1 => A_neg(27), A2 => n152, B1 => A_signal(27), B2
                           => n143, ZN => n226);
   U58 : AOI222_X1 port map( A1 => A_shifted(27), A2 => n178, B1 => 
                           zeroSignal(27), B2 => n169, C1 => A_neg_shifted(27),
                           C2 => n163, ZN => n225);
   U59 : NAND2_X1 port map( A1 => n224, A2 => n223, ZN => Y(26));
   U60 : AOI222_X1 port map( A1 => A_shifted(26), A2 => n178, B1 => 
                           zeroSignal(26), B2 => n169, C1 => A_neg_shifted(26),
                           C2 => n163, ZN => n223);
   U61 : AOI22_X1 port map( A1 => A_neg(26), A2 => n152, B1 => A_signal(26), B2
                           => n143, ZN => n224);
   U62 : NAND2_X1 port map( A1 => n228, A2 => n227, ZN => Y(28));
   U63 : AOI22_X1 port map( A1 => A_neg(28), A2 => n152, B1 => A_signal(28), B2
                           => n143, ZN => n228);
   U64 : AOI222_X1 port map( A1 => A_shifted(28), A2 => n178, B1 => 
                           zeroSignal(28), B2 => n169, C1 => A_neg_shifted(28),
                           C2 => n163, ZN => n227);
   U65 : NAND2_X1 port map( A1 => n258, A2 => n257, ZN => Y(41));
   U66 : AOI222_X1 port map( A1 => A_shifted(41), A2 => n180, B1 => 
                           zeroSignal(41), B2 => n170, C1 => A_neg_shifted(41),
                           C2 => n162, ZN => n257);
   U67 : AOI22_X1 port map( A1 => A_neg(41), A2 => n153, B1 => A_signal(41), B2
                           => n144, ZN => n258);
   U68 : NAND2_X1 port map( A1 => n252, A2 => n251, ZN => Y(39));
   U69 : AOI222_X1 port map( A1 => A_shifted(39), A2 => n179, B1 => 
                           zeroSignal(39), B2 => n170, C1 => A_neg_shifted(39),
                           C2 => n162, ZN => n251);
   U70 : AOI22_X1 port map( A1 => A_neg(39), A2 => n153, B1 => A_signal(39), B2
                           => n144, ZN => n252);
   U71 : NAND2_X1 port map( A1 => n256, A2 => n255, ZN => Y(40));
   U72 : AOI222_X1 port map( A1 => A_shifted(40), A2 => n180, B1 => 
                           zeroSignal(40), B2 => n170, C1 => A_neg_shifted(40),
                           C2 => n162, ZN => n255);
   U73 : AOI22_X1 port map( A1 => A_neg(40), A2 => n153, B1 => A_signal(40), B2
                           => n144, ZN => n256);
   U74 : NAND2_X1 port map( A1 => n262, A2 => n261, ZN => Y(43));
   U75 : AOI222_X1 port map( A1 => A_shifted(43), A2 => n180, B1 => 
                           zeroSignal(43), B2 => n171, C1 => A_neg_shifted(43),
                           C2 => n162, ZN => n261);
   U76 : AOI22_X1 port map( A1 => A_neg(43), A2 => n154, B1 => A_signal(43), B2
                           => n145, ZN => n262);
   U77 : NAND2_X1 port map( A1 => n266, A2 => n265, ZN => Y(45));
   U78 : AOI222_X1 port map( A1 => A_shifted(45), A2 => n180, B1 => 
                           zeroSignal(45), B2 => n171, C1 => A_neg_shifted(45),
                           C2 => n162, ZN => n265);
   U79 : AOI22_X1 port map( A1 => A_neg(45), A2 => n154, B1 => A_signal(45), B2
                           => n145, ZN => n266);
   U80 : NAND2_X1 port map( A1 => n268, A2 => n267, ZN => Y(46));
   U81 : AOI222_X1 port map( A1 => A_shifted(46), A2 => n180, B1 => 
                           zeroSignal(46), B2 => n171, C1 => A_neg_shifted(46),
                           C2 => n161, ZN => n267);
   U82 : AOI22_X1 port map( A1 => A_neg(46), A2 => n154, B1 => A_signal(46), B2
                           => n145, ZN => n268);
   U83 : NAND2_X1 port map( A1 => n270, A2 => n269, ZN => Y(47));
   U84 : AOI222_X1 port map( A1 => A_shifted(47), A2 => n180, B1 => 
                           zeroSignal(47), B2 => n171, C1 => A_neg_shifted(47),
                           C2 => n161, ZN => n269);
   U85 : AOI22_X1 port map( A1 => A_neg(47), A2 => n154, B1 => A_signal(47), B2
                           => n145, ZN => n270);
   U86 : NAND2_X1 port map( A1 => n272, A2 => n271, ZN => Y(48));
   U87 : AOI222_X1 port map( A1 => A_shifted(48), A2 => n180, B1 => 
                           zeroSignal(48), B2 => n171, C1 => A_neg_shifted(48),
                           C2 => n161, ZN => n271);
   U88 : AOI22_X1 port map( A1 => A_neg(48), A2 => n154, B1 => A_signal(48), B2
                           => n145, ZN => n272);
   U89 : NAND2_X1 port map( A1 => n274, A2 => n273, ZN => Y(49));
   U90 : AOI222_X1 port map( A1 => A_shifted(49), A2 => n180, B1 => 
                           zeroSignal(49), B2 => n171, C1 => A_neg_shifted(49),
                           C2 => n161, ZN => n273);
   U91 : AOI22_X1 port map( A1 => A_neg(49), A2 => n154, B1 => A_signal(49), B2
                           => n145, ZN => n274);
   U92 : NAND2_X1 port map( A1 => n278, A2 => n277, ZN => Y(50));
   U93 : AOI222_X1 port map( A1 => A_shifted(50), A2 => n181, B1 => 
                           zeroSignal(50), B2 => n171, C1 => A_neg_shifted(50),
                           C2 => n161, ZN => n277);
   U94 : AOI22_X1 port map( A1 => A_neg(50), A2 => n154, B1 => A_signal(50), B2
                           => n145, ZN => n278);
   U95 : NAND2_X1 port map( A1 => n280, A2 => n279, ZN => Y(51));
   U96 : AOI222_X1 port map( A1 => A_shifted(51), A2 => n181, B1 => 
                           zeroSignal(51), B2 => n171, C1 => A_neg_shifted(51),
                           C2 => n161, ZN => n279);
   U97 : AOI22_X1 port map( A1 => A_neg(51), A2 => n154, B1 => A_signal(51), B2
                           => n145, ZN => n280);
   U98 : NAND2_X1 port map( A1 => n230, A2 => n229, ZN => Y(29));
   U99 : AOI222_X1 port map( A1 => A_shifted(29), A2 => n178, B1 => 
                           zeroSignal(29), B2 => n169, C1 => A_neg_shifted(29),
                           C2 => n163, ZN => n229);
   U100 : NAND2_X1 port map( A1 => n282, A2 => n281, ZN => Y(52));
   U101 : AOI222_X1 port map( A1 => A_shifted(52), A2 => n181, B1 => 
                           zeroSignal(52), B2 => n171, C1 => A_neg_shifted(52),
                           C2 => n161, ZN => n281);
   U102 : AOI22_X1 port map( A1 => A_neg(52), A2 => n154, B1 => A_signal(52), 
                           B2 => n145, ZN => n282);
   U103 : NAND2_X1 port map( A1 => n284, A2 => n283, ZN => Y(53));
   U104 : AOI222_X1 port map( A1 => A_shifted(53), A2 => n181, B1 => 
                           zeroSignal(53), B2 => n172, C1 => A_neg_shifted(53),
                           C2 => n161, ZN => n283);
   U105 : AOI22_X1 port map( A1 => A_neg(53), A2 => n155, B1 => A_signal(53), 
                           B2 => n146, ZN => n284);
   U106 : NAND2_X1 port map( A1 => n286, A2 => n285, ZN => Y(54));
   U107 : AOI222_X1 port map( A1 => A_shifted(54), A2 => n181, B1 => 
                           zeroSignal(54), B2 => n172, C1 => A_neg_shifted(54),
                           C2 => n161, ZN => n285);
   U108 : AOI22_X1 port map( A1 => A_neg(54), A2 => n155, B1 => A_signal(54), 
                           B2 => n146, ZN => n286);
   U109 : NAND2_X1 port map( A1 => n264, A2 => n263, ZN => Y(44));
   U110 : AOI22_X1 port map( A1 => A_neg(44), A2 => n154, B1 => A_signal(44), 
                           B2 => n145, ZN => n264);
   U111 : AOI222_X1 port map( A1 => A_shifted(44), A2 => n180, B1 => 
                           zeroSignal(44), B2 => n171, C1 => A_neg_shifted(44),
                           C2 => n162, ZN => n263);
   U112 : NAND2_X1 port map( A1 => n290, A2 => n289, ZN => Y(56));
   U113 : AOI222_X1 port map( A1 => A_shifted(56), A2 => n181, B1 => 
                           zeroSignal(56), B2 => n172, C1 => A_neg_shifted(56),
                           C2 => n161, ZN => n289);
   U114 : AOI22_X1 port map( A1 => A_neg(56), A2 => n155, B1 => A_signal(56), 
                           B2 => n146, ZN => n290);
   U115 : NAND2_X1 port map( A1 => n292, A2 => n291, ZN => Y(57));
   U116 : AOI222_X1 port map( A1 => A_shifted(57), A2 => n181, B1 => 
                           zeroSignal(57), B2 => n172, C1 => A_neg_shifted(57),
                           C2 => n160, ZN => n291);
   U117 : AOI22_X1 port map( A1 => A_neg(57), A2 => n155, B1 => A_signal(57), 
                           B2 => n146, ZN => n292);
   U118 : NAND2_X1 port map( A1 => n294, A2 => n293, ZN => Y(58));
   U119 : AOI222_X1 port map( A1 => A_shifted(58), A2 => n181, B1 => 
                           zeroSignal(58), B2 => n172, C1 => A_neg_shifted(58),
                           C2 => n160, ZN => n293);
   U120 : AOI22_X1 port map( A1 => A_neg(58), A2 => n155, B1 => A_signal(58), 
                           B2 => n146, ZN => n294);
   U121 : NAND2_X1 port map( A1 => n246, A2 => n245, ZN => Y(36));
   U122 : AOI222_X1 port map( A1 => A_shifted(36), A2 => n179, B1 => 
                           zeroSignal(36), B2 => n170, C1 => A_neg_shifted(36),
                           C2 => n162, ZN => n245);
   U123 : AOI22_X1 port map( A1 => A_neg(36), A2 => n153, B1 => A_signal(36), 
                           B2 => n144, ZN => n246);
   U124 : NAND2_X1 port map( A1 => n234, A2 => n233, ZN => Y(30));
   U125 : AOI22_X1 port map( A1 => A_neg(30), A2 => n152, B1 => A_signal(30), 
                           B2 => n143, ZN => n234);
   U126 : AOI222_X1 port map( A1 => A_shifted(30), A2 => n179, B1 => 
                           zeroSignal(30), B2 => n169, C1 => A_neg_shifted(30),
                           C2 => n163, ZN => n233);
   U127 : NAND2_X1 port map( A1 => n250, A2 => n249, ZN => Y(38));
   U128 : AOI222_X1 port map( A1 => A_shifted(38), A2 => n179, B1 => 
                           zeroSignal(38), B2 => n170, C1 => A_neg_shifted(38),
                           C2 => n162, ZN => n249);
   U129 : AOI22_X1 port map( A1 => A_neg(38), A2 => n153, B1 => A_signal(38), 
                           B2 => n144, ZN => n250);
   U130 : NAND2_X1 port map( A1 => n296, A2 => n295, ZN => Y(59));
   U131 : AOI222_X1 port map( A1 => A_shifted(59), A2 => n181, B1 => 
                           zeroSignal(59), B2 => n172, C1 => A_neg_shifted(59),
                           C2 => n160, ZN => n295);
   U132 : AOI22_X1 port map( A1 => A_neg(59), A2 => n155, B1 => A_signal(59), 
                           B2 => n146, ZN => n296);
   U133 : NAND2_X1 port map( A1 => n288, A2 => n287, ZN => Y(55));
   U134 : AOI22_X1 port map( A1 => A_neg(55), A2 => n155, B1 => A_signal(55), 
                           B2 => n146, ZN => n288);
   U135 : AOI222_X1 port map( A1 => A_shifted(55), A2 => n181, B1 => 
                           zeroSignal(55), B2 => n172, C1 => A_neg_shifted(55),
                           C2 => n161, ZN => n287);
   U136 : NAND2_X1 port map( A1 => n248, A2 => n247, ZN => Y(37));
   U137 : AOI22_X1 port map( A1 => A_neg(37), A2 => n153, B1 => A_signal(37), 
                           B2 => n144, ZN => n248);
   U138 : AOI222_X1 port map( A1 => A_shifted(37), A2 => n179, B1 => 
                           zeroSignal(37), B2 => n170, C1 => A_neg_shifted(37),
                           C2 => n162, ZN => n247);
   U139 : NAND2_X1 port map( A1 => n300, A2 => n299, ZN => Y(60));
   U140 : AOI222_X1 port map( A1 => A_shifted(60), A2 => n182, B1 => 
                           zeroSignal(60), B2 => n172, C1 => A_neg_shifted(60),
                           C2 => n160, ZN => n299);
   U141 : AOI22_X1 port map( A1 => A_neg(60), A2 => n155, B1 => A_signal(60), 
                           B2 => n146, ZN => n300);
   U142 : NAND2_X1 port map( A1 => n302, A2 => n301, ZN => Y(61));
   U143 : AOI222_X1 port map( A1 => A_shifted(61), A2 => n182, B1 => 
                           zeroSignal(61), B2 => n172, C1 => A_neg_shifted(61),
                           C2 => n160, ZN => n301);
   U144 : AOI22_X1 port map( A1 => A_neg(61), A2 => n155, B1 => A_signal(61), 
                           B2 => n146, ZN => n302);
   U145 : NAND2_X1 port map( A1 => n304, A2 => n303, ZN => Y(62));
   U146 : AOI222_X1 port map( A1 => A_shifted(62), A2 => n182, B1 => 
                           zeroSignal(62), B2 => n172, C1 => A_neg_shifted(62),
                           C2 => n160, ZN => n303);
   U147 : AOI22_X1 port map( A1 => A_neg(62), A2 => n155, B1 => A_signal(62), 
                           B2 => n146, ZN => n304);
   U148 : NAND2_X1 port map( A1 => n242, A2 => n241, ZN => Y(34));
   U149 : AOI222_X1 port map( A1 => A_shifted(34), A2 => n179, B1 => 
                           zeroSignal(34), B2 => n170, C1 => A_neg_shifted(34),
                           C2 => n163, ZN => n241);
   U150 : AOI22_X1 port map( A1 => A_neg(34), A2 => n153, B1 => A_signal(34), 
                           B2 => n144, ZN => n242);
   U151 : NAND2_X1 port map( A1 => n236, A2 => n235, ZN => Y(31));
   U152 : AOI222_X1 port map( A1 => A_shifted(31), A2 => n179, B1 => 
                           zeroSignal(31), B2 => n170, C1 => A_neg_shifted(31),
                           C2 => n163, ZN => n235);
   U153 : NAND2_X1 port map( A1 => n306, A2 => n305, ZN => Y(63));
   U154 : AOI222_X1 port map( A1 => A_shifted(63), A2 => n182, B1 => 
                           zeroSignal(63), B2 => n172, C1 => A_neg_shifted(63),
                           C2 => n160, ZN => n305);
   U155 : AOI22_X1 port map( A1 => A_neg(63), A2 => n155, B1 => A_signal(63), 
                           B2 => n146, ZN => n306);
   U156 : NAND2_X1 port map( A1 => n240, A2 => n239, ZN => Y(33));
   U157 : AOI222_X1 port map( A1 => A_shifted(33), A2 => n179, B1 => 
                           zeroSignal(33), B2 => n170, C1 => A_neg_shifted(33),
                           C2 => n163, ZN => n239);
   U158 : AOI22_X1 port map( A1 => A_neg(33), A2 => n153, B1 => A_signal(33), 
                           B2 => n144, ZN => n240);
   U159 : NAND2_X1 port map( A1 => n244, A2 => n243, ZN => Y(35));
   U160 : AOI222_X1 port map( A1 => A_shifted(35), A2 => n179, B1 => 
                           zeroSignal(35), B2 => n170, C1 => A_neg_shifted(35),
                           C2 => n162, ZN => n243);
   U161 : AOI22_X1 port map( A1 => A_neg(35), A2 => n153, B1 => A_signal(35), 
                           B2 => n144, ZN => n244);
   U162 : NAND2_X1 port map( A1 => n238, A2 => n237, ZN => Y(32));
   U163 : AOI222_X1 port map( A1 => A_shifted(32), A2 => n179, B1 => 
                           zeroSignal(32), B2 => n170, C1 => A_neg_shifted(32),
                           C2 => n163, ZN => n237);
   U164 : NAND2_X1 port map( A1 => n188, A2 => n187, ZN => Y(0));
   U165 : AOI22_X1 port map( A1 => A_neg(0), A2 => n151, B1 => A_signal(0), B2 
                           => n142, ZN => n188);
   U166 : AOI222_X1 port map( A1 => A_shifted(0), A2 => n177, B1 => 
                           zeroSignal(0), B2 => n168, C1 => A_neg_shifted(0), 
                           C2 => n165, ZN => n187);
   U167 : NAND2_X1 port map( A1 => n210, A2 => n209, ZN => Y(1));
   U168 : AOI22_X1 port map( A1 => A_neg(1), A2 => n151, B1 => A_signal(1), B2 
                           => n142, ZN => n210);
   U169 : AOI222_X1 port map( A1 => A_shifted(1), A2 => n178, B1 => 
                           zeroSignal(1), B2 => n168, C1 => A_neg_shifted(1), 
                           C2 => n164, ZN => n209);
   U170 : NAND2_X1 port map( A1 => n232, A2 => n231, ZN => Y(2));
   U171 : AOI22_X1 port map( A1 => A_neg(2), A2 => n152, B1 => A_signal(2), B2 
                           => n143, ZN => n232);
   U172 : AOI222_X1 port map( A1 => A_shifted(2), A2 => n179, B1 => 
                           zeroSignal(2), B2 => n169, C1 => A_neg_shifted(2), 
                           C2 => n163, ZN => n231);
   U173 : NAND2_X1 port map( A1 => n254, A2 => n253, ZN => Y(3));
   U174 : AOI22_X1 port map( A1 => A_neg(3), A2 => n153, B1 => A_signal(3), B2 
                           => n144, ZN => n254);
   U175 : AOI222_X1 port map( A1 => A_shifted(3), A2 => n180, B1 => 
                           zeroSignal(3), B2 => n170, C1 => A_neg_shifted(3), 
                           C2 => n162, ZN => n253);
   U176 : NAND2_X1 port map( A1 => n276, A2 => n275, ZN => Y(4));
   U177 : AOI22_X1 port map( A1 => A_neg(4), A2 => n154, B1 => A_signal(4), B2 
                           => n145, ZN => n276);
   U178 : AOI222_X1 port map( A1 => A_shifted(4), A2 => n181, B1 => 
                           zeroSignal(4), B2 => n171, C1 => A_neg_shifted(4), 
                           C2 => n161, ZN => n275);
   U179 : NAND2_X1 port map( A1 => n298, A2 => n297, ZN => Y(5));
   U180 : AOI22_X1 port map( A1 => A_neg(5), A2 => n155, B1 => A_signal(5), B2 
                           => n146, ZN => n298);
   U181 : AOI222_X1 port map( A1 => A_shifted(5), A2 => n182, B1 => 
                           zeroSignal(5), B2 => n172, C1 => A_neg_shifted(5), 
                           C2 => n160, ZN => n297);
   U182 : NAND2_X1 port map( A1 => n308, A2 => n307, ZN => Y(6));
   U183 : AOI22_X1 port map( A1 => A_neg(6), A2 => n156, B1 => A_signal(6), B2 
                           => n147, ZN => n308);
   U184 : AOI222_X1 port map( A1 => A_shifted(6), A2 => n182, B1 => 
                           zeroSignal(6), B2 => n173, C1 => A_neg_shifted(6), 
                           C2 => n160, ZN => n307);
   U185 : NAND2_X1 port map( A1 => n310, A2 => n309, ZN => Y(7));
   U186 : AOI22_X1 port map( A1 => A_neg(7), A2 => n156, B1 => A_signal(7), B2 
                           => n147, ZN => n310);
   U187 : AOI222_X1 port map( A1 => A_shifted(7), A2 => n182, B1 => 
                           zeroSignal(7), B2 => n173, C1 => A_neg_shifted(7), 
                           C2 => n160, ZN => n309);
   U188 : NAND2_X1 port map( A1 => n312, A2 => n311, ZN => Y(8));
   U189 : AOI22_X1 port map( A1 => A_neg(8), A2 => n156, B1 => A_signal(8), B2 
                           => n147, ZN => n312);
   U190 : AOI222_X1 port map( A1 => A_shifted(8), A2 => n182, B1 => 
                           zeroSignal(8), B2 => n173, C1 => A_neg_shifted(8), 
                           C2 => n160, ZN => n311);
   U191 : NAND2_X1 port map( A1 => n318, A2 => n317, ZN => Y(9));
   U192 : AOI22_X1 port map( A1 => A_neg(9), A2 => n156, B1 => A_signal(9), B2 
                           => n147, ZN => n318);
   U193 : AOI222_X1 port map( A1 => A_shifted(9), A2 => n182, B1 => 
                           zeroSignal(9), B2 => n173, C1 => A_neg_shifted(9), 
                           C2 => n160, ZN => n317);
   U194 : NAND2_X1 port map( A1 => n190, A2 => n189, ZN => Y(10));
   U195 : AOI22_X1 port map( A1 => A_neg(10), A2 => n151, B1 => A_signal(10), 
                           B2 => n142, ZN => n190);
   U196 : AOI222_X1 port map( A1 => A_shifted(10), A2 => n177, B1 => 
                           zeroSignal(10), B2 => n168, C1 => A_neg_shifted(10),
                           C2 => n165, ZN => n189);
   U197 : NAND2_X1 port map( A1 => n192, A2 => n191, ZN => Y(11));
   U198 : AOI22_X1 port map( A1 => A_neg(11), A2 => n151, B1 => A_signal(11), 
                           B2 => n142, ZN => n192);
   U199 : AOI222_X1 port map( A1 => A_shifted(11), A2 => n177, B1 => 
                           zeroSignal(11), B2 => n168, C1 => A_neg_shifted(11),
                           C2 => n165, ZN => n191);
   U200 : NAND2_X1 port map( A1 => n194, A2 => n193, ZN => Y(12));
   U201 : AOI22_X1 port map( A1 => A_neg(12), A2 => n151, B1 => A_signal(12), 
                           B2 => n142, ZN => n194);
   U202 : AOI222_X1 port map( A1 => A_shifted(12), A2 => n177, B1 => 
                           zeroSignal(12), B2 => n168, C1 => A_neg_shifted(12),
                           C2 => n165, ZN => n193);
   U203 : NAND2_X1 port map( A1 => n196, A2 => n195, ZN => Y(13));
   U204 : AOI22_X1 port map( A1 => A_neg(13), A2 => n151, B1 => A_signal(13), 
                           B2 => n142, ZN => n196);
   U205 : AOI222_X1 port map( A1 => A_shifted(13), A2 => n177, B1 => 
                           zeroSignal(13), B2 => n168, C1 => A_neg_shifted(13),
                           C2 => n164, ZN => n195);
   U206 : NAND2_X1 port map( A1 => n198, A2 => n197, ZN => Y(14));
   U207 : AOI22_X1 port map( A1 => A_neg(14), A2 => n151, B1 => A_signal(14), 
                           B2 => n142, ZN => n198);
   U208 : AOI222_X1 port map( A1 => A_shifted(14), A2 => n177, B1 => 
                           zeroSignal(14), B2 => n168, C1 => A_neg_shifted(14),
                           C2 => n164, ZN => n197);
   U209 : NAND2_X1 port map( A1 => n200, A2 => n199, ZN => Y(15));
   U210 : AOI22_X1 port map( A1 => A_neg(15), A2 => n151, B1 => A_signal(15), 
                           B2 => n142, ZN => n200);
   U211 : AOI222_X1 port map( A1 => A_shifted(15), A2 => n177, B1 => 
                           zeroSignal(15), B2 => n168, C1 => A_neg_shifted(15),
                           C2 => n164, ZN => n199);
   U212 : NAND2_X1 port map( A1 => n202, A2 => n201, ZN => Y(16));
   U213 : AOI22_X1 port map( A1 => A_neg(16), A2 => n151, B1 => A_signal(16), 
                           B2 => n142, ZN => n202);
   U214 : AOI222_X1 port map( A1 => A_shifted(16), A2 => n177, B1 => 
                           zeroSignal(16), B2 => n168, C1 => A_neg_shifted(16),
                           C2 => n164, ZN => n201);
   U215 : NAND2_X1 port map( A1 => n204, A2 => n203, ZN => Y(17));
   U216 : AOI22_X1 port map( A1 => A_neg(17), A2 => n151, B1 => A_signal(17), 
                           B2 => n142, ZN => n204);
   U217 : AOI222_X1 port map( A1 => A_shifted(17), A2 => n177, B1 => 
                           zeroSignal(17), B2 => n168, C1 => A_neg_shifted(17),
                           C2 => n164, ZN => n203);
   U218 : NAND2_X1 port map( A1 => n206, A2 => n205, ZN => Y(18));
   U219 : AOI22_X1 port map( A1 => A_neg(18), A2 => n151, B1 => A_signal(18), 
                           B2 => n142, ZN => n206);
   U220 : AOI222_X1 port map( A1 => A_shifted(18), A2 => n177, B1 => 
                           zeroSignal(18), B2 => n168, C1 => A_neg_shifted(18),
                           C2 => n164, ZN => n205);
   U221 : NAND2_X1 port map( A1 => n208, A2 => n207, ZN => Y(19));
   U222 : AOI22_X1 port map( A1 => A_neg(19), A2 => n151, B1 => A_signal(19), 
                           B2 => n142, ZN => n208);
   U223 : AOI222_X1 port map( A1 => A_shifted(19), A2 => n177, B1 => 
                           zeroSignal(19), B2 => n168, C1 => A_neg_shifted(19),
                           C2 => n164, ZN => n207);
   U224 : NAND2_X1 port map( A1 => n212, A2 => n211, ZN => Y(20));
   U225 : AOI22_X1 port map( A1 => A_neg(20), A2 => n152, B1 => A_signal(20), 
                           B2 => n143, ZN => n212);
   U226 : AOI222_X1 port map( A1 => A_shifted(20), A2 => n178, B1 => 
                           zeroSignal(20), B2 => n169, C1 => A_neg_shifted(20),
                           C2 => n164, ZN => n211);
   U227 : NAND2_X1 port map( A1 => n214, A2 => n213, ZN => Y(21));
   U228 : AOI22_X1 port map( A1 => A_neg(21), A2 => n152, B1 => A_signal(21), 
                           B2 => n143, ZN => n214);
   U229 : AOI222_X1 port map( A1 => A_shifted(21), A2 => n178, B1 => 
                           zeroSignal(21), B2 => n169, C1 => A_neg_shifted(21),
                           C2 => n164, ZN => n213);
   U230 : NAND2_X1 port map( A1 => n216, A2 => n215, ZN => Y(22));
   U231 : AOI22_X1 port map( A1 => A_neg(22), A2 => n152, B1 => A_signal(22), 
                           B2 => n143, ZN => n216);
   U232 : AOI222_X1 port map( A1 => A_shifted(22), A2 => n178, B1 => 
                           zeroSignal(22), B2 => n169, C1 => A_neg_shifted(22),
                           C2 => n164, ZN => n215);
   U233 : NAND2_X1 port map( A1 => n218, A2 => n217, ZN => Y(23));
   U234 : AOI22_X1 port map( A1 => A_neg(23), A2 => n152, B1 => A_signal(23), 
                           B2 => n143, ZN => n218);
   U235 : AOI222_X1 port map( A1 => A_shifted(23), A2 => n178, B1 => 
                           zeroSignal(23), B2 => n169, C1 => A_neg_shifted(23),
                           C2 => n164, ZN => n217);
   U236 : NAND2_X1 port map( A1 => n220, A2 => n219, ZN => Y(24));
   U237 : AOI22_X1 port map( A1 => A_neg(24), A2 => n152, B1 => A_signal(24), 
                           B2 => n143, ZN => n220);
   U238 : AOI222_X1 port map( A1 => A_shifted(24), A2 => n178, B1 => 
                           zeroSignal(24), B2 => n169, C1 => A_neg_shifted(24),
                           C2 => n163, ZN => n219);
   U239 : NAND2_X1 port map( A1 => n222, A2 => n221, ZN => Y(25));
   U240 : AOI22_X1 port map( A1 => A_neg(25), A2 => n152, B1 => A_signal(25), 
                           B2 => n143, ZN => n222);
   U241 : AOI222_X1 port map( A1 => A_shifted(25), A2 => n178, B1 => 
                           zeroSignal(25), B2 => n169, C1 => A_neg_shifted(25),
                           C2 => n163, ZN => n221);
   U242 : AOI22_X1 port map( A1 => A_neg(32), A2 => n153, B1 => A_signal(32), 
                           B2 => n144, ZN => n238);
   U243 : AOI22_X1 port map( A1 => A_neg(31), A2 => n153, B1 => A_signal(31), 
                           B2 => n144, ZN => n236);
   U244 : AOI22_X1 port map( A1 => A_neg(29), A2 => n152, B1 => A_signal(29), 
                           B2 => n143, ZN => n230);

end SYN_BEHAVIORAL_2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity MUX51_MuxNbit64_2 is

   port( zeroSignal, A_signal, A_neg, A_shifted, A_neg_shifted : in 
         std_logic_vector (63 downto 0);  Sel : in std_logic_vector (2 downto 
         0);  Y : out std_logic_vector (63 downto 0));

end MUX51_MuxNbit64_2;

architecture SYN_BEHAVIORAL_2 of MUX51_MuxNbit64_2 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, 
      n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, 
      n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, 
      n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, 
      n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, 
      n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, 
      n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, 
      n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, 
      n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, 
      n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, 
      n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, 
      n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, 
      n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, 
      n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, 
      n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, 
      n320 : std_logic;

begin
   
   U1 : AND3_X1 port map( A1 => n319, A2 => n320, A3 => Sel(2), ZN => n141);
   U2 : BUF_X1 port map( A => n141, Z => n166);
   U3 : BUF_X1 port map( A => n159, Z => n158);
   U4 : BUF_X1 port map( A => n185, Z => n184);
   U5 : BUF_X1 port map( A => n150, Z => n149);
   U6 : BUF_X1 port map( A => n141, Z => n167);
   U7 : BUF_X1 port map( A => n185, Z => n183);
   U8 : BUF_X1 port map( A => n159, Z => n157);
   U9 : BUF_X1 port map( A => n150, Z => n148);
   U10 : BUF_X1 port map( A => n176, Z => n175);
   U11 : BUF_X1 port map( A => n176, Z => n174);
   U12 : BUF_X1 port map( A => n184, Z => n178);
   U13 : BUF_X1 port map( A => n158, Z => n152);
   U14 : BUF_X1 port map( A => n149, Z => n143);
   U15 : BUF_X1 port map( A => n166, Z => n163);
   U16 : BUF_X1 port map( A => n184, Z => n179);
   U17 : BUF_X1 port map( A => n158, Z => n153);
   U18 : BUF_X1 port map( A => n149, Z => n144);
   U19 : BUF_X1 port map( A => n167, Z => n162);
   U20 : BUF_X1 port map( A => n183, Z => n180);
   U21 : BUF_X1 port map( A => n157, Z => n154);
   U22 : BUF_X1 port map( A => n148, Z => n145);
   U23 : BUF_X1 port map( A => n167, Z => n161);
   U24 : BUF_X1 port map( A => n183, Z => n181);
   U25 : BUF_X1 port map( A => n157, Z => n155);
   U26 : BUF_X1 port map( A => n148, Z => n146);
   U27 : BUF_X1 port map( A => n167, Z => n160);
   U28 : BUF_X1 port map( A => n183, Z => n182);
   U29 : BUF_X1 port map( A => n158, Z => n151);
   U30 : BUF_X1 port map( A => n149, Z => n142);
   U31 : BUF_X1 port map( A => n175, Z => n168);
   U32 : BUF_X1 port map( A => n175, Z => n169);
   U33 : BUF_X1 port map( A => n175, Z => n170);
   U34 : BUF_X1 port map( A => n174, Z => n171);
   U35 : BUF_X1 port map( A => n174, Z => n172);
   U36 : BUF_X1 port map( A => n166, Z => n164);
   U37 : BUF_X1 port map( A => n184, Z => n177);
   U38 : BUF_X1 port map( A => n166, Z => n165);
   U39 : BUF_X1 port map( A => n157, Z => n156);
   U40 : BUF_X1 port map( A => n148, Z => n147);
   U41 : BUF_X1 port map( A => n174, Z => n173);
   U42 : INV_X1 port map( A => Sel(1), ZN => n320);
   U43 : BUF_X1 port map( A => n316, Z => n185);
   U44 : NOR3_X1 port map( A1 => n319, A2 => Sel(2), A3 => n320, ZN => n316);
   U45 : BUF_X1 port map( A => n314, Z => n159);
   U46 : NOR3_X1 port map( A1 => Sel(0), A2 => Sel(2), A3 => n320, ZN => n314);
   U47 : INV_X1 port map( A => Sel(0), ZN => n319);
   U48 : BUF_X1 port map( A => n313, Z => n150);
   U49 : NOR3_X1 port map( A1 => Sel(1), A2 => Sel(2), A3 => n319, ZN => n313);
   U50 : BUF_X1 port map( A => n315, Z => n176);
   U51 : NOR2_X1 port map( A1 => n165, A2 => n186, ZN => n315);
   U52 : AOI21_X1 port map( B1 => n319, B2 => n320, A => Sel(2), ZN => n186);
   U53 : NAND2_X1 port map( A1 => n260, A2 => n259, ZN => Y(42));
   U54 : AOI222_X1 port map( A1 => A_shifted(42), A2 => n180, B1 => 
                           zeroSignal(42), B2 => n171, C1 => A_neg_shifted(42),
                           C2 => n162, ZN => n259);
   U55 : AOI22_X1 port map( A1 => A_neg(42), A2 => n154, B1 => A_signal(42), B2
                           => n145, ZN => n260);
   U56 : NAND2_X1 port map( A1 => n230, A2 => n229, ZN => Y(29));
   U57 : AOI22_X1 port map( A1 => A_neg(29), A2 => n152, B1 => A_signal(29), B2
                           => n143, ZN => n230);
   U58 : AOI222_X1 port map( A1 => A_shifted(29), A2 => n178, B1 => 
                           zeroSignal(29), B2 => n169, C1 => A_neg_shifted(29),
                           C2 => n163, ZN => n229);
   U59 : NAND2_X1 port map( A1 => n228, A2 => n227, ZN => Y(28));
   U60 : AOI222_X1 port map( A1 => A_shifted(28), A2 => n178, B1 => 
                           zeroSignal(28), B2 => n169, C1 => A_neg_shifted(28),
                           C2 => n163, ZN => n227);
   U61 : AOI22_X1 port map( A1 => A_neg(28), A2 => n152, B1 => A_signal(28), B2
                           => n143, ZN => n228);
   U62 : NAND2_X1 port map( A1 => n234, A2 => n233, ZN => Y(30));
   U63 : AOI22_X1 port map( A1 => A_neg(30), A2 => n152, B1 => A_signal(30), B2
                           => n143, ZN => n234);
   U64 : AOI222_X1 port map( A1 => A_shifted(30), A2 => n179, B1 => 
                           zeroSignal(30), B2 => n169, C1 => A_neg_shifted(30),
                           C2 => n163, ZN => n233);
   U65 : NAND2_X1 port map( A1 => n262, A2 => n261, ZN => Y(43));
   U66 : AOI222_X1 port map( A1 => A_shifted(43), A2 => n180, B1 => 
                           zeroSignal(43), B2 => n171, C1 => A_neg_shifted(43),
                           C2 => n162, ZN => n261);
   U67 : AOI22_X1 port map( A1 => A_neg(43), A2 => n154, B1 => A_signal(43), B2
                           => n145, ZN => n262);
   U68 : NAND2_X1 port map( A1 => n258, A2 => n257, ZN => Y(41));
   U69 : AOI222_X1 port map( A1 => A_shifted(41), A2 => n180, B1 => 
                           zeroSignal(41), B2 => n170, C1 => A_neg_shifted(41),
                           C2 => n162, ZN => n257);
   U70 : AOI22_X1 port map( A1 => A_neg(41), A2 => n153, B1 => A_signal(41), B2
                           => n144, ZN => n258);
   U71 : NAND2_X1 port map( A1 => n264, A2 => n263, ZN => Y(44));
   U72 : AOI222_X1 port map( A1 => A_shifted(44), A2 => n180, B1 => 
                           zeroSignal(44), B2 => n171, C1 => A_neg_shifted(44),
                           C2 => n162, ZN => n263);
   U73 : AOI22_X1 port map( A1 => A_neg(44), A2 => n154, B1 => A_signal(44), B2
                           => n145, ZN => n264);
   U74 : NAND2_X1 port map( A1 => n266, A2 => n265, ZN => Y(45));
   U75 : AOI222_X1 port map( A1 => A_shifted(45), A2 => n180, B1 => 
                           zeroSignal(45), B2 => n171, C1 => A_neg_shifted(45),
                           C2 => n162, ZN => n265);
   U76 : AOI22_X1 port map( A1 => A_neg(45), A2 => n154, B1 => A_signal(45), B2
                           => n145, ZN => n266);
   U77 : NAND2_X1 port map( A1 => n270, A2 => n269, ZN => Y(47));
   U78 : AOI222_X1 port map( A1 => A_shifted(47), A2 => n180, B1 => 
                           zeroSignal(47), B2 => n171, C1 => A_neg_shifted(47),
                           C2 => n161, ZN => n269);
   U79 : AOI22_X1 port map( A1 => A_neg(47), A2 => n154, B1 => A_signal(47), B2
                           => n145, ZN => n270);
   U80 : NAND2_X1 port map( A1 => n272, A2 => n271, ZN => Y(48));
   U81 : AOI222_X1 port map( A1 => A_shifted(48), A2 => n180, B1 => 
                           zeroSignal(48), B2 => n171, C1 => A_neg_shifted(48),
                           C2 => n161, ZN => n271);
   U82 : AOI22_X1 port map( A1 => A_neg(48), A2 => n154, B1 => A_signal(48), B2
                           => n145, ZN => n272);
   U83 : NAND2_X1 port map( A1 => n274, A2 => n273, ZN => Y(49));
   U84 : AOI222_X1 port map( A1 => A_shifted(49), A2 => n180, B1 => 
                           zeroSignal(49), B2 => n171, C1 => A_neg_shifted(49),
                           C2 => n161, ZN => n273);
   U85 : AOI22_X1 port map( A1 => A_neg(49), A2 => n154, B1 => A_signal(49), B2
                           => n145, ZN => n274);
   U86 : NAND2_X1 port map( A1 => n278, A2 => n277, ZN => Y(50));
   U87 : AOI222_X1 port map( A1 => A_shifted(50), A2 => n181, B1 => 
                           zeroSignal(50), B2 => n171, C1 => A_neg_shifted(50),
                           C2 => n161, ZN => n277);
   U88 : AOI22_X1 port map( A1 => A_neg(50), A2 => n154, B1 => A_signal(50), B2
                           => n145, ZN => n278);
   U89 : NAND2_X1 port map( A1 => n280, A2 => n279, ZN => Y(51));
   U90 : AOI222_X1 port map( A1 => A_shifted(51), A2 => n181, B1 => 
                           zeroSignal(51), B2 => n171, C1 => A_neg_shifted(51),
                           C2 => n161, ZN => n279);
   U91 : AOI22_X1 port map( A1 => A_neg(51), A2 => n154, B1 => A_signal(51), B2
                           => n145, ZN => n280);
   U92 : NAND2_X1 port map( A1 => n282, A2 => n281, ZN => Y(52));
   U93 : AOI222_X1 port map( A1 => A_shifted(52), A2 => n181, B1 => 
                           zeroSignal(52), B2 => n171, C1 => A_neg_shifted(52),
                           C2 => n161, ZN => n281);
   U94 : AOI22_X1 port map( A1 => A_neg(52), A2 => n154, B1 => A_signal(52), B2
                           => n145, ZN => n282);
   U95 : NAND2_X1 port map( A1 => n284, A2 => n283, ZN => Y(53));
   U96 : AOI222_X1 port map( A1 => A_shifted(53), A2 => n181, B1 => 
                           zeroSignal(53), B2 => n172, C1 => A_neg_shifted(53),
                           C2 => n161, ZN => n283);
   U97 : AOI22_X1 port map( A1 => A_neg(53), A2 => n155, B1 => A_signal(53), B2
                           => n146, ZN => n284);
   U98 : NAND2_X1 port map( A1 => n236, A2 => n235, ZN => Y(31));
   U99 : AOI222_X1 port map( A1 => A_shifted(31), A2 => n179, B1 => 
                           zeroSignal(31), B2 => n170, C1 => A_neg_shifted(31),
                           C2 => n163, ZN => n235);
   U100 : NAND2_X1 port map( A1 => n286, A2 => n285, ZN => Y(54));
   U101 : AOI222_X1 port map( A1 => A_shifted(54), A2 => n181, B1 => 
                           zeroSignal(54), B2 => n172, C1 => A_neg_shifted(54),
                           C2 => n161, ZN => n285);
   U102 : AOI22_X1 port map( A1 => A_neg(54), A2 => n155, B1 => A_signal(54), 
                           B2 => n146, ZN => n286);
   U103 : NAND2_X1 port map( A1 => n288, A2 => n287, ZN => Y(55));
   U104 : AOI222_X1 port map( A1 => A_shifted(55), A2 => n181, B1 => 
                           zeroSignal(55), B2 => n172, C1 => A_neg_shifted(55),
                           C2 => n161, ZN => n287);
   U105 : AOI22_X1 port map( A1 => A_neg(55), A2 => n155, B1 => A_signal(55), 
                           B2 => n146, ZN => n288);
   U106 : NAND2_X1 port map( A1 => n290, A2 => n289, ZN => Y(56));
   U107 : AOI222_X1 port map( A1 => A_shifted(56), A2 => n181, B1 => 
                           zeroSignal(56), B2 => n172, C1 => A_neg_shifted(56),
                           C2 => n161, ZN => n289);
   U108 : AOI22_X1 port map( A1 => A_neg(56), A2 => n155, B1 => A_signal(56), 
                           B2 => n146, ZN => n290);
   U109 : NAND2_X1 port map( A1 => n268, A2 => n267, ZN => Y(46));
   U110 : AOI22_X1 port map( A1 => A_neg(46), A2 => n154, B1 => A_signal(46), 
                           B2 => n145, ZN => n268);
   U111 : AOI222_X1 port map( A1 => A_shifted(46), A2 => n180, B1 => 
                           zeroSignal(46), B2 => n171, C1 => A_neg_shifted(46),
                           C2 => n161, ZN => n267);
   U112 : NAND2_X1 port map( A1 => n294, A2 => n293, ZN => Y(58));
   U113 : AOI222_X1 port map( A1 => A_shifted(58), A2 => n181, B1 => 
                           zeroSignal(58), B2 => n172, C1 => A_neg_shifted(58),
                           C2 => n160, ZN => n293);
   U114 : AOI22_X1 port map( A1 => A_neg(58), A2 => n155, B1 => A_signal(58), 
                           B2 => n146, ZN => n294);
   U115 : NAND2_X1 port map( A1 => n296, A2 => n295, ZN => Y(59));
   U116 : AOI222_X1 port map( A1 => A_shifted(59), A2 => n181, B1 => 
                           zeroSignal(59), B2 => n172, C1 => A_neg_shifted(59),
                           C2 => n160, ZN => n295);
   U117 : AOI22_X1 port map( A1 => A_neg(59), A2 => n155, B1 => A_signal(59), 
                           B2 => n146, ZN => n296);
   U118 : NAND2_X1 port map( A1 => n300, A2 => n299, ZN => Y(60));
   U119 : AOI222_X1 port map( A1 => A_shifted(60), A2 => n182, B1 => 
                           zeroSignal(60), B2 => n172, C1 => A_neg_shifted(60),
                           C2 => n160, ZN => n299);
   U120 : AOI22_X1 port map( A1 => A_neg(60), A2 => n155, B1 => A_signal(60), 
                           B2 => n146, ZN => n300);
   U121 : NAND2_X1 port map( A1 => n250, A2 => n249, ZN => Y(38));
   U122 : AOI222_X1 port map( A1 => A_shifted(38), A2 => n179, B1 => 
                           zeroSignal(38), B2 => n170, C1 => A_neg_shifted(38),
                           C2 => n162, ZN => n249);
   U123 : AOI22_X1 port map( A1 => A_neg(38), A2 => n153, B1 => A_signal(38), 
                           B2 => n144, ZN => n250);
   U124 : NAND2_X1 port map( A1 => n256, A2 => n255, ZN => Y(40));
   U125 : AOI222_X1 port map( A1 => A_shifted(40), A2 => n180, B1 => 
                           zeroSignal(40), B2 => n170, C1 => A_neg_shifted(40),
                           C2 => n162, ZN => n255);
   U126 : AOI22_X1 port map( A1 => A_neg(40), A2 => n153, B1 => A_signal(40), 
                           B2 => n144, ZN => n256);
   U127 : NAND2_X1 port map( A1 => n302, A2 => n301, ZN => Y(61));
   U128 : AOI222_X1 port map( A1 => A_shifted(61), A2 => n182, B1 => 
                           zeroSignal(61), B2 => n172, C1 => A_neg_shifted(61),
                           C2 => n160, ZN => n301);
   U129 : AOI22_X1 port map( A1 => A_neg(61), A2 => n155, B1 => A_signal(61), 
                           B2 => n146, ZN => n302);
   U130 : NAND2_X1 port map( A1 => n238, A2 => n237, ZN => Y(32));
   U131 : AOI22_X1 port map( A1 => A_neg(32), A2 => n153, B1 => A_signal(32), 
                           B2 => n144, ZN => n238);
   U132 : AOI222_X1 port map( A1 => A_shifted(32), A2 => n179, B1 => 
                           zeroSignal(32), B2 => n170, C1 => A_neg_shifted(32),
                           C2 => n163, ZN => n237);
   U133 : NAND2_X1 port map( A1 => n292, A2 => n291, ZN => Y(57));
   U134 : AOI22_X1 port map( A1 => A_neg(57), A2 => n155, B1 => A_signal(57), 
                           B2 => n146, ZN => n292);
   U135 : AOI222_X1 port map( A1 => A_shifted(57), A2 => n181, B1 => 
                           zeroSignal(57), B2 => n172, C1 => A_neg_shifted(57),
                           C2 => n160, ZN => n291);
   U136 : NAND2_X1 port map( A1 => n252, A2 => n251, ZN => Y(39));
   U137 : AOI22_X1 port map( A1 => A_neg(39), A2 => n153, B1 => A_signal(39), 
                           B2 => n144, ZN => n252);
   U138 : AOI222_X1 port map( A1 => A_shifted(39), A2 => n179, B1 => 
                           zeroSignal(39), B2 => n170, C1 => A_neg_shifted(39),
                           C2 => n162, ZN => n251);
   U139 : NAND2_X1 port map( A1 => n304, A2 => n303, ZN => Y(62));
   U140 : AOI222_X1 port map( A1 => A_shifted(62), A2 => n182, B1 => 
                           zeroSignal(62), B2 => n172, C1 => A_neg_shifted(62),
                           C2 => n160, ZN => n303);
   U141 : AOI22_X1 port map( A1 => A_neg(62), A2 => n155, B1 => A_signal(62), 
                           B2 => n146, ZN => n304);
   U142 : NAND2_X1 port map( A1 => n306, A2 => n305, ZN => Y(63));
   U143 : AOI222_X1 port map( A1 => A_shifted(63), A2 => n182, B1 => 
                           zeroSignal(63), B2 => n172, C1 => A_neg_shifted(63),
                           C2 => n160, ZN => n305);
   U144 : AOI22_X1 port map( A1 => A_neg(63), A2 => n155, B1 => A_signal(63), 
                           B2 => n146, ZN => n306);
   U145 : NAND2_X1 port map( A1 => n244, A2 => n243, ZN => Y(35));
   U146 : AOI222_X1 port map( A1 => A_shifted(35), A2 => n179, B1 => 
                           zeroSignal(35), B2 => n170, C1 => A_neg_shifted(35),
                           C2 => n162, ZN => n243);
   U147 : AOI22_X1 port map( A1 => A_neg(35), A2 => n153, B1 => A_signal(35), 
                           B2 => n144, ZN => n244);
   U148 : NAND2_X1 port map( A1 => n246, A2 => n245, ZN => Y(36));
   U149 : AOI222_X1 port map( A1 => A_shifted(36), A2 => n179, B1 => 
                           zeroSignal(36), B2 => n170, C1 => A_neg_shifted(36),
                           C2 => n162, ZN => n245);
   U150 : AOI22_X1 port map( A1 => A_neg(36), A2 => n153, B1 => A_signal(36), 
                           B2 => n144, ZN => n246);
   U151 : NAND2_X1 port map( A1 => n240, A2 => n239, ZN => Y(33));
   U152 : AOI222_X1 port map( A1 => A_shifted(33), A2 => n179, B1 => 
                           zeroSignal(33), B2 => n170, C1 => A_neg_shifted(33),
                           C2 => n163, ZN => n239);
   U153 : NAND2_X1 port map( A1 => n248, A2 => n247, ZN => Y(37));
   U154 : AOI222_X1 port map( A1 => A_shifted(37), A2 => n179, B1 => 
                           zeroSignal(37), B2 => n170, C1 => A_neg_shifted(37),
                           C2 => n162, ZN => n247);
   U155 : AOI22_X1 port map( A1 => A_neg(37), A2 => n153, B1 => A_signal(37), 
                           B2 => n144, ZN => n248);
   U156 : NAND2_X1 port map( A1 => n242, A2 => n241, ZN => Y(34));
   U157 : AOI222_X1 port map( A1 => A_shifted(34), A2 => n179, B1 => 
                           zeroSignal(34), B2 => n170, C1 => A_neg_shifted(34),
                           C2 => n163, ZN => n241);
   U158 : NAND2_X1 port map( A1 => n188, A2 => n187, ZN => Y(0));
   U159 : AOI22_X1 port map( A1 => A_neg(0), A2 => n151, B1 => A_signal(0), B2 
                           => n142, ZN => n188);
   U160 : AOI222_X1 port map( A1 => A_shifted(0), A2 => n177, B1 => 
                           zeroSignal(0), B2 => n168, C1 => A_neg_shifted(0), 
                           C2 => n165, ZN => n187);
   U161 : NAND2_X1 port map( A1 => n210, A2 => n209, ZN => Y(1));
   U162 : AOI22_X1 port map( A1 => A_neg(1), A2 => n151, B1 => A_signal(1), B2 
                           => n142, ZN => n210);
   U163 : AOI222_X1 port map( A1 => A_shifted(1), A2 => n178, B1 => 
                           zeroSignal(1), B2 => n168, C1 => A_neg_shifted(1), 
                           C2 => n164, ZN => n209);
   U164 : NAND2_X1 port map( A1 => n232, A2 => n231, ZN => Y(2));
   U165 : AOI22_X1 port map( A1 => A_neg(2), A2 => n152, B1 => A_signal(2), B2 
                           => n143, ZN => n232);
   U166 : AOI222_X1 port map( A1 => A_shifted(2), A2 => n179, B1 => 
                           zeroSignal(2), B2 => n169, C1 => A_neg_shifted(2), 
                           C2 => n163, ZN => n231);
   U167 : NAND2_X1 port map( A1 => n254, A2 => n253, ZN => Y(3));
   U168 : AOI22_X1 port map( A1 => A_neg(3), A2 => n153, B1 => A_signal(3), B2 
                           => n144, ZN => n254);
   U169 : AOI222_X1 port map( A1 => A_shifted(3), A2 => n180, B1 => 
                           zeroSignal(3), B2 => n170, C1 => A_neg_shifted(3), 
                           C2 => n162, ZN => n253);
   U170 : NAND2_X1 port map( A1 => n276, A2 => n275, ZN => Y(4));
   U171 : AOI22_X1 port map( A1 => A_neg(4), A2 => n154, B1 => A_signal(4), B2 
                           => n145, ZN => n276);
   U172 : AOI222_X1 port map( A1 => A_shifted(4), A2 => n181, B1 => 
                           zeroSignal(4), B2 => n171, C1 => A_neg_shifted(4), 
                           C2 => n161, ZN => n275);
   U173 : NAND2_X1 port map( A1 => n298, A2 => n297, ZN => Y(5));
   U174 : AOI22_X1 port map( A1 => A_neg(5), A2 => n155, B1 => A_signal(5), B2 
                           => n146, ZN => n298);
   U175 : AOI222_X1 port map( A1 => A_shifted(5), A2 => n182, B1 => 
                           zeroSignal(5), B2 => n172, C1 => A_neg_shifted(5), 
                           C2 => n160, ZN => n297);
   U176 : NAND2_X1 port map( A1 => n308, A2 => n307, ZN => Y(6));
   U177 : AOI22_X1 port map( A1 => A_neg(6), A2 => n156, B1 => A_signal(6), B2 
                           => n147, ZN => n308);
   U178 : AOI222_X1 port map( A1 => A_shifted(6), A2 => n182, B1 => 
                           zeroSignal(6), B2 => n173, C1 => A_neg_shifted(6), 
                           C2 => n160, ZN => n307);
   U179 : NAND2_X1 port map( A1 => n310, A2 => n309, ZN => Y(7));
   U180 : AOI22_X1 port map( A1 => A_neg(7), A2 => n156, B1 => A_signal(7), B2 
                           => n147, ZN => n310);
   U181 : AOI222_X1 port map( A1 => A_shifted(7), A2 => n182, B1 => 
                           zeroSignal(7), B2 => n173, C1 => A_neg_shifted(7), 
                           C2 => n160, ZN => n309);
   U182 : NAND2_X1 port map( A1 => n312, A2 => n311, ZN => Y(8));
   U183 : AOI22_X1 port map( A1 => A_neg(8), A2 => n156, B1 => A_signal(8), B2 
                           => n147, ZN => n312);
   U184 : AOI222_X1 port map( A1 => A_shifted(8), A2 => n182, B1 => 
                           zeroSignal(8), B2 => n173, C1 => A_neg_shifted(8), 
                           C2 => n160, ZN => n311);
   U185 : NAND2_X1 port map( A1 => n318, A2 => n317, ZN => Y(9));
   U186 : AOI22_X1 port map( A1 => A_neg(9), A2 => n156, B1 => A_signal(9), B2 
                           => n147, ZN => n318);
   U187 : AOI222_X1 port map( A1 => A_shifted(9), A2 => n182, B1 => 
                           zeroSignal(9), B2 => n173, C1 => A_neg_shifted(9), 
                           C2 => n160, ZN => n317);
   U188 : NAND2_X1 port map( A1 => n190, A2 => n189, ZN => Y(10));
   U189 : AOI22_X1 port map( A1 => A_neg(10), A2 => n151, B1 => A_signal(10), 
                           B2 => n142, ZN => n190);
   U190 : AOI222_X1 port map( A1 => A_shifted(10), A2 => n177, B1 => 
                           zeroSignal(10), B2 => n168, C1 => A_neg_shifted(10),
                           C2 => n165, ZN => n189);
   U191 : NAND2_X1 port map( A1 => n192, A2 => n191, ZN => Y(11));
   U192 : AOI22_X1 port map( A1 => A_neg(11), A2 => n151, B1 => A_signal(11), 
                           B2 => n142, ZN => n192);
   U193 : AOI222_X1 port map( A1 => A_shifted(11), A2 => n177, B1 => 
                           zeroSignal(11), B2 => n168, C1 => A_neg_shifted(11),
                           C2 => n165, ZN => n191);
   U194 : NAND2_X1 port map( A1 => n194, A2 => n193, ZN => Y(12));
   U195 : AOI22_X1 port map( A1 => A_neg(12), A2 => n151, B1 => A_signal(12), 
                           B2 => n142, ZN => n194);
   U196 : AOI222_X1 port map( A1 => A_shifted(12), A2 => n177, B1 => 
                           zeroSignal(12), B2 => n168, C1 => A_neg_shifted(12),
                           C2 => n165, ZN => n193);
   U197 : NAND2_X1 port map( A1 => n196, A2 => n195, ZN => Y(13));
   U198 : AOI22_X1 port map( A1 => A_neg(13), A2 => n151, B1 => A_signal(13), 
                           B2 => n142, ZN => n196);
   U199 : AOI222_X1 port map( A1 => A_shifted(13), A2 => n177, B1 => 
                           zeroSignal(13), B2 => n168, C1 => A_neg_shifted(13),
                           C2 => n164, ZN => n195);
   U200 : NAND2_X1 port map( A1 => n198, A2 => n197, ZN => Y(14));
   U201 : AOI22_X1 port map( A1 => A_neg(14), A2 => n151, B1 => A_signal(14), 
                           B2 => n142, ZN => n198);
   U202 : AOI222_X1 port map( A1 => A_shifted(14), A2 => n177, B1 => 
                           zeroSignal(14), B2 => n168, C1 => A_neg_shifted(14),
                           C2 => n164, ZN => n197);
   U203 : NAND2_X1 port map( A1 => n200, A2 => n199, ZN => Y(15));
   U204 : AOI22_X1 port map( A1 => A_neg(15), A2 => n151, B1 => A_signal(15), 
                           B2 => n142, ZN => n200);
   U205 : AOI222_X1 port map( A1 => A_shifted(15), A2 => n177, B1 => 
                           zeroSignal(15), B2 => n168, C1 => A_neg_shifted(15),
                           C2 => n164, ZN => n199);
   U206 : NAND2_X1 port map( A1 => n202, A2 => n201, ZN => Y(16));
   U207 : AOI22_X1 port map( A1 => A_neg(16), A2 => n151, B1 => A_signal(16), 
                           B2 => n142, ZN => n202);
   U208 : AOI222_X1 port map( A1 => A_shifted(16), A2 => n177, B1 => 
                           zeroSignal(16), B2 => n168, C1 => A_neg_shifted(16),
                           C2 => n164, ZN => n201);
   U209 : NAND2_X1 port map( A1 => n204, A2 => n203, ZN => Y(17));
   U210 : AOI22_X1 port map( A1 => A_neg(17), A2 => n151, B1 => A_signal(17), 
                           B2 => n142, ZN => n204);
   U211 : AOI222_X1 port map( A1 => A_shifted(17), A2 => n177, B1 => 
                           zeroSignal(17), B2 => n168, C1 => A_neg_shifted(17),
                           C2 => n164, ZN => n203);
   U212 : NAND2_X1 port map( A1 => n206, A2 => n205, ZN => Y(18));
   U213 : AOI22_X1 port map( A1 => A_neg(18), A2 => n151, B1 => A_signal(18), 
                           B2 => n142, ZN => n206);
   U214 : AOI222_X1 port map( A1 => A_shifted(18), A2 => n177, B1 => 
                           zeroSignal(18), B2 => n168, C1 => A_neg_shifted(18),
                           C2 => n164, ZN => n205);
   U215 : NAND2_X1 port map( A1 => n208, A2 => n207, ZN => Y(19));
   U216 : AOI22_X1 port map( A1 => A_neg(19), A2 => n151, B1 => A_signal(19), 
                           B2 => n142, ZN => n208);
   U217 : AOI222_X1 port map( A1 => A_shifted(19), A2 => n177, B1 => 
                           zeroSignal(19), B2 => n168, C1 => A_neg_shifted(19),
                           C2 => n164, ZN => n207);
   U218 : NAND2_X1 port map( A1 => n212, A2 => n211, ZN => Y(20));
   U219 : AOI22_X1 port map( A1 => A_neg(20), A2 => n152, B1 => A_signal(20), 
                           B2 => n143, ZN => n212);
   U220 : AOI222_X1 port map( A1 => A_shifted(20), A2 => n178, B1 => 
                           zeroSignal(20), B2 => n169, C1 => A_neg_shifted(20),
                           C2 => n164, ZN => n211);
   U221 : NAND2_X1 port map( A1 => n214, A2 => n213, ZN => Y(21));
   U222 : AOI22_X1 port map( A1 => A_neg(21), A2 => n152, B1 => A_signal(21), 
                           B2 => n143, ZN => n214);
   U223 : AOI222_X1 port map( A1 => A_shifted(21), A2 => n178, B1 => 
                           zeroSignal(21), B2 => n169, C1 => A_neg_shifted(21),
                           C2 => n164, ZN => n213);
   U224 : NAND2_X1 port map( A1 => n216, A2 => n215, ZN => Y(22));
   U225 : AOI22_X1 port map( A1 => A_neg(22), A2 => n152, B1 => A_signal(22), 
                           B2 => n143, ZN => n216);
   U226 : AOI222_X1 port map( A1 => A_shifted(22), A2 => n178, B1 => 
                           zeroSignal(22), B2 => n169, C1 => A_neg_shifted(22),
                           C2 => n164, ZN => n215);
   U227 : NAND2_X1 port map( A1 => n218, A2 => n217, ZN => Y(23));
   U228 : AOI22_X1 port map( A1 => A_neg(23), A2 => n152, B1 => A_signal(23), 
                           B2 => n143, ZN => n218);
   U229 : AOI222_X1 port map( A1 => A_shifted(23), A2 => n178, B1 => 
                           zeroSignal(23), B2 => n169, C1 => A_neg_shifted(23),
                           C2 => n164, ZN => n217);
   U230 : NAND2_X1 port map( A1 => n220, A2 => n219, ZN => Y(24));
   U231 : AOI22_X1 port map( A1 => A_neg(24), A2 => n152, B1 => A_signal(24), 
                           B2 => n143, ZN => n220);
   U232 : AOI222_X1 port map( A1 => A_shifted(24), A2 => n178, B1 => 
                           zeroSignal(24), B2 => n169, C1 => A_neg_shifted(24),
                           C2 => n163, ZN => n219);
   U233 : NAND2_X1 port map( A1 => n222, A2 => n221, ZN => Y(25));
   U234 : AOI22_X1 port map( A1 => A_neg(25), A2 => n152, B1 => A_signal(25), 
                           B2 => n143, ZN => n222);
   U235 : AOI222_X1 port map( A1 => A_shifted(25), A2 => n178, B1 => 
                           zeroSignal(25), B2 => n169, C1 => A_neg_shifted(25),
                           C2 => n163, ZN => n221);
   U236 : NAND2_X1 port map( A1 => n224, A2 => n223, ZN => Y(26));
   U237 : AOI22_X1 port map( A1 => A_neg(26), A2 => n152, B1 => A_signal(26), 
                           B2 => n143, ZN => n224);
   U238 : AOI222_X1 port map( A1 => A_shifted(26), A2 => n178, B1 => 
                           zeroSignal(26), B2 => n169, C1 => A_neg_shifted(26),
                           C2 => n163, ZN => n223);
   U239 : NAND2_X1 port map( A1 => n226, A2 => n225, ZN => Y(27));
   U240 : AOI22_X1 port map( A1 => A_neg(27), A2 => n152, B1 => A_signal(27), 
                           B2 => n143, ZN => n226);
   U241 : AOI222_X1 port map( A1 => A_shifted(27), A2 => n178, B1 => 
                           zeroSignal(27), B2 => n169, C1 => A_neg_shifted(27),
                           C2 => n163, ZN => n225);
   U242 : AOI22_X1 port map( A1 => A_neg(34), A2 => n153, B1 => A_signal(34), 
                           B2 => n144, ZN => n242);
   U243 : AOI22_X1 port map( A1 => A_neg(33), A2 => n153, B1 => A_signal(33), 
                           B2 => n144, ZN => n240);
   U244 : AOI22_X1 port map( A1 => A_neg(31), A2 => n153, B1 => A_signal(31), 
                           B2 => n144, ZN => n236);

end SYN_BEHAVIORAL_2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity MUX51_MuxNbit64_1 is

   port( zeroSignal, A_signal, A_neg, A_shifted, A_neg_shifted : in 
         std_logic_vector (63 downto 0);  Sel : in std_logic_vector (2 downto 
         0);  Y : out std_logic_vector (63 downto 0));

end MUX51_MuxNbit64_1;

architecture SYN_BEHAVIORAL_2 of MUX51_MuxNbit64_1 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, 
      n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, 
      n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, 
      n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, 
      n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, 
      n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, 
      n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, 
      n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, 
      n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, 
      n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, 
      n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, 
      n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, 
      n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, 
      n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, 
      n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, 
      n320 : std_logic;

begin
   
   U1 : AND3_X1 port map( A1 => n319, A2 => n320, A3 => Sel(2), ZN => n141);
   U2 : BUF_X1 port map( A => n141, Z => n166);
   U3 : BUF_X1 port map( A => n159, Z => n158);
   U4 : BUF_X1 port map( A => n185, Z => n184);
   U5 : BUF_X1 port map( A => n150, Z => n149);
   U6 : BUF_X1 port map( A => n141, Z => n167);
   U7 : BUF_X1 port map( A => n185, Z => n183);
   U8 : BUF_X1 port map( A => n159, Z => n157);
   U9 : BUF_X1 port map( A => n150, Z => n148);
   U10 : BUF_X1 port map( A => n176, Z => n175);
   U11 : BUF_X1 port map( A => n176, Z => n174);
   U12 : BUF_X1 port map( A => n184, Z => n179);
   U13 : BUF_X1 port map( A => n158, Z => n153);
   U14 : BUF_X1 port map( A => n149, Z => n144);
   U15 : BUF_X1 port map( A => n166, Z => n163);
   U16 : BUF_X1 port map( A => n149, Z => n143);
   U17 : BUF_X1 port map( A => n158, Z => n152);
   U18 : BUF_X1 port map( A => n167, Z => n162);
   U19 : BUF_X1 port map( A => n183, Z => n180);
   U20 : BUF_X1 port map( A => n157, Z => n154);
   U21 : BUF_X1 port map( A => n148, Z => n145);
   U22 : BUF_X1 port map( A => n167, Z => n161);
   U23 : BUF_X1 port map( A => n183, Z => n181);
   U24 : BUF_X1 port map( A => n157, Z => n155);
   U25 : BUF_X1 port map( A => n148, Z => n146);
   U26 : BUF_X1 port map( A => n167, Z => n160);
   U27 : BUF_X1 port map( A => n183, Z => n182);
   U28 : BUF_X1 port map( A => n158, Z => n151);
   U29 : BUF_X1 port map( A => n149, Z => n142);
   U30 : BUF_X1 port map( A => n175, Z => n168);
   U31 : BUF_X1 port map( A => n175, Z => n169);
   U32 : BUF_X1 port map( A => n175, Z => n170);
   U33 : BUF_X1 port map( A => n174, Z => n171);
   U34 : BUF_X1 port map( A => n174, Z => n172);
   U35 : BUF_X1 port map( A => n166, Z => n164);
   U36 : BUF_X1 port map( A => n184, Z => n177);
   U37 : BUF_X1 port map( A => n184, Z => n178);
   U38 : BUF_X1 port map( A => n166, Z => n165);
   U39 : BUF_X1 port map( A => n157, Z => n156);
   U40 : BUF_X1 port map( A => n148, Z => n147);
   U41 : BUF_X1 port map( A => n174, Z => n173);
   U42 : INV_X1 port map( A => Sel(1), ZN => n320);
   U43 : BUF_X1 port map( A => n316, Z => n185);
   U44 : NOR3_X1 port map( A1 => n319, A2 => Sel(2), A3 => n320, ZN => n316);
   U45 : BUF_X1 port map( A => n314, Z => n159);
   U46 : NOR3_X1 port map( A1 => Sel(0), A2 => Sel(2), A3 => n320, ZN => n314);
   U47 : INV_X1 port map( A => Sel(0), ZN => n319);
   U48 : BUF_X1 port map( A => n313, Z => n150);
   U49 : NOR3_X1 port map( A1 => Sel(1), A2 => Sel(2), A3 => n319, ZN => n313);
   U50 : BUF_X1 port map( A => n315, Z => n176);
   U51 : NOR2_X1 port map( A1 => n165, A2 => n186, ZN => n315);
   U52 : AOI21_X1 port map( B1 => n319, B2 => n320, A => Sel(2), ZN => n186);
   U53 : NAND2_X1 port map( A1 => n236, A2 => n235, ZN => Y(31));
   U54 : AOI22_X1 port map( A1 => A_neg(31), A2 => n153, B1 => A_signal(31), B2
                           => n144, ZN => n236);
   U55 : AOI222_X1 port map( A1 => A_shifted(31), A2 => n179, B1 => 
                           zeroSignal(31), B2 => n170, C1 => A_neg_shifted(31),
                           C2 => n163, ZN => n235);
   U56 : NAND2_X1 port map( A1 => n238, A2 => n237, ZN => Y(32));
   U57 : AOI22_X1 port map( A1 => A_neg(32), A2 => n153, B1 => A_signal(32), B2
                           => n144, ZN => n238);
   U58 : AOI222_X1 port map( A1 => A_shifted(32), A2 => n179, B1 => 
                           zeroSignal(32), B2 => n170, C1 => A_neg_shifted(32),
                           C2 => n163, ZN => n237);
   U59 : NAND2_X1 port map( A1 => n266, A2 => n265, ZN => Y(45));
   U60 : AOI222_X1 port map( A1 => A_shifted(45), A2 => n180, B1 => 
                           zeroSignal(45), B2 => n171, C1 => A_neg_shifted(45),
                           C2 => n162, ZN => n265);
   U61 : AOI22_X1 port map( A1 => A_neg(45), A2 => n154, B1 => A_signal(45), B2
                           => n145, ZN => n266);
   U62 : NAND2_X1 port map( A1 => n262, A2 => n261, ZN => Y(43));
   U63 : AOI222_X1 port map( A1 => A_shifted(43), A2 => n180, B1 => 
                           zeroSignal(43), B2 => n171, C1 => A_neg_shifted(43),
                           C2 => n162, ZN => n261);
   U64 : AOI22_X1 port map( A1 => A_neg(43), A2 => n154, B1 => A_signal(43), B2
                           => n145, ZN => n262);
   U65 : NAND2_X1 port map( A1 => n264, A2 => n263, ZN => Y(44));
   U66 : AOI222_X1 port map( A1 => A_shifted(44), A2 => n180, B1 => 
                           zeroSignal(44), B2 => n171, C1 => A_neg_shifted(44),
                           C2 => n162, ZN => n263);
   U67 : AOI22_X1 port map( A1 => A_neg(44), A2 => n154, B1 => A_signal(44), B2
                           => n145, ZN => n264);
   U68 : NAND2_X1 port map( A1 => n268, A2 => n267, ZN => Y(46));
   U69 : AOI222_X1 port map( A1 => A_shifted(46), A2 => n180, B1 => 
                           zeroSignal(46), B2 => n171, C1 => A_neg_shifted(46),
                           C2 => n161, ZN => n267);
   U70 : AOI22_X1 port map( A1 => A_neg(46), A2 => n154, B1 => A_signal(46), B2
                           => n145, ZN => n268);
   U71 : NAND2_X1 port map( A1 => n234, A2 => n233, ZN => Y(30));
   U72 : AOI222_X1 port map( A1 => A_shifted(30), A2 => n179, B1 => 
                           zeroSignal(30), B2 => n169, C1 => A_neg_shifted(30),
                           C2 => n163, ZN => n233);
   U73 : AOI22_X1 port map( A1 => A_neg(30), A2 => n152, B1 => A_signal(30), B2
                           => n143, ZN => n234);
   U74 : NAND2_X1 port map( A1 => n270, A2 => n269, ZN => Y(47));
   U75 : AOI222_X1 port map( A1 => A_shifted(47), A2 => n180, B1 => 
                           zeroSignal(47), B2 => n171, C1 => A_neg_shifted(47),
                           C2 => n161, ZN => n269);
   U76 : AOI22_X1 port map( A1 => A_neg(47), A2 => n154, B1 => A_signal(47), B2
                           => n145, ZN => n270);
   U77 : NAND2_X1 port map( A1 => n274, A2 => n273, ZN => Y(49));
   U78 : AOI222_X1 port map( A1 => A_shifted(49), A2 => n180, B1 => 
                           zeroSignal(49), B2 => n171, C1 => A_neg_shifted(49),
                           C2 => n161, ZN => n273);
   U79 : AOI22_X1 port map( A1 => A_neg(49), A2 => n154, B1 => A_signal(49), B2
                           => n145, ZN => n274);
   U80 : NAND2_X1 port map( A1 => n278, A2 => n277, ZN => Y(50));
   U81 : AOI222_X1 port map( A1 => A_shifted(50), A2 => n181, B1 => 
                           zeroSignal(50), B2 => n171, C1 => A_neg_shifted(50),
                           C2 => n161, ZN => n277);
   U82 : AOI22_X1 port map( A1 => A_neg(50), A2 => n154, B1 => A_signal(50), B2
                           => n145, ZN => n278);
   U83 : NAND2_X1 port map( A1 => n280, A2 => n279, ZN => Y(51));
   U84 : AOI222_X1 port map( A1 => A_shifted(51), A2 => n181, B1 => 
                           zeroSignal(51), B2 => n171, C1 => A_neg_shifted(51),
                           C2 => n161, ZN => n279);
   U85 : AOI22_X1 port map( A1 => A_neg(51), A2 => n154, B1 => A_signal(51), B2
                           => n145, ZN => n280);
   U86 : NAND2_X1 port map( A1 => n282, A2 => n281, ZN => Y(52));
   U87 : AOI222_X1 port map( A1 => A_shifted(52), A2 => n181, B1 => 
                           zeroSignal(52), B2 => n171, C1 => A_neg_shifted(52),
                           C2 => n161, ZN => n281);
   U88 : AOI22_X1 port map( A1 => A_neg(52), A2 => n154, B1 => A_signal(52), B2
                           => n145, ZN => n282);
   U89 : NAND2_X1 port map( A1 => n284, A2 => n283, ZN => Y(53));
   U90 : AOI222_X1 port map( A1 => A_shifted(53), A2 => n181, B1 => 
                           zeroSignal(53), B2 => n172, C1 => A_neg_shifted(53),
                           C2 => n161, ZN => n283);
   U91 : AOI22_X1 port map( A1 => A_neg(53), A2 => n155, B1 => A_signal(53), B2
                           => n146, ZN => n284);
   U92 : NAND2_X1 port map( A1 => n286, A2 => n285, ZN => Y(54));
   U93 : AOI222_X1 port map( A1 => A_shifted(54), A2 => n181, B1 => 
                           zeroSignal(54), B2 => n172, C1 => A_neg_shifted(54),
                           C2 => n161, ZN => n285);
   U94 : AOI22_X1 port map( A1 => A_neg(54), A2 => n155, B1 => A_signal(54), B2
                           => n146, ZN => n286);
   U95 : NAND2_X1 port map( A1 => n288, A2 => n287, ZN => Y(55));
   U96 : AOI222_X1 port map( A1 => A_shifted(55), A2 => n181, B1 => 
                           zeroSignal(55), B2 => n172, C1 => A_neg_shifted(55),
                           C2 => n161, ZN => n287);
   U97 : AOI22_X1 port map( A1 => A_neg(55), A2 => n155, B1 => A_signal(55), B2
                           => n146, ZN => n288);
   U98 : NAND2_X1 port map( A1 => n290, A2 => n289, ZN => Y(56));
   U99 : AOI222_X1 port map( A1 => A_shifted(56), A2 => n181, B1 => 
                           zeroSignal(56), B2 => n172, C1 => A_neg_shifted(56),
                           C2 => n161, ZN => n289);
   U100 : AOI22_X1 port map( A1 => A_neg(56), A2 => n155, B1 => A_signal(56), 
                           B2 => n146, ZN => n290);
   U101 : NAND2_X1 port map( A1 => n240, A2 => n239, ZN => Y(33));
   U102 : AOI222_X1 port map( A1 => A_shifted(33), A2 => n179, B1 => 
                           zeroSignal(33), B2 => n170, C1 => A_neg_shifted(33),
                           C2 => n163, ZN => n239);
   U103 : NAND2_X1 port map( A1 => n292, A2 => n291, ZN => Y(57));
   U104 : AOI222_X1 port map( A1 => A_shifted(57), A2 => n181, B1 => 
                           zeroSignal(57), B2 => n172, C1 => A_neg_shifted(57),
                           C2 => n160, ZN => n291);
   U105 : AOI22_X1 port map( A1 => A_neg(57), A2 => n155, B1 => A_signal(57), 
                           B2 => n146, ZN => n292);
   U106 : NAND2_X1 port map( A1 => n304, A2 => n303, ZN => Y(62));
   U107 : AOI222_X1 port map( A1 => A_shifted(62), A2 => n182, B1 => 
                           zeroSignal(62), B2 => n172, C1 => A_neg_shifted(62),
                           C2 => n160, ZN => n303);
   U108 : AOI22_X1 port map( A1 => A_neg(62), A2 => n155, B1 => A_signal(62), 
                           B2 => n146, ZN => n304);
   U109 : NAND2_X1 port map( A1 => n294, A2 => n293, ZN => Y(58));
   U110 : AOI222_X1 port map( A1 => A_shifted(58), A2 => n181, B1 => 
                           zeroSignal(58), B2 => n172, C1 => A_neg_shifted(58),
                           C2 => n160, ZN => n293);
   U111 : AOI22_X1 port map( A1 => A_neg(58), A2 => n155, B1 => A_signal(58), 
                           B2 => n146, ZN => n294);
   U112 : NAND2_X1 port map( A1 => n272, A2 => n271, ZN => Y(48));
   U113 : AOI22_X1 port map( A1 => A_neg(48), A2 => n154, B1 => A_signal(48), 
                           B2 => n145, ZN => n272);
   U114 : AOI222_X1 port map( A1 => A_shifted(48), A2 => n180, B1 => 
                           zeroSignal(48), B2 => n171, C1 => A_neg_shifted(48),
                           C2 => n161, ZN => n271);
   U115 : NAND2_X1 port map( A1 => n302, A2 => n301, ZN => Y(61));
   U116 : AOI222_X1 port map( A1 => A_shifted(61), A2 => n182, B1 => 
                           zeroSignal(61), B2 => n172, C1 => A_neg_shifted(61),
                           C2 => n160, ZN => n301);
   U117 : AOI22_X1 port map( A1 => A_neg(61), A2 => n155, B1 => A_signal(61), 
                           B2 => n146, ZN => n302);
   U118 : NAND2_X1 port map( A1 => n300, A2 => n299, ZN => Y(60));
   U119 : AOI222_X1 port map( A1 => A_shifted(60), A2 => n182, B1 => 
                           zeroSignal(60), B2 => n172, C1 => A_neg_shifted(60),
                           C2 => n160, ZN => n299);
   U120 : AOI22_X1 port map( A1 => A_neg(60), A2 => n155, B1 => A_signal(60), 
                           B2 => n146, ZN => n300);
   U121 : NAND2_X1 port map( A1 => n306, A2 => n305, ZN => Y(63));
   U122 : AOI222_X1 port map( A1 => A_shifted(63), A2 => n182, B1 => 
                           zeroSignal(63), B2 => n172, C1 => A_neg_shifted(63),
                           C2 => n160, ZN => n305);
   U123 : AOI22_X1 port map( A1 => A_neg(63), A2 => n155, B1 => A_signal(63), 
                           B2 => n146, ZN => n306);
   U124 : NAND2_X1 port map( A1 => n256, A2 => n255, ZN => Y(40));
   U125 : AOI222_X1 port map( A1 => A_shifted(40), A2 => n180, B1 => 
                           zeroSignal(40), B2 => n170, C1 => A_neg_shifted(40),
                           C2 => n162, ZN => n255);
   U126 : AOI22_X1 port map( A1 => A_neg(40), A2 => n153, B1 => A_signal(40), 
                           B2 => n144, ZN => n256);
   U127 : NAND2_X1 port map( A1 => n296, A2 => n295, ZN => Y(59));
   U128 : AOI22_X1 port map( A1 => A_neg(59), A2 => n155, B1 => A_signal(59), 
                           B2 => n146, ZN => n296);
   U129 : AOI222_X1 port map( A1 => A_shifted(59), A2 => n181, B1 => 
                           zeroSignal(59), B2 => n172, C1 => A_neg_shifted(59),
                           C2 => n160, ZN => n295);
   U130 : NAND2_X1 port map( A1 => n260, A2 => n259, ZN => Y(42));
   U131 : AOI222_X1 port map( A1 => A_shifted(42), A2 => n180, B1 => 
                           zeroSignal(42), B2 => n171, C1 => A_neg_shifted(42),
                           C2 => n162, ZN => n259);
   U132 : AOI22_X1 port map( A1 => A_neg(42), A2 => n154, B1 => A_signal(42), 
                           B2 => n145, ZN => n260);
   U133 : NAND2_X1 port map( A1 => n242, A2 => n241, ZN => Y(34));
   U134 : AOI22_X1 port map( A1 => A_neg(34), A2 => n153, B1 => A_signal(34), 
                           B2 => n144, ZN => n242);
   U135 : AOI222_X1 port map( A1 => A_shifted(34), A2 => n179, B1 => 
                           zeroSignal(34), B2 => n170, C1 => A_neg_shifted(34),
                           C2 => n163, ZN => n241);
   U136 : NAND2_X1 port map( A1 => n258, A2 => n257, ZN => Y(41));
   U137 : AOI22_X1 port map( A1 => A_neg(41), A2 => n153, B1 => A_signal(41), 
                           B2 => n144, ZN => n258);
   U138 : AOI222_X1 port map( A1 => A_shifted(41), A2 => n180, B1 => 
                           zeroSignal(41), B2 => n170, C1 => A_neg_shifted(41),
                           C2 => n162, ZN => n257);
   U139 : NAND2_X1 port map( A1 => n244, A2 => n243, ZN => Y(35));
   U140 : AOI222_X1 port map( A1 => A_shifted(35), A2 => n179, B1 => 
                           zeroSignal(35), B2 => n170, C1 => A_neg_shifted(35),
                           C2 => n162, ZN => n243);
   U141 : NAND2_X1 port map( A1 => n248, A2 => n247, ZN => Y(37));
   U142 : AOI222_X1 port map( A1 => A_shifted(37), A2 => n179, B1 => 
                           zeroSignal(37), B2 => n170, C1 => A_neg_shifted(37),
                           C2 => n162, ZN => n247);
   U143 : AOI22_X1 port map( A1 => A_neg(37), A2 => n153, B1 => A_signal(37), 
                           B2 => n144, ZN => n248);
   U144 : NAND2_X1 port map( A1 => n250, A2 => n249, ZN => Y(38));
   U145 : AOI222_X1 port map( A1 => A_shifted(38), A2 => n179, B1 => 
                           zeroSignal(38), B2 => n170, C1 => A_neg_shifted(38),
                           C2 => n162, ZN => n249);
   U146 : AOI22_X1 port map( A1 => A_neg(38), A2 => n153, B1 => A_signal(38), 
                           B2 => n144, ZN => n250);
   U147 : NAND2_X1 port map( A1 => n252, A2 => n251, ZN => Y(39));
   U148 : AOI222_X1 port map( A1 => A_shifted(39), A2 => n179, B1 => 
                           zeroSignal(39), B2 => n170, C1 => A_neg_shifted(39),
                           C2 => n162, ZN => n251);
   U149 : AOI22_X1 port map( A1 => A_neg(39), A2 => n153, B1 => A_signal(39), 
                           B2 => n144, ZN => n252);
   U150 : NAND2_X1 port map( A1 => n246, A2 => n245, ZN => Y(36));
   U151 : AOI222_X1 port map( A1 => A_shifted(36), A2 => n179, B1 => 
                           zeroSignal(36), B2 => n170, C1 => A_neg_shifted(36),
                           C2 => n162, ZN => n245);
   U152 : NAND2_X1 port map( A1 => n188, A2 => n187, ZN => Y(0));
   U153 : AOI22_X1 port map( A1 => A_neg(0), A2 => n151, B1 => A_signal(0), B2 
                           => n142, ZN => n188);
   U154 : AOI222_X1 port map( A1 => A_shifted(0), A2 => n177, B1 => 
                           zeroSignal(0), B2 => n168, C1 => A_neg_shifted(0), 
                           C2 => n165, ZN => n187);
   U155 : NAND2_X1 port map( A1 => n210, A2 => n209, ZN => Y(1));
   U156 : AOI22_X1 port map( A1 => A_neg(1), A2 => n151, B1 => A_signal(1), B2 
                           => n142, ZN => n210);
   U157 : AOI222_X1 port map( A1 => A_shifted(1), A2 => n178, B1 => 
                           zeroSignal(1), B2 => n168, C1 => A_neg_shifted(1), 
                           C2 => n164, ZN => n209);
   U158 : NAND2_X1 port map( A1 => n232, A2 => n231, ZN => Y(2));
   U159 : AOI22_X1 port map( A1 => A_neg(2), A2 => n152, B1 => A_signal(2), B2 
                           => n143, ZN => n232);
   U160 : AOI222_X1 port map( A1 => A_shifted(2), A2 => n179, B1 => 
                           zeroSignal(2), B2 => n169, C1 => A_neg_shifted(2), 
                           C2 => n163, ZN => n231);
   U161 : NAND2_X1 port map( A1 => n254, A2 => n253, ZN => Y(3));
   U162 : AOI22_X1 port map( A1 => A_neg(3), A2 => n153, B1 => A_signal(3), B2 
                           => n144, ZN => n254);
   U163 : AOI222_X1 port map( A1 => A_shifted(3), A2 => n180, B1 => 
                           zeroSignal(3), B2 => n170, C1 => A_neg_shifted(3), 
                           C2 => n162, ZN => n253);
   U164 : NAND2_X1 port map( A1 => n276, A2 => n275, ZN => Y(4));
   U165 : AOI22_X1 port map( A1 => A_neg(4), A2 => n154, B1 => A_signal(4), B2 
                           => n145, ZN => n276);
   U166 : AOI222_X1 port map( A1 => A_shifted(4), A2 => n181, B1 => 
                           zeroSignal(4), B2 => n171, C1 => A_neg_shifted(4), 
                           C2 => n161, ZN => n275);
   U167 : NAND2_X1 port map( A1 => n298, A2 => n297, ZN => Y(5));
   U168 : AOI22_X1 port map( A1 => A_neg(5), A2 => n155, B1 => A_signal(5), B2 
                           => n146, ZN => n298);
   U169 : AOI222_X1 port map( A1 => A_shifted(5), A2 => n182, B1 => 
                           zeroSignal(5), B2 => n172, C1 => A_neg_shifted(5), 
                           C2 => n160, ZN => n297);
   U170 : NAND2_X1 port map( A1 => n308, A2 => n307, ZN => Y(6));
   U171 : AOI22_X1 port map( A1 => A_neg(6), A2 => n156, B1 => A_signal(6), B2 
                           => n147, ZN => n308);
   U172 : AOI222_X1 port map( A1 => A_shifted(6), A2 => n182, B1 => 
                           zeroSignal(6), B2 => n173, C1 => A_neg_shifted(6), 
                           C2 => n160, ZN => n307);
   U173 : NAND2_X1 port map( A1 => n310, A2 => n309, ZN => Y(7));
   U174 : AOI22_X1 port map( A1 => A_neg(7), A2 => n156, B1 => A_signal(7), B2 
                           => n147, ZN => n310);
   U175 : AOI222_X1 port map( A1 => A_shifted(7), A2 => n182, B1 => 
                           zeroSignal(7), B2 => n173, C1 => A_neg_shifted(7), 
                           C2 => n160, ZN => n309);
   U176 : NAND2_X1 port map( A1 => n312, A2 => n311, ZN => Y(8));
   U177 : AOI22_X1 port map( A1 => A_neg(8), A2 => n156, B1 => A_signal(8), B2 
                           => n147, ZN => n312);
   U178 : AOI222_X1 port map( A1 => A_shifted(8), A2 => n182, B1 => 
                           zeroSignal(8), B2 => n173, C1 => A_neg_shifted(8), 
                           C2 => n160, ZN => n311);
   U179 : NAND2_X1 port map( A1 => n318, A2 => n317, ZN => Y(9));
   U180 : AOI22_X1 port map( A1 => A_neg(9), A2 => n156, B1 => A_signal(9), B2 
                           => n147, ZN => n318);
   U181 : AOI222_X1 port map( A1 => A_shifted(9), A2 => n182, B1 => 
                           zeroSignal(9), B2 => n173, C1 => A_neg_shifted(9), 
                           C2 => n160, ZN => n317);
   U182 : NAND2_X1 port map( A1 => n190, A2 => n189, ZN => Y(10));
   U183 : AOI22_X1 port map( A1 => A_neg(10), A2 => n151, B1 => A_signal(10), 
                           B2 => n142, ZN => n190);
   U184 : AOI222_X1 port map( A1 => A_shifted(10), A2 => n177, B1 => 
                           zeroSignal(10), B2 => n168, C1 => A_neg_shifted(10),
                           C2 => n165, ZN => n189);
   U185 : NAND2_X1 port map( A1 => n192, A2 => n191, ZN => Y(11));
   U186 : AOI22_X1 port map( A1 => A_neg(11), A2 => n151, B1 => A_signal(11), 
                           B2 => n142, ZN => n192);
   U187 : AOI222_X1 port map( A1 => A_shifted(11), A2 => n177, B1 => 
                           zeroSignal(11), B2 => n168, C1 => A_neg_shifted(11),
                           C2 => n165, ZN => n191);
   U188 : NAND2_X1 port map( A1 => n194, A2 => n193, ZN => Y(12));
   U189 : AOI22_X1 port map( A1 => A_neg(12), A2 => n151, B1 => A_signal(12), 
                           B2 => n142, ZN => n194);
   U190 : AOI222_X1 port map( A1 => A_shifted(12), A2 => n177, B1 => 
                           zeroSignal(12), B2 => n168, C1 => A_neg_shifted(12),
                           C2 => n165, ZN => n193);
   U191 : NAND2_X1 port map( A1 => n196, A2 => n195, ZN => Y(13));
   U192 : AOI22_X1 port map( A1 => A_neg(13), A2 => n151, B1 => A_signal(13), 
                           B2 => n142, ZN => n196);
   U193 : AOI222_X1 port map( A1 => A_shifted(13), A2 => n177, B1 => 
                           zeroSignal(13), B2 => n168, C1 => A_neg_shifted(13),
                           C2 => n164, ZN => n195);
   U194 : NAND2_X1 port map( A1 => n198, A2 => n197, ZN => Y(14));
   U195 : AOI22_X1 port map( A1 => A_neg(14), A2 => n151, B1 => A_signal(14), 
                           B2 => n142, ZN => n198);
   U196 : AOI222_X1 port map( A1 => A_shifted(14), A2 => n177, B1 => 
                           zeroSignal(14), B2 => n168, C1 => A_neg_shifted(14),
                           C2 => n164, ZN => n197);
   U197 : NAND2_X1 port map( A1 => n200, A2 => n199, ZN => Y(15));
   U198 : AOI22_X1 port map( A1 => A_neg(15), A2 => n151, B1 => A_signal(15), 
                           B2 => n142, ZN => n200);
   U199 : AOI222_X1 port map( A1 => A_shifted(15), A2 => n177, B1 => 
                           zeroSignal(15), B2 => n168, C1 => A_neg_shifted(15),
                           C2 => n164, ZN => n199);
   U200 : NAND2_X1 port map( A1 => n202, A2 => n201, ZN => Y(16));
   U201 : AOI22_X1 port map( A1 => A_neg(16), A2 => n151, B1 => A_signal(16), 
                           B2 => n142, ZN => n202);
   U202 : AOI222_X1 port map( A1 => A_shifted(16), A2 => n177, B1 => 
                           zeroSignal(16), B2 => n168, C1 => A_neg_shifted(16),
                           C2 => n164, ZN => n201);
   U203 : NAND2_X1 port map( A1 => n204, A2 => n203, ZN => Y(17));
   U204 : AOI22_X1 port map( A1 => A_neg(17), A2 => n151, B1 => A_signal(17), 
                           B2 => n142, ZN => n204);
   U205 : AOI222_X1 port map( A1 => A_shifted(17), A2 => n177, B1 => 
                           zeroSignal(17), B2 => n168, C1 => A_neg_shifted(17),
                           C2 => n164, ZN => n203);
   U206 : NAND2_X1 port map( A1 => n206, A2 => n205, ZN => Y(18));
   U207 : AOI22_X1 port map( A1 => A_neg(18), A2 => n151, B1 => A_signal(18), 
                           B2 => n142, ZN => n206);
   U208 : AOI222_X1 port map( A1 => A_shifted(18), A2 => n177, B1 => 
                           zeroSignal(18), B2 => n168, C1 => A_neg_shifted(18),
                           C2 => n164, ZN => n205);
   U209 : NAND2_X1 port map( A1 => n208, A2 => n207, ZN => Y(19));
   U210 : AOI22_X1 port map( A1 => A_neg(19), A2 => n151, B1 => A_signal(19), 
                           B2 => n142, ZN => n208);
   U211 : AOI222_X1 port map( A1 => A_shifted(19), A2 => n177, B1 => 
                           zeroSignal(19), B2 => n168, C1 => A_neg_shifted(19),
                           C2 => n164, ZN => n207);
   U212 : NAND2_X1 port map( A1 => n212, A2 => n211, ZN => Y(20));
   U213 : AOI22_X1 port map( A1 => A_neg(20), A2 => n152, B1 => A_signal(20), 
                           B2 => n143, ZN => n212);
   U214 : AOI222_X1 port map( A1 => A_shifted(20), A2 => n178, B1 => 
                           zeroSignal(20), B2 => n169, C1 => A_neg_shifted(20),
                           C2 => n164, ZN => n211);
   U215 : NAND2_X1 port map( A1 => n214, A2 => n213, ZN => Y(21));
   U216 : AOI22_X1 port map( A1 => A_neg(21), A2 => n152, B1 => A_signal(21), 
                           B2 => n143, ZN => n214);
   U217 : AOI222_X1 port map( A1 => A_shifted(21), A2 => n178, B1 => 
                           zeroSignal(21), B2 => n169, C1 => A_neg_shifted(21),
                           C2 => n164, ZN => n213);
   U218 : NAND2_X1 port map( A1 => n216, A2 => n215, ZN => Y(22));
   U219 : AOI22_X1 port map( A1 => A_neg(22), A2 => n152, B1 => A_signal(22), 
                           B2 => n143, ZN => n216);
   U220 : AOI222_X1 port map( A1 => A_shifted(22), A2 => n178, B1 => 
                           zeroSignal(22), B2 => n169, C1 => A_neg_shifted(22),
                           C2 => n164, ZN => n215);
   U221 : NAND2_X1 port map( A1 => n218, A2 => n217, ZN => Y(23));
   U222 : AOI22_X1 port map( A1 => A_neg(23), A2 => n152, B1 => A_signal(23), 
                           B2 => n143, ZN => n218);
   U223 : AOI222_X1 port map( A1 => A_shifted(23), A2 => n178, B1 => 
                           zeroSignal(23), B2 => n169, C1 => A_neg_shifted(23),
                           C2 => n164, ZN => n217);
   U224 : NAND2_X1 port map( A1 => n220, A2 => n219, ZN => Y(24));
   U225 : AOI22_X1 port map( A1 => A_neg(24), A2 => n152, B1 => A_signal(24), 
                           B2 => n143, ZN => n220);
   U226 : AOI222_X1 port map( A1 => A_shifted(24), A2 => n178, B1 => 
                           zeroSignal(24), B2 => n169, C1 => A_neg_shifted(24),
                           C2 => n163, ZN => n219);
   U227 : NAND2_X1 port map( A1 => n222, A2 => n221, ZN => Y(25));
   U228 : AOI22_X1 port map( A1 => A_neg(25), A2 => n152, B1 => A_signal(25), 
                           B2 => n143, ZN => n222);
   U229 : AOI222_X1 port map( A1 => A_shifted(25), A2 => n178, B1 => 
                           zeroSignal(25), B2 => n169, C1 => A_neg_shifted(25),
                           C2 => n163, ZN => n221);
   U230 : NAND2_X1 port map( A1 => n224, A2 => n223, ZN => Y(26));
   U231 : AOI22_X1 port map( A1 => A_neg(26), A2 => n152, B1 => A_signal(26), 
                           B2 => n143, ZN => n224);
   U232 : AOI222_X1 port map( A1 => A_shifted(26), A2 => n178, B1 => 
                           zeroSignal(26), B2 => n169, C1 => A_neg_shifted(26),
                           C2 => n163, ZN => n223);
   U233 : NAND2_X1 port map( A1 => n226, A2 => n225, ZN => Y(27));
   U234 : AOI22_X1 port map( A1 => A_neg(27), A2 => n152, B1 => A_signal(27), 
                           B2 => n143, ZN => n226);
   U235 : AOI222_X1 port map( A1 => A_shifted(27), A2 => n178, B1 => 
                           zeroSignal(27), B2 => n169, C1 => A_neg_shifted(27),
                           C2 => n163, ZN => n225);
   U236 : NAND2_X1 port map( A1 => n228, A2 => n227, ZN => Y(28));
   U237 : AOI22_X1 port map( A1 => A_neg(28), A2 => n152, B1 => A_signal(28), 
                           B2 => n143, ZN => n228);
   U238 : AOI222_X1 port map( A1 => A_shifted(28), A2 => n178, B1 => 
                           zeroSignal(28), B2 => n169, C1 => A_neg_shifted(28),
                           C2 => n163, ZN => n227);
   U239 : NAND2_X1 port map( A1 => n230, A2 => n229, ZN => Y(29));
   U240 : AOI22_X1 port map( A1 => A_neg(29), A2 => n152, B1 => A_signal(29), 
                           B2 => n143, ZN => n230);
   U241 : AOI222_X1 port map( A1 => A_shifted(29), A2 => n178, B1 => 
                           zeroSignal(29), B2 => n169, C1 => A_neg_shifted(29),
                           C2 => n163, ZN => n229);
   U242 : AOI22_X1 port map( A1 => A_neg(36), A2 => n153, B1 => A_signal(36), 
                           B2 => n144, ZN => n246);
   U243 : AOI22_X1 port map( A1 => A_neg(35), A2 => n153, B1 => A_signal(35), 
                           B2 => n144, ZN => n244);
   U244 : AOI22_X1 port map( A1 => A_neg(33), A2 => n153, B1 => A_signal(33), 
                           B2 => n144, ZN => n240);

end SYN_BEHAVIORAL_2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity encoder_15 is

   port( pieceofB : in std_logic_vector (2 downto 0);  sel : out 
         std_logic_vector (2 downto 0));

end encoder_15;

architecture SYN_behavioral of encoder_15 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n7, n8, n9 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => pieceofB(1), A2 => pieceofB(0), ZN => n4);
   U4 : OR2_X1 port map( A1 => pieceofB(0), A2 => pieceofB(1), ZN => n5);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n8, ZN => n7);
   U6 : AND3_X2 port map( A1 => n7, A2 => n4, A3 => pieceofB(2), ZN => sel(2));
   U7 : INV_X1 port map( A => pieceofB(2), ZN => n9);
   U8 : AOI21_X1 port map( B1 => n7, B2 => n4, A => pieceofB(2), ZN => sel(0));
   U9 : OAI22_X1 port map( A1 => n7, A2 => n9, B1 => n4, B2 => pieceofB(2), ZN 
                           => sel(1));
   U10 : NAND2_X1 port map( A1 => pieceofB(1), A2 => pieceofB(0), ZN => n8);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity encoder_14 is

   port( pieceofB : in std_logic_vector (2 downto 0);  sel : out 
         std_logic_vector (2 downto 0));

end encoder_14;

architecture SYN_behavioral of encoder_14 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n6, n7 : std_logic;

begin
   
   U3 : INV_X1 port map( A => pieceofB(2), ZN => n7);
   U4 : AOI21_X1 port map( B1 => n5, B2 => n6, A => pieceofB(2), ZN => sel(0));
   U5 : AND3_X1 port map( A1 => pieceofB(2), A2 => n6, A3 => n5, ZN => sel(2));
   U6 : NAND2_X1 port map( A1 => pieceofB(1), A2 => pieceofB(0), ZN => n6);
   U7 : OAI22_X1 port map( A1 => n7, A2 => n5, B1 => pieceofB(2), B2 => n6, ZN 
                           => sel(1));
   U8 : OAI21_X1 port map( B1 => pieceofB(1), B2 => pieceofB(0), A => n6, ZN =>
                           n5);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity encoder_13 is

   port( pieceofB : in std_logic_vector (2 downto 0);  sel : out 
         std_logic_vector (2 downto 0));

end encoder_13;

architecture SYN_behavioral of encoder_13 is

   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n6, n7 : std_logic;

begin
   
   U3 : OAI22_X1 port map( A1 => n7, A2 => n5, B1 => pieceofB(2), B2 => n6, ZN 
                           => sel(1));
   U4 : INV_X1 port map( A => pieceofB(2), ZN => n7);
   U5 : OAI21_X1 port map( B1 => pieceofB(1), B2 => pieceofB(0), A => n6, ZN =>
                           n5);
   U6 : NAND2_X1 port map( A1 => pieceofB(1), A2 => pieceofB(0), ZN => n6);
   U7 : AOI21_X1 port map( B1 => n5, B2 => n6, A => pieceofB(2), ZN => sel(0));
   U8 : AND3_X1 port map( A1 => pieceofB(2), A2 => n6, A3 => n5, ZN => sel(2));

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity encoder_12 is

   port( pieceofB : in std_logic_vector (2 downto 0);  sel : out 
         std_logic_vector (2 downto 0));

end encoder_12;

architecture SYN_behavioral of encoder_12 is

   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n6, n7 : std_logic;

begin
   
   U3 : OAI22_X1 port map( A1 => n7, A2 => n5, B1 => pieceofB(2), B2 => n6, ZN 
                           => sel(1));
   U4 : INV_X1 port map( A => pieceofB(2), ZN => n7);
   U5 : OAI21_X1 port map( B1 => pieceofB(1), B2 => pieceofB(0), A => n6, ZN =>
                           n5);
   U6 : NAND2_X1 port map( A1 => pieceofB(1), A2 => pieceofB(0), ZN => n6);
   U7 : AOI21_X1 port map( B1 => n5, B2 => n6, A => pieceofB(2), ZN => sel(0));
   U8 : AND3_X1 port map( A1 => pieceofB(2), A2 => n6, A3 => n5, ZN => sel(2));

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity encoder_11 is

   port( pieceofB : in std_logic_vector (2 downto 0);  sel : out 
         std_logic_vector (2 downto 0));

end encoder_11;

architecture SYN_behavioral of encoder_11 is

   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n6, n7 : std_logic;

begin
   
   U3 : OAI22_X1 port map( A1 => n7, A2 => n5, B1 => pieceofB(2), B2 => n6, ZN 
                           => sel(1));
   U4 : INV_X1 port map( A => pieceofB(2), ZN => n7);
   U5 : OAI21_X1 port map( B1 => pieceofB(1), B2 => pieceofB(0), A => n6, ZN =>
                           n5);
   U6 : NAND2_X1 port map( A1 => pieceofB(1), A2 => pieceofB(0), ZN => n6);
   U7 : AOI21_X1 port map( B1 => n5, B2 => n6, A => pieceofB(2), ZN => sel(0));
   U8 : AND3_X1 port map( A1 => pieceofB(2), A2 => n6, A3 => n5, ZN => sel(2));

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity encoder_10 is

   port( pieceofB : in std_logic_vector (2 downto 0);  sel : out 
         std_logic_vector (2 downto 0));

end encoder_10;

architecture SYN_behavioral of encoder_10 is

   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n6, n7 : std_logic;

begin
   
   U3 : OAI22_X1 port map( A1 => n7, A2 => n5, B1 => pieceofB(2), B2 => n6, ZN 
                           => sel(1));
   U4 : INV_X1 port map( A => pieceofB(2), ZN => n7);
   U5 : OAI21_X1 port map( B1 => pieceofB(1), B2 => pieceofB(0), A => n6, ZN =>
                           n5);
   U6 : NAND2_X1 port map( A1 => pieceofB(1), A2 => pieceofB(0), ZN => n6);
   U7 : AOI21_X1 port map( B1 => n5, B2 => n6, A => pieceofB(2), ZN => sel(0));
   U8 : AND3_X1 port map( A1 => pieceofB(2), A2 => n6, A3 => n5, ZN => sel(2));

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity encoder_9 is

   port( pieceofB : in std_logic_vector (2 downto 0);  sel : out 
         std_logic_vector (2 downto 0));

end encoder_9;

architecture SYN_behavioral of encoder_9 is

   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n6, n7 : std_logic;

begin
   
   U3 : OAI22_X1 port map( A1 => n7, A2 => n5, B1 => pieceofB(2), B2 => n6, ZN 
                           => sel(1));
   U4 : INV_X1 port map( A => pieceofB(2), ZN => n7);
   U5 : OAI21_X1 port map( B1 => pieceofB(1), B2 => pieceofB(0), A => n6, ZN =>
                           n5);
   U6 : NAND2_X1 port map( A1 => pieceofB(1), A2 => pieceofB(0), ZN => n6);
   U7 : AOI21_X1 port map( B1 => n5, B2 => n6, A => pieceofB(2), ZN => sel(0));
   U8 : AND3_X1 port map( A1 => pieceofB(2), A2 => n6, A3 => n5, ZN => sel(2));

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity encoder_8 is

   port( pieceofB : in std_logic_vector (2 downto 0);  sel : out 
         std_logic_vector (2 downto 0));

end encoder_8;

architecture SYN_behavioral of encoder_8 is

   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n6, n7 : std_logic;

begin
   
   U3 : OAI22_X1 port map( A1 => n7, A2 => n5, B1 => pieceofB(2), B2 => n6, ZN 
                           => sel(1));
   U4 : INV_X1 port map( A => pieceofB(2), ZN => n7);
   U5 : OAI21_X1 port map( B1 => pieceofB(1), B2 => pieceofB(0), A => n6, ZN =>
                           n5);
   U6 : NAND2_X1 port map( A1 => pieceofB(1), A2 => pieceofB(0), ZN => n6);
   U7 : AOI21_X1 port map( B1 => n5, B2 => n6, A => pieceofB(2), ZN => sel(0));
   U8 : AND3_X1 port map( A1 => pieceofB(2), A2 => n6, A3 => n5, ZN => sel(2));

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity encoder_7 is

   port( pieceofB : in std_logic_vector (2 downto 0);  sel : out 
         std_logic_vector (2 downto 0));

end encoder_7;

architecture SYN_behavioral of encoder_7 is

   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n6, n7 : std_logic;

begin
   
   U3 : OAI22_X1 port map( A1 => n7, A2 => n5, B1 => pieceofB(2), B2 => n6, ZN 
                           => sel(1));
   U4 : INV_X1 port map( A => pieceofB(2), ZN => n7);
   U5 : OAI21_X1 port map( B1 => pieceofB(1), B2 => pieceofB(0), A => n6, ZN =>
                           n5);
   U6 : NAND2_X1 port map( A1 => pieceofB(1), A2 => pieceofB(0), ZN => n6);
   U7 : AOI21_X1 port map( B1 => n5, B2 => n6, A => pieceofB(2), ZN => sel(0));
   U8 : AND3_X1 port map( A1 => pieceofB(2), A2 => n6, A3 => n5, ZN => sel(2));

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity encoder_6 is

   port( pieceofB : in std_logic_vector (2 downto 0);  sel : out 
         std_logic_vector (2 downto 0));

end encoder_6;

architecture SYN_behavioral of encoder_6 is

   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n6, n7 : std_logic;

begin
   
   U3 : OAI22_X1 port map( A1 => n7, A2 => n5, B1 => pieceofB(2), B2 => n6, ZN 
                           => sel(1));
   U4 : INV_X1 port map( A => pieceofB(2), ZN => n7);
   U5 : OAI21_X1 port map( B1 => pieceofB(1), B2 => pieceofB(0), A => n6, ZN =>
                           n5);
   U6 : NAND2_X1 port map( A1 => pieceofB(1), A2 => pieceofB(0), ZN => n6);
   U7 : AOI21_X1 port map( B1 => n5, B2 => n6, A => pieceofB(2), ZN => sel(0));
   U8 : AND3_X1 port map( A1 => pieceofB(2), A2 => n6, A3 => n5, ZN => sel(2));

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity encoder_5 is

   port( pieceofB : in std_logic_vector (2 downto 0);  sel : out 
         std_logic_vector (2 downto 0));

end encoder_5;

architecture SYN_behavioral of encoder_5 is

   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n6, n7 : std_logic;

begin
   
   U3 : OAI22_X1 port map( A1 => n7, A2 => n5, B1 => pieceofB(2), B2 => n6, ZN 
                           => sel(1));
   U4 : INV_X1 port map( A => pieceofB(2), ZN => n7);
   U5 : OAI21_X1 port map( B1 => pieceofB(1), B2 => pieceofB(0), A => n6, ZN =>
                           n5);
   U6 : NAND2_X1 port map( A1 => pieceofB(1), A2 => pieceofB(0), ZN => n6);
   U7 : AOI21_X1 port map( B1 => n5, B2 => n6, A => pieceofB(2), ZN => sel(0));
   U8 : AND3_X1 port map( A1 => pieceofB(2), A2 => n6, A3 => n5, ZN => sel(2));

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity encoder_4 is

   port( pieceofB : in std_logic_vector (2 downto 0);  sel : out 
         std_logic_vector (2 downto 0));

end encoder_4;

architecture SYN_behavioral of encoder_4 is

   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n6, n7 : std_logic;

begin
   
   U3 : OAI22_X1 port map( A1 => n7, A2 => n5, B1 => pieceofB(2), B2 => n6, ZN 
                           => sel(1));
   U4 : INV_X1 port map( A => pieceofB(2), ZN => n7);
   U5 : OAI21_X1 port map( B1 => pieceofB(1), B2 => pieceofB(0), A => n6, ZN =>
                           n5);
   U6 : NAND2_X1 port map( A1 => pieceofB(1), A2 => pieceofB(0), ZN => n6);
   U7 : AOI21_X1 port map( B1 => n5, B2 => n6, A => pieceofB(2), ZN => sel(0));
   U8 : AND3_X1 port map( A1 => pieceofB(2), A2 => n6, A3 => n5, ZN => sel(2));

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity encoder_3 is

   port( pieceofB : in std_logic_vector (2 downto 0);  sel : out 
         std_logic_vector (2 downto 0));

end encoder_3;

architecture SYN_behavioral of encoder_3 is

   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n6, n7 : std_logic;

begin
   
   U3 : OAI22_X1 port map( A1 => n7, A2 => n5, B1 => pieceofB(2), B2 => n6, ZN 
                           => sel(1));
   U4 : INV_X1 port map( A => pieceofB(2), ZN => n7);
   U5 : OAI21_X1 port map( B1 => pieceofB(1), B2 => pieceofB(0), A => n6, ZN =>
                           n5);
   U6 : NAND2_X1 port map( A1 => pieceofB(1), A2 => pieceofB(0), ZN => n6);
   U7 : AOI21_X1 port map( B1 => n5, B2 => n6, A => pieceofB(2), ZN => sel(0));
   U8 : AND3_X1 port map( A1 => pieceofB(2), A2 => n6, A3 => n5, ZN => sel(2));

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity encoder_2 is

   port( pieceofB : in std_logic_vector (2 downto 0);  sel : out 
         std_logic_vector (2 downto 0));

end encoder_2;

architecture SYN_behavioral of encoder_2 is

   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n6, n7 : std_logic;

begin
   
   U3 : OAI22_X1 port map( A1 => n7, A2 => n5, B1 => pieceofB(2), B2 => n6, ZN 
                           => sel(1));
   U4 : INV_X1 port map( A => pieceofB(2), ZN => n7);
   U5 : OAI21_X1 port map( B1 => pieceofB(1), B2 => pieceofB(0), A => n6, ZN =>
                           n5);
   U6 : NAND2_X1 port map( A1 => pieceofB(1), A2 => pieceofB(0), ZN => n6);
   U7 : AOI21_X1 port map( B1 => n5, B2 => n6, A => pieceofB(2), ZN => sel(0));
   U8 : AND3_X1 port map( A1 => pieceofB(2), A2 => n6, A3 => n5, ZN => sel(2));

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity encoder_1 is

   port( pieceofB : in std_logic_vector (2 downto 0);  sel : out 
         std_logic_vector (2 downto 0));

end encoder_1;

architecture SYN_behavioral of encoder_1 is

   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n6, n7 : std_logic;

begin
   
   U3 : OAI22_X1 port map( A1 => n7, A2 => n5, B1 => pieceofB(2), B2 => n6, ZN 
                           => sel(1));
   U4 : INV_X1 port map( A => pieceofB(2), ZN => n7);
   U5 : OAI21_X1 port map( B1 => pieceofB(1), B2 => pieceofB(0), A => n6, ZN =>
                           n5);
   U6 : NAND2_X1 port map( A1 => pieceofB(1), A2 => pieceofB(0), ZN => n6);
   U7 : AOI21_X1 port map( B1 => n5, B2 => n6, A => pieceofB(2), ZN => sel(0));
   U8 : AND3_X1 port map( A1 => pieceofB(2), A2 => n6, A3 => n5, ZN => sel(2));

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity leftshifter_NbitShifter64_62 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_62;

architecture SYN_behavioral of leftshifter_NbitShifter64_62 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity leftshifter_NbitShifter64_61 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_61;

architecture SYN_behavioral of leftshifter_NbitShifter64_61 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity leftshifter_NbitShifter64_60 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_60;

architecture SYN_behavioral of leftshifter_NbitShifter64_60 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity leftshifter_NbitShifter64_59 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_59;

architecture SYN_behavioral of leftshifter_NbitShifter64_59 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity leftshifter_NbitShifter64_58 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_58;

architecture SYN_behavioral of leftshifter_NbitShifter64_58 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity leftshifter_NbitShifter64_57 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_57;

architecture SYN_behavioral of leftshifter_NbitShifter64_57 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity leftshifter_NbitShifter64_56 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_56;

architecture SYN_behavioral of leftshifter_NbitShifter64_56 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity leftshifter_NbitShifter64_55 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_55;

architecture SYN_behavioral of leftshifter_NbitShifter64_55 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity leftshifter_NbitShifter64_54 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_54;

architecture SYN_behavioral of leftshifter_NbitShifter64_54 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity leftshifter_NbitShifter64_53 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_53;

architecture SYN_behavioral of leftshifter_NbitShifter64_53 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity leftshifter_NbitShifter64_52 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_52;

architecture SYN_behavioral of leftshifter_NbitShifter64_52 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity leftshifter_NbitShifter64_51 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_51;

architecture SYN_behavioral of leftshifter_NbitShifter64_51 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity leftshifter_NbitShifter64_50 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_50;

architecture SYN_behavioral of leftshifter_NbitShifter64_50 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity leftshifter_NbitShifter64_49 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_49;

architecture SYN_behavioral of leftshifter_NbitShifter64_49 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity leftshifter_NbitShifter64_48 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_48;

architecture SYN_behavioral of leftshifter_NbitShifter64_48 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity leftshifter_NbitShifter64_47 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_47;

architecture SYN_behavioral of leftshifter_NbitShifter64_47 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity leftshifter_NbitShifter64_46 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_46;

architecture SYN_behavioral of leftshifter_NbitShifter64_46 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity leftshifter_NbitShifter64_45 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_45;

architecture SYN_behavioral of leftshifter_NbitShifter64_45 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity leftshifter_NbitShifter64_44 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_44;

architecture SYN_behavioral of leftshifter_NbitShifter64_44 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity leftshifter_NbitShifter64_43 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_43;

architecture SYN_behavioral of leftshifter_NbitShifter64_43 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity leftshifter_NbitShifter64_42 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_42;

architecture SYN_behavioral of leftshifter_NbitShifter64_42 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity leftshifter_NbitShifter64_41 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_41;

architecture SYN_behavioral of leftshifter_NbitShifter64_41 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity leftshifter_NbitShifter64_40 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_40;

architecture SYN_behavioral of leftshifter_NbitShifter64_40 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity leftshifter_NbitShifter64_39 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_39;

architecture SYN_behavioral of leftshifter_NbitShifter64_39 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity leftshifter_NbitShifter64_38 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_38;

architecture SYN_behavioral of leftshifter_NbitShifter64_38 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity leftshifter_NbitShifter64_37 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_37;

architecture SYN_behavioral of leftshifter_NbitShifter64_37 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity leftshifter_NbitShifter64_36 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_36;

architecture SYN_behavioral of leftshifter_NbitShifter64_36 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity leftshifter_NbitShifter64_35 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_35;

architecture SYN_behavioral of leftshifter_NbitShifter64_35 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity leftshifter_NbitShifter64_34 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_34;

architecture SYN_behavioral of leftshifter_NbitShifter64_34 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity leftshifter_NbitShifter64_33 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_33;

architecture SYN_behavioral of leftshifter_NbitShifter64_33 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity leftshifter_NbitShifter64_32 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_32;

architecture SYN_behavioral of leftshifter_NbitShifter64_32 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity leftshifter_NbitShifter64_31 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_31;

architecture SYN_behavioral of leftshifter_NbitShifter64_31 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity leftshifter_NbitShifter64_30 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_30;

architecture SYN_behavioral of leftshifter_NbitShifter64_30 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity leftshifter_NbitShifter64_29 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_29;

architecture SYN_behavioral of leftshifter_NbitShifter64_29 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity leftshifter_NbitShifter64_28 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_28;

architecture SYN_behavioral of leftshifter_NbitShifter64_28 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity leftshifter_NbitShifter64_27 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_27;

architecture SYN_behavioral of leftshifter_NbitShifter64_27 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity leftshifter_NbitShifter64_26 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_26;

architecture SYN_behavioral of leftshifter_NbitShifter64_26 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity leftshifter_NbitShifter64_25 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_25;

architecture SYN_behavioral of leftshifter_NbitShifter64_25 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity leftshifter_NbitShifter64_24 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_24;

architecture SYN_behavioral of leftshifter_NbitShifter64_24 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity leftshifter_NbitShifter64_23 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_23;

architecture SYN_behavioral of leftshifter_NbitShifter64_23 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity leftshifter_NbitShifter64_22 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_22;

architecture SYN_behavioral of leftshifter_NbitShifter64_22 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity leftshifter_NbitShifter64_21 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_21;

architecture SYN_behavioral of leftshifter_NbitShifter64_21 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity leftshifter_NbitShifter64_20 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_20;

architecture SYN_behavioral of leftshifter_NbitShifter64_20 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity leftshifter_NbitShifter64_19 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_19;

architecture SYN_behavioral of leftshifter_NbitShifter64_19 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity leftshifter_NbitShifter64_18 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_18;

architecture SYN_behavioral of leftshifter_NbitShifter64_18 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity leftshifter_NbitShifter64_17 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_17;

architecture SYN_behavioral of leftshifter_NbitShifter64_17 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity leftshifter_NbitShifter64_16 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_16;

architecture SYN_behavioral of leftshifter_NbitShifter64_16 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity leftshifter_NbitShifter64_15 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_15;

architecture SYN_behavioral of leftshifter_NbitShifter64_15 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity leftshifter_NbitShifter64_14 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_14;

architecture SYN_behavioral of leftshifter_NbitShifter64_14 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity leftshifter_NbitShifter64_13 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_13;

architecture SYN_behavioral of leftshifter_NbitShifter64_13 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity leftshifter_NbitShifter64_12 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_12;

architecture SYN_behavioral of leftshifter_NbitShifter64_12 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity leftshifter_NbitShifter64_11 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_11;

architecture SYN_behavioral of leftshifter_NbitShifter64_11 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity leftshifter_NbitShifter64_10 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_10;

architecture SYN_behavioral of leftshifter_NbitShifter64_10 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity leftshifter_NbitShifter64_9 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_9;

architecture SYN_behavioral of leftshifter_NbitShifter64_9 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity leftshifter_NbitShifter64_8 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_8;

architecture SYN_behavioral of leftshifter_NbitShifter64_8 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity leftshifter_NbitShifter64_7 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_7;

architecture SYN_behavioral of leftshifter_NbitShifter64_7 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity leftshifter_NbitShifter64_6 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_6;

architecture SYN_behavioral of leftshifter_NbitShifter64_6 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity leftshifter_NbitShifter64_5 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_5;

architecture SYN_behavioral of leftshifter_NbitShifter64_5 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity leftshifter_NbitShifter64_4 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_4;

architecture SYN_behavioral of leftshifter_NbitShifter64_4 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity leftshifter_NbitShifter64_3 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_3;

architecture SYN_behavioral of leftshifter_NbitShifter64_3 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity leftshifter_NbitShifter64_2 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_2;

architecture SYN_behavioral of leftshifter_NbitShifter64_2 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity leftshifter_NbitShifter64_1 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_1;

architecture SYN_behavioral of leftshifter_NbitShifter64_1 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity RCA_NbitRca64_14 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_NbitRca64_14;

architecture SYN_STRUCTURAL of RCA_NbitRca64_14 is

   component FA_833
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_834
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_835
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_836
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_837
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_838
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_839
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_840
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_841
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_842
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_843
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_844
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_845
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_846
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_847
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_848
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_849
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_850
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_851
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_852
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_853
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_854
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_855
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_856
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_857
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_858
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_859
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_860
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_861
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_862
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_863
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_864
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_865
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_866
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_867
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_868
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_869
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_870
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_871
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_872
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_873
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_874
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_875
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_876
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_877
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_878
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_879
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_880
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_881
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_882
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_883
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_884
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_885
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_886
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_887
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_888
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_889
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_890
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_891
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_892
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_893
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_894
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_895
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_896
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_63_port, CTMP_62_port, CTMP_61_port, CTMP_60_port, CTMP_59_port,
      CTMP_58_port, CTMP_57_port, CTMP_56_port, CTMP_55_port, CTMP_54_port, 
      CTMP_53_port, CTMP_52_port, CTMP_51_port, CTMP_50_port, CTMP_49_port, 
      CTMP_48_port, CTMP_47_port, CTMP_46_port, CTMP_45_port, CTMP_44_port, 
      CTMP_43_port, CTMP_42_port, CTMP_41_port, CTMP_40_port, CTMP_39_port, 
      CTMP_38_port, CTMP_37_port, CTMP_36_port, CTMP_35_port, CTMP_34_port, 
      CTMP_33_port, CTMP_32_port, CTMP_31_port, CTMP_30_port, CTMP_29_port, 
      CTMP_28_port, CTMP_27_port, CTMP_26_port, CTMP_25_port, CTMP_24_port, 
      CTMP_23_port, CTMP_22_port, CTMP_21_port, CTMP_20_port, CTMP_19_port, 
      CTMP_18_port, CTMP_17_port, CTMP_16_port, CTMP_15_port, CTMP_14_port, 
      CTMP_13_port, CTMP_12_port, CTMP_11_port, CTMP_10_port, CTMP_9_port, 
      CTMP_8_port, CTMP_7_port, CTMP_6_port, CTMP_5_port, CTMP_4_port, 
      CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_896 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_895 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_894 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_893 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => CTMP_4_port);
   FAI_5 : FA_892 port map( A => A(4), B => B(4), Ci => CTMP_4_port, S => S(4),
                           Co => CTMP_5_port);
   FAI_6 : FA_891 port map( A => A(5), B => B(5), Ci => CTMP_5_port, S => S(5),
                           Co => CTMP_6_port);
   FAI_7 : FA_890 port map( A => A(6), B => B(6), Ci => CTMP_6_port, S => S(6),
                           Co => CTMP_7_port);
   FAI_8 : FA_889 port map( A => A(7), B => B(7), Ci => CTMP_7_port, S => S(7),
                           Co => CTMP_8_port);
   FAI_9 : FA_888 port map( A => A(8), B => B(8), Ci => CTMP_8_port, S => S(8),
                           Co => CTMP_9_port);
   FAI_10 : FA_887 port map( A => A(9), B => B(9), Ci => CTMP_9_port, S => S(9)
                           , Co => CTMP_10_port);
   FAI_11 : FA_886 port map( A => A(10), B => B(10), Ci => CTMP_10_port, S => 
                           S(10), Co => CTMP_11_port);
   FAI_12 : FA_885 port map( A => A(11), B => B(11), Ci => CTMP_11_port, S => 
                           S(11), Co => CTMP_12_port);
   FAI_13 : FA_884 port map( A => A(12), B => B(12), Ci => CTMP_12_port, S => 
                           S(12), Co => CTMP_13_port);
   FAI_14 : FA_883 port map( A => A(13), B => B(13), Ci => CTMP_13_port, S => 
                           S(13), Co => CTMP_14_port);
   FAI_15 : FA_882 port map( A => A(14), B => B(14), Ci => CTMP_14_port, S => 
                           S(14), Co => CTMP_15_port);
   FAI_16 : FA_881 port map( A => A(15), B => B(15), Ci => CTMP_15_port, S => 
                           S(15), Co => CTMP_16_port);
   FAI_17 : FA_880 port map( A => A(16), B => B(16), Ci => CTMP_16_port, S => 
                           S(16), Co => CTMP_17_port);
   FAI_18 : FA_879 port map( A => A(17), B => B(17), Ci => CTMP_17_port, S => 
                           S(17), Co => CTMP_18_port);
   FAI_19 : FA_878 port map( A => A(18), B => B(18), Ci => CTMP_18_port, S => 
                           S(18), Co => CTMP_19_port);
   FAI_20 : FA_877 port map( A => A(19), B => B(19), Ci => CTMP_19_port, S => 
                           S(19), Co => CTMP_20_port);
   FAI_21 : FA_876 port map( A => A(20), B => B(20), Ci => CTMP_20_port, S => 
                           S(20), Co => CTMP_21_port);
   FAI_22 : FA_875 port map( A => A(21), B => B(21), Ci => CTMP_21_port, S => 
                           S(21), Co => CTMP_22_port);
   FAI_23 : FA_874 port map( A => A(22), B => B(22), Ci => CTMP_22_port, S => 
                           S(22), Co => CTMP_23_port);
   FAI_24 : FA_873 port map( A => A(23), B => B(23), Ci => CTMP_23_port, S => 
                           S(23), Co => CTMP_24_port);
   FAI_25 : FA_872 port map( A => A(24), B => B(24), Ci => CTMP_24_port, S => 
                           S(24), Co => CTMP_25_port);
   FAI_26 : FA_871 port map( A => A(25), B => B(25), Ci => CTMP_25_port, S => 
                           S(25), Co => CTMP_26_port);
   FAI_27 : FA_870 port map( A => A(26), B => B(26), Ci => CTMP_26_port, S => 
                           S(26), Co => CTMP_27_port);
   FAI_28 : FA_869 port map( A => A(27), B => B(27), Ci => CTMP_27_port, S => 
                           S(27), Co => CTMP_28_port);
   FAI_29 : FA_868 port map( A => A(28), B => B(28), Ci => CTMP_28_port, S => 
                           S(28), Co => CTMP_29_port);
   FAI_30 : FA_867 port map( A => A(29), B => B(29), Ci => CTMP_29_port, S => 
                           S(29), Co => CTMP_30_port);
   FAI_31 : FA_866 port map( A => A(30), B => B(30), Ci => CTMP_30_port, S => 
                           S(30), Co => CTMP_31_port);
   FAI_32 : FA_865 port map( A => A(31), B => B(31), Ci => CTMP_31_port, S => 
                           S(31), Co => CTMP_32_port);
   FAI_33 : FA_864 port map( A => A(32), B => B(32), Ci => CTMP_32_port, S => 
                           S(32), Co => CTMP_33_port);
   FAI_34 : FA_863 port map( A => A(33), B => B(33), Ci => CTMP_33_port, S => 
                           S(33), Co => CTMP_34_port);
   FAI_35 : FA_862 port map( A => A(34), B => B(34), Ci => CTMP_34_port, S => 
                           S(34), Co => CTMP_35_port);
   FAI_36 : FA_861 port map( A => A(35), B => B(35), Ci => CTMP_35_port, S => 
                           S(35), Co => CTMP_36_port);
   FAI_37 : FA_860 port map( A => A(36), B => B(36), Ci => CTMP_36_port, S => 
                           S(36), Co => CTMP_37_port);
   FAI_38 : FA_859 port map( A => A(37), B => B(37), Ci => CTMP_37_port, S => 
                           S(37), Co => CTMP_38_port);
   FAI_39 : FA_858 port map( A => A(38), B => B(38), Ci => CTMP_38_port, S => 
                           S(38), Co => CTMP_39_port);
   FAI_40 : FA_857 port map( A => A(39), B => B(39), Ci => CTMP_39_port, S => 
                           S(39), Co => CTMP_40_port);
   FAI_41 : FA_856 port map( A => A(40), B => B(40), Ci => CTMP_40_port, S => 
                           S(40), Co => CTMP_41_port);
   FAI_42 : FA_855 port map( A => A(41), B => B(41), Ci => CTMP_41_port, S => 
                           S(41), Co => CTMP_42_port);
   FAI_43 : FA_854 port map( A => A(42), B => B(42), Ci => CTMP_42_port, S => 
                           S(42), Co => CTMP_43_port);
   FAI_44 : FA_853 port map( A => A(43), B => B(43), Ci => CTMP_43_port, S => 
                           S(43), Co => CTMP_44_port);
   FAI_45 : FA_852 port map( A => A(44), B => B(44), Ci => CTMP_44_port, S => 
                           S(44), Co => CTMP_45_port);
   FAI_46 : FA_851 port map( A => A(45), B => B(45), Ci => CTMP_45_port, S => 
                           S(45), Co => CTMP_46_port);
   FAI_47 : FA_850 port map( A => A(46), B => B(46), Ci => CTMP_46_port, S => 
                           S(46), Co => CTMP_47_port);
   FAI_48 : FA_849 port map( A => A(47), B => B(47), Ci => CTMP_47_port, S => 
                           S(47), Co => CTMP_48_port);
   FAI_49 : FA_848 port map( A => A(48), B => B(48), Ci => CTMP_48_port, S => 
                           S(48), Co => CTMP_49_port);
   FAI_50 : FA_847 port map( A => A(49), B => B(49), Ci => CTMP_49_port, S => 
                           S(49), Co => CTMP_50_port);
   FAI_51 : FA_846 port map( A => A(50), B => B(50), Ci => CTMP_50_port, S => 
                           S(50), Co => CTMP_51_port);
   FAI_52 : FA_845 port map( A => A(51), B => B(51), Ci => CTMP_51_port, S => 
                           S(51), Co => CTMP_52_port);
   FAI_53 : FA_844 port map( A => A(52), B => B(52), Ci => CTMP_52_port, S => 
                           S(52), Co => CTMP_53_port);
   FAI_54 : FA_843 port map( A => A(53), B => B(53), Ci => CTMP_53_port, S => 
                           S(53), Co => CTMP_54_port);
   FAI_55 : FA_842 port map( A => A(54), B => B(54), Ci => CTMP_54_port, S => 
                           S(54), Co => CTMP_55_port);
   FAI_56 : FA_841 port map( A => A(55), B => B(55), Ci => CTMP_55_port, S => 
                           S(55), Co => CTMP_56_port);
   FAI_57 : FA_840 port map( A => A(56), B => B(56), Ci => CTMP_56_port, S => 
                           S(56), Co => CTMP_57_port);
   FAI_58 : FA_839 port map( A => A(57), B => B(57), Ci => CTMP_57_port, S => 
                           S(57), Co => CTMP_58_port);
   FAI_59 : FA_838 port map( A => A(58), B => B(58), Ci => CTMP_58_port, S => 
                           S(58), Co => CTMP_59_port);
   FAI_60 : FA_837 port map( A => A(59), B => B(59), Ci => CTMP_59_port, S => 
                           S(59), Co => CTMP_60_port);
   FAI_61 : FA_836 port map( A => A(60), B => B(60), Ci => CTMP_60_port, S => 
                           S(60), Co => CTMP_61_port);
   FAI_62 : FA_835 port map( A => A(61), B => B(61), Ci => CTMP_61_port, S => 
                           S(61), Co => CTMP_62_port);
   FAI_63 : FA_834 port map( A => A(62), B => B(62), Ci => CTMP_62_port, S => 
                           S(62), Co => CTMP_63_port);
   FAI_64 : FA_833 port map( A => A(63), B => B(63), Ci => CTMP_63_port, S => 
                           S(63), Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity RCA_NbitRca64_13 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_NbitRca64_13;

architecture SYN_STRUCTURAL of RCA_NbitRca64_13 is

   component FA_769
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_770
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_771
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_772
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_773
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_774
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_775
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_776
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_777
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_778
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_779
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_780
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_781
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_782
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_783
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_784
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_785
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_786
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_787
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_788
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_789
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_790
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_791
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_792
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_793
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_794
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_795
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_796
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_797
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_798
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_799
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_800
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_801
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_802
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_803
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_804
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_805
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_806
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_807
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_808
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_809
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_810
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_811
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_812
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_813
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_814
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_815
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_816
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_817
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_818
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_819
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_820
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_821
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_822
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_823
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_824
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_825
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_826
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_827
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_828
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_829
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_830
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_831
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_832
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_63_port, CTMP_62_port, CTMP_61_port, CTMP_60_port, CTMP_59_port,
      CTMP_58_port, CTMP_57_port, CTMP_56_port, CTMP_55_port, CTMP_54_port, 
      CTMP_53_port, CTMP_52_port, CTMP_51_port, CTMP_50_port, CTMP_49_port, 
      CTMP_48_port, CTMP_47_port, CTMP_46_port, CTMP_45_port, CTMP_44_port, 
      CTMP_43_port, CTMP_42_port, CTMP_41_port, CTMP_40_port, CTMP_39_port, 
      CTMP_38_port, CTMP_37_port, CTMP_36_port, CTMP_35_port, CTMP_34_port, 
      CTMP_33_port, CTMP_32_port, CTMP_31_port, CTMP_30_port, CTMP_29_port, 
      CTMP_28_port, CTMP_27_port, CTMP_26_port, CTMP_25_port, CTMP_24_port, 
      CTMP_23_port, CTMP_22_port, CTMP_21_port, CTMP_20_port, CTMP_19_port, 
      CTMP_18_port, CTMP_17_port, CTMP_16_port, CTMP_15_port, CTMP_14_port, 
      CTMP_13_port, CTMP_12_port, CTMP_11_port, CTMP_10_port, CTMP_9_port, 
      CTMP_8_port, CTMP_7_port, CTMP_6_port, CTMP_5_port, CTMP_4_port, 
      CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_832 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_831 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_830 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_829 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => CTMP_4_port);
   FAI_5 : FA_828 port map( A => A(4), B => B(4), Ci => CTMP_4_port, S => S(4),
                           Co => CTMP_5_port);
   FAI_6 : FA_827 port map( A => A(5), B => B(5), Ci => CTMP_5_port, S => S(5),
                           Co => CTMP_6_port);
   FAI_7 : FA_826 port map( A => A(6), B => B(6), Ci => CTMP_6_port, S => S(6),
                           Co => CTMP_7_port);
   FAI_8 : FA_825 port map( A => A(7), B => B(7), Ci => CTMP_7_port, S => S(7),
                           Co => CTMP_8_port);
   FAI_9 : FA_824 port map( A => A(8), B => B(8), Ci => CTMP_8_port, S => S(8),
                           Co => CTMP_9_port);
   FAI_10 : FA_823 port map( A => A(9), B => B(9), Ci => CTMP_9_port, S => S(9)
                           , Co => CTMP_10_port);
   FAI_11 : FA_822 port map( A => A(10), B => B(10), Ci => CTMP_10_port, S => 
                           S(10), Co => CTMP_11_port);
   FAI_12 : FA_821 port map( A => A(11), B => B(11), Ci => CTMP_11_port, S => 
                           S(11), Co => CTMP_12_port);
   FAI_13 : FA_820 port map( A => A(12), B => B(12), Ci => CTMP_12_port, S => 
                           S(12), Co => CTMP_13_port);
   FAI_14 : FA_819 port map( A => A(13), B => B(13), Ci => CTMP_13_port, S => 
                           S(13), Co => CTMP_14_port);
   FAI_15 : FA_818 port map( A => A(14), B => B(14), Ci => CTMP_14_port, S => 
                           S(14), Co => CTMP_15_port);
   FAI_16 : FA_817 port map( A => A(15), B => B(15), Ci => CTMP_15_port, S => 
                           S(15), Co => CTMP_16_port);
   FAI_17 : FA_816 port map( A => A(16), B => B(16), Ci => CTMP_16_port, S => 
                           S(16), Co => CTMP_17_port);
   FAI_18 : FA_815 port map( A => A(17), B => B(17), Ci => CTMP_17_port, S => 
                           S(17), Co => CTMP_18_port);
   FAI_19 : FA_814 port map( A => A(18), B => B(18), Ci => CTMP_18_port, S => 
                           S(18), Co => CTMP_19_port);
   FAI_20 : FA_813 port map( A => A(19), B => B(19), Ci => CTMP_19_port, S => 
                           S(19), Co => CTMP_20_port);
   FAI_21 : FA_812 port map( A => A(20), B => B(20), Ci => CTMP_20_port, S => 
                           S(20), Co => CTMP_21_port);
   FAI_22 : FA_811 port map( A => A(21), B => B(21), Ci => CTMP_21_port, S => 
                           S(21), Co => CTMP_22_port);
   FAI_23 : FA_810 port map( A => A(22), B => B(22), Ci => CTMP_22_port, S => 
                           S(22), Co => CTMP_23_port);
   FAI_24 : FA_809 port map( A => A(23), B => B(23), Ci => CTMP_23_port, S => 
                           S(23), Co => CTMP_24_port);
   FAI_25 : FA_808 port map( A => A(24), B => B(24), Ci => CTMP_24_port, S => 
                           S(24), Co => CTMP_25_port);
   FAI_26 : FA_807 port map( A => A(25), B => B(25), Ci => CTMP_25_port, S => 
                           S(25), Co => CTMP_26_port);
   FAI_27 : FA_806 port map( A => A(26), B => B(26), Ci => CTMP_26_port, S => 
                           S(26), Co => CTMP_27_port);
   FAI_28 : FA_805 port map( A => A(27), B => B(27), Ci => CTMP_27_port, S => 
                           S(27), Co => CTMP_28_port);
   FAI_29 : FA_804 port map( A => A(28), B => B(28), Ci => CTMP_28_port, S => 
                           S(28), Co => CTMP_29_port);
   FAI_30 : FA_803 port map( A => A(29), B => B(29), Ci => CTMP_29_port, S => 
                           S(29), Co => CTMP_30_port);
   FAI_31 : FA_802 port map( A => A(30), B => B(30), Ci => CTMP_30_port, S => 
                           S(30), Co => CTMP_31_port);
   FAI_32 : FA_801 port map( A => A(31), B => B(31), Ci => CTMP_31_port, S => 
                           S(31), Co => CTMP_32_port);
   FAI_33 : FA_800 port map( A => A(32), B => B(32), Ci => CTMP_32_port, S => 
                           S(32), Co => CTMP_33_port);
   FAI_34 : FA_799 port map( A => A(33), B => B(33), Ci => CTMP_33_port, S => 
                           S(33), Co => CTMP_34_port);
   FAI_35 : FA_798 port map( A => A(34), B => B(34), Ci => CTMP_34_port, S => 
                           S(34), Co => CTMP_35_port);
   FAI_36 : FA_797 port map( A => A(35), B => B(35), Ci => CTMP_35_port, S => 
                           S(35), Co => CTMP_36_port);
   FAI_37 : FA_796 port map( A => A(36), B => B(36), Ci => CTMP_36_port, S => 
                           S(36), Co => CTMP_37_port);
   FAI_38 : FA_795 port map( A => A(37), B => B(37), Ci => CTMP_37_port, S => 
                           S(37), Co => CTMP_38_port);
   FAI_39 : FA_794 port map( A => A(38), B => B(38), Ci => CTMP_38_port, S => 
                           S(38), Co => CTMP_39_port);
   FAI_40 : FA_793 port map( A => A(39), B => B(39), Ci => CTMP_39_port, S => 
                           S(39), Co => CTMP_40_port);
   FAI_41 : FA_792 port map( A => A(40), B => B(40), Ci => CTMP_40_port, S => 
                           S(40), Co => CTMP_41_port);
   FAI_42 : FA_791 port map( A => A(41), B => B(41), Ci => CTMP_41_port, S => 
                           S(41), Co => CTMP_42_port);
   FAI_43 : FA_790 port map( A => A(42), B => B(42), Ci => CTMP_42_port, S => 
                           S(42), Co => CTMP_43_port);
   FAI_44 : FA_789 port map( A => A(43), B => B(43), Ci => CTMP_43_port, S => 
                           S(43), Co => CTMP_44_port);
   FAI_45 : FA_788 port map( A => A(44), B => B(44), Ci => CTMP_44_port, S => 
                           S(44), Co => CTMP_45_port);
   FAI_46 : FA_787 port map( A => A(45), B => B(45), Ci => CTMP_45_port, S => 
                           S(45), Co => CTMP_46_port);
   FAI_47 : FA_786 port map( A => A(46), B => B(46), Ci => CTMP_46_port, S => 
                           S(46), Co => CTMP_47_port);
   FAI_48 : FA_785 port map( A => A(47), B => B(47), Ci => CTMP_47_port, S => 
                           S(47), Co => CTMP_48_port);
   FAI_49 : FA_784 port map( A => A(48), B => B(48), Ci => CTMP_48_port, S => 
                           S(48), Co => CTMP_49_port);
   FAI_50 : FA_783 port map( A => A(49), B => B(49), Ci => CTMP_49_port, S => 
                           S(49), Co => CTMP_50_port);
   FAI_51 : FA_782 port map( A => A(50), B => B(50), Ci => CTMP_50_port, S => 
                           S(50), Co => CTMP_51_port);
   FAI_52 : FA_781 port map( A => A(51), B => B(51), Ci => CTMP_51_port, S => 
                           S(51), Co => CTMP_52_port);
   FAI_53 : FA_780 port map( A => A(52), B => B(52), Ci => CTMP_52_port, S => 
                           S(52), Co => CTMP_53_port);
   FAI_54 : FA_779 port map( A => A(53), B => B(53), Ci => CTMP_53_port, S => 
                           S(53), Co => CTMP_54_port);
   FAI_55 : FA_778 port map( A => A(54), B => B(54), Ci => CTMP_54_port, S => 
                           S(54), Co => CTMP_55_port);
   FAI_56 : FA_777 port map( A => A(55), B => B(55), Ci => CTMP_55_port, S => 
                           S(55), Co => CTMP_56_port);
   FAI_57 : FA_776 port map( A => A(56), B => B(56), Ci => CTMP_56_port, S => 
                           S(56), Co => CTMP_57_port);
   FAI_58 : FA_775 port map( A => A(57), B => B(57), Ci => CTMP_57_port, S => 
                           S(57), Co => CTMP_58_port);
   FAI_59 : FA_774 port map( A => A(58), B => B(58), Ci => CTMP_58_port, S => 
                           S(58), Co => CTMP_59_port);
   FAI_60 : FA_773 port map( A => A(59), B => B(59), Ci => CTMP_59_port, S => 
                           S(59), Co => CTMP_60_port);
   FAI_61 : FA_772 port map( A => A(60), B => B(60), Ci => CTMP_60_port, S => 
                           S(60), Co => CTMP_61_port);
   FAI_62 : FA_771 port map( A => A(61), B => B(61), Ci => CTMP_61_port, S => 
                           S(61), Co => CTMP_62_port);
   FAI_63 : FA_770 port map( A => A(62), B => B(62), Ci => CTMP_62_port, S => 
                           S(62), Co => CTMP_63_port);
   FAI_64 : FA_769 port map( A => A(63), B => B(63), Ci => CTMP_63_port, S => 
                           S(63), Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity RCA_NbitRca64_12 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_NbitRca64_12;

architecture SYN_STRUCTURAL of RCA_NbitRca64_12 is

   component FA_705
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_706
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_707
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_708
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_709
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_710
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_711
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_712
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_713
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_714
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_715
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_716
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_717
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_718
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_719
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_720
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_721
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_722
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_723
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_724
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_725
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_726
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_727
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_728
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_729
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_730
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_731
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_732
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_733
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_734
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_735
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_736
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_737
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_738
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_739
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_740
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_741
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_742
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_743
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_744
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_745
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_746
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_747
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_748
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_749
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_750
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_751
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_752
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_753
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_754
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_755
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_756
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_757
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_758
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_759
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_760
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_761
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_762
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_763
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_764
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_765
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_766
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_767
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_768
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_63_port, CTMP_62_port, CTMP_61_port, CTMP_60_port, CTMP_59_port,
      CTMP_58_port, CTMP_57_port, CTMP_56_port, CTMP_55_port, CTMP_54_port, 
      CTMP_53_port, CTMP_52_port, CTMP_51_port, CTMP_50_port, CTMP_49_port, 
      CTMP_48_port, CTMP_47_port, CTMP_46_port, CTMP_45_port, CTMP_44_port, 
      CTMP_43_port, CTMP_42_port, CTMP_41_port, CTMP_40_port, CTMP_39_port, 
      CTMP_38_port, CTMP_37_port, CTMP_36_port, CTMP_35_port, CTMP_34_port, 
      CTMP_33_port, CTMP_32_port, CTMP_31_port, CTMP_30_port, CTMP_29_port, 
      CTMP_28_port, CTMP_27_port, CTMP_26_port, CTMP_25_port, CTMP_24_port, 
      CTMP_23_port, CTMP_22_port, CTMP_21_port, CTMP_20_port, CTMP_19_port, 
      CTMP_18_port, CTMP_17_port, CTMP_16_port, CTMP_15_port, CTMP_14_port, 
      CTMP_13_port, CTMP_12_port, CTMP_11_port, CTMP_10_port, CTMP_9_port, 
      CTMP_8_port, CTMP_7_port, CTMP_6_port, CTMP_5_port, CTMP_4_port, 
      CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_768 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_767 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_766 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_765 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => CTMP_4_port);
   FAI_5 : FA_764 port map( A => A(4), B => B(4), Ci => CTMP_4_port, S => S(4),
                           Co => CTMP_5_port);
   FAI_6 : FA_763 port map( A => A(5), B => B(5), Ci => CTMP_5_port, S => S(5),
                           Co => CTMP_6_port);
   FAI_7 : FA_762 port map( A => A(6), B => B(6), Ci => CTMP_6_port, S => S(6),
                           Co => CTMP_7_port);
   FAI_8 : FA_761 port map( A => A(7), B => B(7), Ci => CTMP_7_port, S => S(7),
                           Co => CTMP_8_port);
   FAI_9 : FA_760 port map( A => A(8), B => B(8), Ci => CTMP_8_port, S => S(8),
                           Co => CTMP_9_port);
   FAI_10 : FA_759 port map( A => A(9), B => B(9), Ci => CTMP_9_port, S => S(9)
                           , Co => CTMP_10_port);
   FAI_11 : FA_758 port map( A => A(10), B => B(10), Ci => CTMP_10_port, S => 
                           S(10), Co => CTMP_11_port);
   FAI_12 : FA_757 port map( A => A(11), B => B(11), Ci => CTMP_11_port, S => 
                           S(11), Co => CTMP_12_port);
   FAI_13 : FA_756 port map( A => A(12), B => B(12), Ci => CTMP_12_port, S => 
                           S(12), Co => CTMP_13_port);
   FAI_14 : FA_755 port map( A => A(13), B => B(13), Ci => CTMP_13_port, S => 
                           S(13), Co => CTMP_14_port);
   FAI_15 : FA_754 port map( A => A(14), B => B(14), Ci => CTMP_14_port, S => 
                           S(14), Co => CTMP_15_port);
   FAI_16 : FA_753 port map( A => A(15), B => B(15), Ci => CTMP_15_port, S => 
                           S(15), Co => CTMP_16_port);
   FAI_17 : FA_752 port map( A => A(16), B => B(16), Ci => CTMP_16_port, S => 
                           S(16), Co => CTMP_17_port);
   FAI_18 : FA_751 port map( A => A(17), B => B(17), Ci => CTMP_17_port, S => 
                           S(17), Co => CTMP_18_port);
   FAI_19 : FA_750 port map( A => A(18), B => B(18), Ci => CTMP_18_port, S => 
                           S(18), Co => CTMP_19_port);
   FAI_20 : FA_749 port map( A => A(19), B => B(19), Ci => CTMP_19_port, S => 
                           S(19), Co => CTMP_20_port);
   FAI_21 : FA_748 port map( A => A(20), B => B(20), Ci => CTMP_20_port, S => 
                           S(20), Co => CTMP_21_port);
   FAI_22 : FA_747 port map( A => A(21), B => B(21), Ci => CTMP_21_port, S => 
                           S(21), Co => CTMP_22_port);
   FAI_23 : FA_746 port map( A => A(22), B => B(22), Ci => CTMP_22_port, S => 
                           S(22), Co => CTMP_23_port);
   FAI_24 : FA_745 port map( A => A(23), B => B(23), Ci => CTMP_23_port, S => 
                           S(23), Co => CTMP_24_port);
   FAI_25 : FA_744 port map( A => A(24), B => B(24), Ci => CTMP_24_port, S => 
                           S(24), Co => CTMP_25_port);
   FAI_26 : FA_743 port map( A => A(25), B => B(25), Ci => CTMP_25_port, S => 
                           S(25), Co => CTMP_26_port);
   FAI_27 : FA_742 port map( A => A(26), B => B(26), Ci => CTMP_26_port, S => 
                           S(26), Co => CTMP_27_port);
   FAI_28 : FA_741 port map( A => A(27), B => B(27), Ci => CTMP_27_port, S => 
                           S(27), Co => CTMP_28_port);
   FAI_29 : FA_740 port map( A => A(28), B => B(28), Ci => CTMP_28_port, S => 
                           S(28), Co => CTMP_29_port);
   FAI_30 : FA_739 port map( A => A(29), B => B(29), Ci => CTMP_29_port, S => 
                           S(29), Co => CTMP_30_port);
   FAI_31 : FA_738 port map( A => A(30), B => B(30), Ci => CTMP_30_port, S => 
                           S(30), Co => CTMP_31_port);
   FAI_32 : FA_737 port map( A => A(31), B => B(31), Ci => CTMP_31_port, S => 
                           S(31), Co => CTMP_32_port);
   FAI_33 : FA_736 port map( A => A(32), B => B(32), Ci => CTMP_32_port, S => 
                           S(32), Co => CTMP_33_port);
   FAI_34 : FA_735 port map( A => A(33), B => B(33), Ci => CTMP_33_port, S => 
                           S(33), Co => CTMP_34_port);
   FAI_35 : FA_734 port map( A => A(34), B => B(34), Ci => CTMP_34_port, S => 
                           S(34), Co => CTMP_35_port);
   FAI_36 : FA_733 port map( A => A(35), B => B(35), Ci => CTMP_35_port, S => 
                           S(35), Co => CTMP_36_port);
   FAI_37 : FA_732 port map( A => A(36), B => B(36), Ci => CTMP_36_port, S => 
                           S(36), Co => CTMP_37_port);
   FAI_38 : FA_731 port map( A => A(37), B => B(37), Ci => CTMP_37_port, S => 
                           S(37), Co => CTMP_38_port);
   FAI_39 : FA_730 port map( A => A(38), B => B(38), Ci => CTMP_38_port, S => 
                           S(38), Co => CTMP_39_port);
   FAI_40 : FA_729 port map( A => A(39), B => B(39), Ci => CTMP_39_port, S => 
                           S(39), Co => CTMP_40_port);
   FAI_41 : FA_728 port map( A => A(40), B => B(40), Ci => CTMP_40_port, S => 
                           S(40), Co => CTMP_41_port);
   FAI_42 : FA_727 port map( A => A(41), B => B(41), Ci => CTMP_41_port, S => 
                           S(41), Co => CTMP_42_port);
   FAI_43 : FA_726 port map( A => A(42), B => B(42), Ci => CTMP_42_port, S => 
                           S(42), Co => CTMP_43_port);
   FAI_44 : FA_725 port map( A => A(43), B => B(43), Ci => CTMP_43_port, S => 
                           S(43), Co => CTMP_44_port);
   FAI_45 : FA_724 port map( A => A(44), B => B(44), Ci => CTMP_44_port, S => 
                           S(44), Co => CTMP_45_port);
   FAI_46 : FA_723 port map( A => A(45), B => B(45), Ci => CTMP_45_port, S => 
                           S(45), Co => CTMP_46_port);
   FAI_47 : FA_722 port map( A => A(46), B => B(46), Ci => CTMP_46_port, S => 
                           S(46), Co => CTMP_47_port);
   FAI_48 : FA_721 port map( A => A(47), B => B(47), Ci => CTMP_47_port, S => 
                           S(47), Co => CTMP_48_port);
   FAI_49 : FA_720 port map( A => A(48), B => B(48), Ci => CTMP_48_port, S => 
                           S(48), Co => CTMP_49_port);
   FAI_50 : FA_719 port map( A => A(49), B => B(49), Ci => CTMP_49_port, S => 
                           S(49), Co => CTMP_50_port);
   FAI_51 : FA_718 port map( A => A(50), B => B(50), Ci => CTMP_50_port, S => 
                           S(50), Co => CTMP_51_port);
   FAI_52 : FA_717 port map( A => A(51), B => B(51), Ci => CTMP_51_port, S => 
                           S(51), Co => CTMP_52_port);
   FAI_53 : FA_716 port map( A => A(52), B => B(52), Ci => CTMP_52_port, S => 
                           S(52), Co => CTMP_53_port);
   FAI_54 : FA_715 port map( A => A(53), B => B(53), Ci => CTMP_53_port, S => 
                           S(53), Co => CTMP_54_port);
   FAI_55 : FA_714 port map( A => A(54), B => B(54), Ci => CTMP_54_port, S => 
                           S(54), Co => CTMP_55_port);
   FAI_56 : FA_713 port map( A => A(55), B => B(55), Ci => CTMP_55_port, S => 
                           S(55), Co => CTMP_56_port);
   FAI_57 : FA_712 port map( A => A(56), B => B(56), Ci => CTMP_56_port, S => 
                           S(56), Co => CTMP_57_port);
   FAI_58 : FA_711 port map( A => A(57), B => B(57), Ci => CTMP_57_port, S => 
                           S(57), Co => CTMP_58_port);
   FAI_59 : FA_710 port map( A => A(58), B => B(58), Ci => CTMP_58_port, S => 
                           S(58), Co => CTMP_59_port);
   FAI_60 : FA_709 port map( A => A(59), B => B(59), Ci => CTMP_59_port, S => 
                           S(59), Co => CTMP_60_port);
   FAI_61 : FA_708 port map( A => A(60), B => B(60), Ci => CTMP_60_port, S => 
                           S(60), Co => CTMP_61_port);
   FAI_62 : FA_707 port map( A => A(61), B => B(61), Ci => CTMP_61_port, S => 
                           S(61), Co => CTMP_62_port);
   FAI_63 : FA_706 port map( A => A(62), B => B(62), Ci => CTMP_62_port, S => 
                           S(62), Co => CTMP_63_port);
   FAI_64 : FA_705 port map( A => A(63), B => B(63), Ci => CTMP_63_port, S => 
                           S(63), Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity RCA_NbitRca64_11 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_NbitRca64_11;

architecture SYN_STRUCTURAL of RCA_NbitRca64_11 is

   component FA_641
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_642
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_643
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_644
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_645
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_646
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_647
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_648
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_649
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_650
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_651
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_652
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_653
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_654
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_655
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_656
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_657
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_658
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_659
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_660
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_661
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_662
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_663
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_664
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_665
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_666
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_667
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_668
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_669
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_670
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_671
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_672
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_673
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_674
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_675
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_676
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_677
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_678
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_679
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_680
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_681
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_682
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_683
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_684
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_685
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_686
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_687
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_688
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_689
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_690
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_691
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_692
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_693
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_694
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_695
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_696
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_697
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_698
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_699
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_700
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_701
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_702
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_703
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_704
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_63_port, CTMP_62_port, CTMP_61_port, CTMP_60_port, CTMP_59_port,
      CTMP_58_port, CTMP_57_port, CTMP_56_port, CTMP_55_port, CTMP_54_port, 
      CTMP_53_port, CTMP_52_port, CTMP_51_port, CTMP_50_port, CTMP_49_port, 
      CTMP_48_port, CTMP_47_port, CTMP_46_port, CTMP_45_port, CTMP_44_port, 
      CTMP_43_port, CTMP_42_port, CTMP_41_port, CTMP_40_port, CTMP_39_port, 
      CTMP_38_port, CTMP_37_port, CTMP_36_port, CTMP_35_port, CTMP_34_port, 
      CTMP_33_port, CTMP_32_port, CTMP_31_port, CTMP_30_port, CTMP_29_port, 
      CTMP_28_port, CTMP_27_port, CTMP_26_port, CTMP_25_port, CTMP_24_port, 
      CTMP_23_port, CTMP_22_port, CTMP_21_port, CTMP_20_port, CTMP_19_port, 
      CTMP_18_port, CTMP_17_port, CTMP_16_port, CTMP_15_port, CTMP_14_port, 
      CTMP_13_port, CTMP_12_port, CTMP_11_port, CTMP_10_port, CTMP_9_port, 
      CTMP_8_port, CTMP_7_port, CTMP_6_port, CTMP_5_port, CTMP_4_port, 
      CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_704 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_703 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_702 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_701 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => CTMP_4_port);
   FAI_5 : FA_700 port map( A => A(4), B => B(4), Ci => CTMP_4_port, S => S(4),
                           Co => CTMP_5_port);
   FAI_6 : FA_699 port map( A => A(5), B => B(5), Ci => CTMP_5_port, S => S(5),
                           Co => CTMP_6_port);
   FAI_7 : FA_698 port map( A => A(6), B => B(6), Ci => CTMP_6_port, S => S(6),
                           Co => CTMP_7_port);
   FAI_8 : FA_697 port map( A => A(7), B => B(7), Ci => CTMP_7_port, S => S(7),
                           Co => CTMP_8_port);
   FAI_9 : FA_696 port map( A => A(8), B => B(8), Ci => CTMP_8_port, S => S(8),
                           Co => CTMP_9_port);
   FAI_10 : FA_695 port map( A => A(9), B => B(9), Ci => CTMP_9_port, S => S(9)
                           , Co => CTMP_10_port);
   FAI_11 : FA_694 port map( A => A(10), B => B(10), Ci => CTMP_10_port, S => 
                           S(10), Co => CTMP_11_port);
   FAI_12 : FA_693 port map( A => A(11), B => B(11), Ci => CTMP_11_port, S => 
                           S(11), Co => CTMP_12_port);
   FAI_13 : FA_692 port map( A => A(12), B => B(12), Ci => CTMP_12_port, S => 
                           S(12), Co => CTMP_13_port);
   FAI_14 : FA_691 port map( A => A(13), B => B(13), Ci => CTMP_13_port, S => 
                           S(13), Co => CTMP_14_port);
   FAI_15 : FA_690 port map( A => A(14), B => B(14), Ci => CTMP_14_port, S => 
                           S(14), Co => CTMP_15_port);
   FAI_16 : FA_689 port map( A => A(15), B => B(15), Ci => CTMP_15_port, S => 
                           S(15), Co => CTMP_16_port);
   FAI_17 : FA_688 port map( A => A(16), B => B(16), Ci => CTMP_16_port, S => 
                           S(16), Co => CTMP_17_port);
   FAI_18 : FA_687 port map( A => A(17), B => B(17), Ci => CTMP_17_port, S => 
                           S(17), Co => CTMP_18_port);
   FAI_19 : FA_686 port map( A => A(18), B => B(18), Ci => CTMP_18_port, S => 
                           S(18), Co => CTMP_19_port);
   FAI_20 : FA_685 port map( A => A(19), B => B(19), Ci => CTMP_19_port, S => 
                           S(19), Co => CTMP_20_port);
   FAI_21 : FA_684 port map( A => A(20), B => B(20), Ci => CTMP_20_port, S => 
                           S(20), Co => CTMP_21_port);
   FAI_22 : FA_683 port map( A => A(21), B => B(21), Ci => CTMP_21_port, S => 
                           S(21), Co => CTMP_22_port);
   FAI_23 : FA_682 port map( A => A(22), B => B(22), Ci => CTMP_22_port, S => 
                           S(22), Co => CTMP_23_port);
   FAI_24 : FA_681 port map( A => A(23), B => B(23), Ci => CTMP_23_port, S => 
                           S(23), Co => CTMP_24_port);
   FAI_25 : FA_680 port map( A => A(24), B => B(24), Ci => CTMP_24_port, S => 
                           S(24), Co => CTMP_25_port);
   FAI_26 : FA_679 port map( A => A(25), B => B(25), Ci => CTMP_25_port, S => 
                           S(25), Co => CTMP_26_port);
   FAI_27 : FA_678 port map( A => A(26), B => B(26), Ci => CTMP_26_port, S => 
                           S(26), Co => CTMP_27_port);
   FAI_28 : FA_677 port map( A => A(27), B => B(27), Ci => CTMP_27_port, S => 
                           S(27), Co => CTMP_28_port);
   FAI_29 : FA_676 port map( A => A(28), B => B(28), Ci => CTMP_28_port, S => 
                           S(28), Co => CTMP_29_port);
   FAI_30 : FA_675 port map( A => A(29), B => B(29), Ci => CTMP_29_port, S => 
                           S(29), Co => CTMP_30_port);
   FAI_31 : FA_674 port map( A => A(30), B => B(30), Ci => CTMP_30_port, S => 
                           S(30), Co => CTMP_31_port);
   FAI_32 : FA_673 port map( A => A(31), B => B(31), Ci => CTMP_31_port, S => 
                           S(31), Co => CTMP_32_port);
   FAI_33 : FA_672 port map( A => A(32), B => B(32), Ci => CTMP_32_port, S => 
                           S(32), Co => CTMP_33_port);
   FAI_34 : FA_671 port map( A => A(33), B => B(33), Ci => CTMP_33_port, S => 
                           S(33), Co => CTMP_34_port);
   FAI_35 : FA_670 port map( A => A(34), B => B(34), Ci => CTMP_34_port, S => 
                           S(34), Co => CTMP_35_port);
   FAI_36 : FA_669 port map( A => A(35), B => B(35), Ci => CTMP_35_port, S => 
                           S(35), Co => CTMP_36_port);
   FAI_37 : FA_668 port map( A => A(36), B => B(36), Ci => CTMP_36_port, S => 
                           S(36), Co => CTMP_37_port);
   FAI_38 : FA_667 port map( A => A(37), B => B(37), Ci => CTMP_37_port, S => 
                           S(37), Co => CTMP_38_port);
   FAI_39 : FA_666 port map( A => A(38), B => B(38), Ci => CTMP_38_port, S => 
                           S(38), Co => CTMP_39_port);
   FAI_40 : FA_665 port map( A => A(39), B => B(39), Ci => CTMP_39_port, S => 
                           S(39), Co => CTMP_40_port);
   FAI_41 : FA_664 port map( A => A(40), B => B(40), Ci => CTMP_40_port, S => 
                           S(40), Co => CTMP_41_port);
   FAI_42 : FA_663 port map( A => A(41), B => B(41), Ci => CTMP_41_port, S => 
                           S(41), Co => CTMP_42_port);
   FAI_43 : FA_662 port map( A => A(42), B => B(42), Ci => CTMP_42_port, S => 
                           S(42), Co => CTMP_43_port);
   FAI_44 : FA_661 port map( A => A(43), B => B(43), Ci => CTMP_43_port, S => 
                           S(43), Co => CTMP_44_port);
   FAI_45 : FA_660 port map( A => A(44), B => B(44), Ci => CTMP_44_port, S => 
                           S(44), Co => CTMP_45_port);
   FAI_46 : FA_659 port map( A => A(45), B => B(45), Ci => CTMP_45_port, S => 
                           S(45), Co => CTMP_46_port);
   FAI_47 : FA_658 port map( A => A(46), B => B(46), Ci => CTMP_46_port, S => 
                           S(46), Co => CTMP_47_port);
   FAI_48 : FA_657 port map( A => A(47), B => B(47), Ci => CTMP_47_port, S => 
                           S(47), Co => CTMP_48_port);
   FAI_49 : FA_656 port map( A => A(48), B => B(48), Ci => CTMP_48_port, S => 
                           S(48), Co => CTMP_49_port);
   FAI_50 : FA_655 port map( A => A(49), B => B(49), Ci => CTMP_49_port, S => 
                           S(49), Co => CTMP_50_port);
   FAI_51 : FA_654 port map( A => A(50), B => B(50), Ci => CTMP_50_port, S => 
                           S(50), Co => CTMP_51_port);
   FAI_52 : FA_653 port map( A => A(51), B => B(51), Ci => CTMP_51_port, S => 
                           S(51), Co => CTMP_52_port);
   FAI_53 : FA_652 port map( A => A(52), B => B(52), Ci => CTMP_52_port, S => 
                           S(52), Co => CTMP_53_port);
   FAI_54 : FA_651 port map( A => A(53), B => B(53), Ci => CTMP_53_port, S => 
                           S(53), Co => CTMP_54_port);
   FAI_55 : FA_650 port map( A => A(54), B => B(54), Ci => CTMP_54_port, S => 
                           S(54), Co => CTMP_55_port);
   FAI_56 : FA_649 port map( A => A(55), B => B(55), Ci => CTMP_55_port, S => 
                           S(55), Co => CTMP_56_port);
   FAI_57 : FA_648 port map( A => A(56), B => B(56), Ci => CTMP_56_port, S => 
                           S(56), Co => CTMP_57_port);
   FAI_58 : FA_647 port map( A => A(57), B => B(57), Ci => CTMP_57_port, S => 
                           S(57), Co => CTMP_58_port);
   FAI_59 : FA_646 port map( A => A(58), B => B(58), Ci => CTMP_58_port, S => 
                           S(58), Co => CTMP_59_port);
   FAI_60 : FA_645 port map( A => A(59), B => B(59), Ci => CTMP_59_port, S => 
                           S(59), Co => CTMP_60_port);
   FAI_61 : FA_644 port map( A => A(60), B => B(60), Ci => CTMP_60_port, S => 
                           S(60), Co => CTMP_61_port);
   FAI_62 : FA_643 port map( A => A(61), B => B(61), Ci => CTMP_61_port, S => 
                           S(61), Co => CTMP_62_port);
   FAI_63 : FA_642 port map( A => A(62), B => B(62), Ci => CTMP_62_port, S => 
                           S(62), Co => CTMP_63_port);
   FAI_64 : FA_641 port map( A => A(63), B => B(63), Ci => CTMP_63_port, S => 
                           S(63), Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity RCA_NbitRca64_10 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_NbitRca64_10;

architecture SYN_STRUCTURAL of RCA_NbitRca64_10 is

   component FA_577
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_578
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_579
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_580
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_581
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_582
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_583
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_584
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_585
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_586
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_587
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_588
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_589
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_590
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_591
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_592
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_593
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_594
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_595
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_596
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_597
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_598
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_599
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_600
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_601
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_602
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_603
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_604
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_605
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_606
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_607
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_608
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_609
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_610
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_611
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_612
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_613
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_614
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_615
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_616
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_617
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_618
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_619
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_620
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_621
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_622
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_623
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_624
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_625
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_626
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_627
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_628
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_629
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_630
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_631
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_632
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_633
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_634
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_635
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_636
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_637
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_638
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_639
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_640
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_63_port, CTMP_62_port, CTMP_61_port, CTMP_60_port, CTMP_59_port,
      CTMP_58_port, CTMP_57_port, CTMP_56_port, CTMP_55_port, CTMP_54_port, 
      CTMP_53_port, CTMP_52_port, CTMP_51_port, CTMP_50_port, CTMP_49_port, 
      CTMP_48_port, CTMP_47_port, CTMP_46_port, CTMP_45_port, CTMP_44_port, 
      CTMP_43_port, CTMP_42_port, CTMP_41_port, CTMP_40_port, CTMP_39_port, 
      CTMP_38_port, CTMP_37_port, CTMP_36_port, CTMP_35_port, CTMP_34_port, 
      CTMP_33_port, CTMP_32_port, CTMP_31_port, CTMP_30_port, CTMP_29_port, 
      CTMP_28_port, CTMP_27_port, CTMP_26_port, CTMP_25_port, CTMP_24_port, 
      CTMP_23_port, CTMP_22_port, CTMP_21_port, CTMP_20_port, CTMP_19_port, 
      CTMP_18_port, CTMP_17_port, CTMP_16_port, CTMP_15_port, CTMP_14_port, 
      CTMP_13_port, CTMP_12_port, CTMP_11_port, CTMP_10_port, CTMP_9_port, 
      CTMP_8_port, CTMP_7_port, CTMP_6_port, CTMP_5_port, CTMP_4_port, 
      CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_640 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_639 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_638 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_637 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => CTMP_4_port);
   FAI_5 : FA_636 port map( A => A(4), B => B(4), Ci => CTMP_4_port, S => S(4),
                           Co => CTMP_5_port);
   FAI_6 : FA_635 port map( A => A(5), B => B(5), Ci => CTMP_5_port, S => S(5),
                           Co => CTMP_6_port);
   FAI_7 : FA_634 port map( A => A(6), B => B(6), Ci => CTMP_6_port, S => S(6),
                           Co => CTMP_7_port);
   FAI_8 : FA_633 port map( A => A(7), B => B(7), Ci => CTMP_7_port, S => S(7),
                           Co => CTMP_8_port);
   FAI_9 : FA_632 port map( A => A(8), B => B(8), Ci => CTMP_8_port, S => S(8),
                           Co => CTMP_9_port);
   FAI_10 : FA_631 port map( A => A(9), B => B(9), Ci => CTMP_9_port, S => S(9)
                           , Co => CTMP_10_port);
   FAI_11 : FA_630 port map( A => A(10), B => B(10), Ci => CTMP_10_port, S => 
                           S(10), Co => CTMP_11_port);
   FAI_12 : FA_629 port map( A => A(11), B => B(11), Ci => CTMP_11_port, S => 
                           S(11), Co => CTMP_12_port);
   FAI_13 : FA_628 port map( A => A(12), B => B(12), Ci => CTMP_12_port, S => 
                           S(12), Co => CTMP_13_port);
   FAI_14 : FA_627 port map( A => A(13), B => B(13), Ci => CTMP_13_port, S => 
                           S(13), Co => CTMP_14_port);
   FAI_15 : FA_626 port map( A => A(14), B => B(14), Ci => CTMP_14_port, S => 
                           S(14), Co => CTMP_15_port);
   FAI_16 : FA_625 port map( A => A(15), B => B(15), Ci => CTMP_15_port, S => 
                           S(15), Co => CTMP_16_port);
   FAI_17 : FA_624 port map( A => A(16), B => B(16), Ci => CTMP_16_port, S => 
                           S(16), Co => CTMP_17_port);
   FAI_18 : FA_623 port map( A => A(17), B => B(17), Ci => CTMP_17_port, S => 
                           S(17), Co => CTMP_18_port);
   FAI_19 : FA_622 port map( A => A(18), B => B(18), Ci => CTMP_18_port, S => 
                           S(18), Co => CTMP_19_port);
   FAI_20 : FA_621 port map( A => A(19), B => B(19), Ci => CTMP_19_port, S => 
                           S(19), Co => CTMP_20_port);
   FAI_21 : FA_620 port map( A => A(20), B => B(20), Ci => CTMP_20_port, S => 
                           S(20), Co => CTMP_21_port);
   FAI_22 : FA_619 port map( A => A(21), B => B(21), Ci => CTMP_21_port, S => 
                           S(21), Co => CTMP_22_port);
   FAI_23 : FA_618 port map( A => A(22), B => B(22), Ci => CTMP_22_port, S => 
                           S(22), Co => CTMP_23_port);
   FAI_24 : FA_617 port map( A => A(23), B => B(23), Ci => CTMP_23_port, S => 
                           S(23), Co => CTMP_24_port);
   FAI_25 : FA_616 port map( A => A(24), B => B(24), Ci => CTMP_24_port, S => 
                           S(24), Co => CTMP_25_port);
   FAI_26 : FA_615 port map( A => A(25), B => B(25), Ci => CTMP_25_port, S => 
                           S(25), Co => CTMP_26_port);
   FAI_27 : FA_614 port map( A => A(26), B => B(26), Ci => CTMP_26_port, S => 
                           S(26), Co => CTMP_27_port);
   FAI_28 : FA_613 port map( A => A(27), B => B(27), Ci => CTMP_27_port, S => 
                           S(27), Co => CTMP_28_port);
   FAI_29 : FA_612 port map( A => A(28), B => B(28), Ci => CTMP_28_port, S => 
                           S(28), Co => CTMP_29_port);
   FAI_30 : FA_611 port map( A => A(29), B => B(29), Ci => CTMP_29_port, S => 
                           S(29), Co => CTMP_30_port);
   FAI_31 : FA_610 port map( A => A(30), B => B(30), Ci => CTMP_30_port, S => 
                           S(30), Co => CTMP_31_port);
   FAI_32 : FA_609 port map( A => A(31), B => B(31), Ci => CTMP_31_port, S => 
                           S(31), Co => CTMP_32_port);
   FAI_33 : FA_608 port map( A => A(32), B => B(32), Ci => CTMP_32_port, S => 
                           S(32), Co => CTMP_33_port);
   FAI_34 : FA_607 port map( A => A(33), B => B(33), Ci => CTMP_33_port, S => 
                           S(33), Co => CTMP_34_port);
   FAI_35 : FA_606 port map( A => A(34), B => B(34), Ci => CTMP_34_port, S => 
                           S(34), Co => CTMP_35_port);
   FAI_36 : FA_605 port map( A => A(35), B => B(35), Ci => CTMP_35_port, S => 
                           S(35), Co => CTMP_36_port);
   FAI_37 : FA_604 port map( A => A(36), B => B(36), Ci => CTMP_36_port, S => 
                           S(36), Co => CTMP_37_port);
   FAI_38 : FA_603 port map( A => A(37), B => B(37), Ci => CTMP_37_port, S => 
                           S(37), Co => CTMP_38_port);
   FAI_39 : FA_602 port map( A => A(38), B => B(38), Ci => CTMP_38_port, S => 
                           S(38), Co => CTMP_39_port);
   FAI_40 : FA_601 port map( A => A(39), B => B(39), Ci => CTMP_39_port, S => 
                           S(39), Co => CTMP_40_port);
   FAI_41 : FA_600 port map( A => A(40), B => B(40), Ci => CTMP_40_port, S => 
                           S(40), Co => CTMP_41_port);
   FAI_42 : FA_599 port map( A => A(41), B => B(41), Ci => CTMP_41_port, S => 
                           S(41), Co => CTMP_42_port);
   FAI_43 : FA_598 port map( A => A(42), B => B(42), Ci => CTMP_42_port, S => 
                           S(42), Co => CTMP_43_port);
   FAI_44 : FA_597 port map( A => A(43), B => B(43), Ci => CTMP_43_port, S => 
                           S(43), Co => CTMP_44_port);
   FAI_45 : FA_596 port map( A => A(44), B => B(44), Ci => CTMP_44_port, S => 
                           S(44), Co => CTMP_45_port);
   FAI_46 : FA_595 port map( A => A(45), B => B(45), Ci => CTMP_45_port, S => 
                           S(45), Co => CTMP_46_port);
   FAI_47 : FA_594 port map( A => A(46), B => B(46), Ci => CTMP_46_port, S => 
                           S(46), Co => CTMP_47_port);
   FAI_48 : FA_593 port map( A => A(47), B => B(47), Ci => CTMP_47_port, S => 
                           S(47), Co => CTMP_48_port);
   FAI_49 : FA_592 port map( A => A(48), B => B(48), Ci => CTMP_48_port, S => 
                           S(48), Co => CTMP_49_port);
   FAI_50 : FA_591 port map( A => A(49), B => B(49), Ci => CTMP_49_port, S => 
                           S(49), Co => CTMP_50_port);
   FAI_51 : FA_590 port map( A => A(50), B => B(50), Ci => CTMP_50_port, S => 
                           S(50), Co => CTMP_51_port);
   FAI_52 : FA_589 port map( A => A(51), B => B(51), Ci => CTMP_51_port, S => 
                           S(51), Co => CTMP_52_port);
   FAI_53 : FA_588 port map( A => A(52), B => B(52), Ci => CTMP_52_port, S => 
                           S(52), Co => CTMP_53_port);
   FAI_54 : FA_587 port map( A => A(53), B => B(53), Ci => CTMP_53_port, S => 
                           S(53), Co => CTMP_54_port);
   FAI_55 : FA_586 port map( A => A(54), B => B(54), Ci => CTMP_54_port, S => 
                           S(54), Co => CTMP_55_port);
   FAI_56 : FA_585 port map( A => A(55), B => B(55), Ci => CTMP_55_port, S => 
                           S(55), Co => CTMP_56_port);
   FAI_57 : FA_584 port map( A => A(56), B => B(56), Ci => CTMP_56_port, S => 
                           S(56), Co => CTMP_57_port);
   FAI_58 : FA_583 port map( A => A(57), B => B(57), Ci => CTMP_57_port, S => 
                           S(57), Co => CTMP_58_port);
   FAI_59 : FA_582 port map( A => A(58), B => B(58), Ci => CTMP_58_port, S => 
                           S(58), Co => CTMP_59_port);
   FAI_60 : FA_581 port map( A => A(59), B => B(59), Ci => CTMP_59_port, S => 
                           S(59), Co => CTMP_60_port);
   FAI_61 : FA_580 port map( A => A(60), B => B(60), Ci => CTMP_60_port, S => 
                           S(60), Co => CTMP_61_port);
   FAI_62 : FA_579 port map( A => A(61), B => B(61), Ci => CTMP_61_port, S => 
                           S(61), Co => CTMP_62_port);
   FAI_63 : FA_578 port map( A => A(62), B => B(62), Ci => CTMP_62_port, S => 
                           S(62), Co => CTMP_63_port);
   FAI_64 : FA_577 port map( A => A(63), B => B(63), Ci => CTMP_63_port, S => 
                           S(63), Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity RCA_NbitRca64_9 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_NbitRca64_9;

architecture SYN_STRUCTURAL of RCA_NbitRca64_9 is

   component FA_513
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_514
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_515
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_516
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_517
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_518
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_519
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_520
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_521
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_522
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_523
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_524
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_525
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_526
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_527
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_528
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_529
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_530
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_531
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_532
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_533
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_534
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_535
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_536
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_537
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_538
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_539
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_540
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_541
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_542
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_543
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_544
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_545
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_546
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_547
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_548
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_549
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_550
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_551
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_552
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_553
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_554
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_555
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_556
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_557
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_558
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_559
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_560
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_561
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_562
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_563
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_564
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_565
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_566
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_567
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_568
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_569
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_570
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_571
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_572
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_573
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_574
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_575
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_576
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_63_port, CTMP_62_port, CTMP_61_port, CTMP_60_port, CTMP_59_port,
      CTMP_58_port, CTMP_57_port, CTMP_56_port, CTMP_55_port, CTMP_54_port, 
      CTMP_53_port, CTMP_52_port, CTMP_51_port, CTMP_50_port, CTMP_49_port, 
      CTMP_48_port, CTMP_47_port, CTMP_46_port, CTMP_45_port, CTMP_44_port, 
      CTMP_43_port, CTMP_42_port, CTMP_41_port, CTMP_40_port, CTMP_39_port, 
      CTMP_38_port, CTMP_37_port, CTMP_36_port, CTMP_35_port, CTMP_34_port, 
      CTMP_33_port, CTMP_32_port, CTMP_31_port, CTMP_30_port, CTMP_29_port, 
      CTMP_28_port, CTMP_27_port, CTMP_26_port, CTMP_25_port, CTMP_24_port, 
      CTMP_23_port, CTMP_22_port, CTMP_21_port, CTMP_20_port, CTMP_19_port, 
      CTMP_18_port, CTMP_17_port, CTMP_16_port, CTMP_15_port, CTMP_14_port, 
      CTMP_13_port, CTMP_12_port, CTMP_11_port, CTMP_10_port, CTMP_9_port, 
      CTMP_8_port, CTMP_7_port, CTMP_6_port, CTMP_5_port, CTMP_4_port, 
      CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_576 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_575 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_574 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_573 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => CTMP_4_port);
   FAI_5 : FA_572 port map( A => A(4), B => B(4), Ci => CTMP_4_port, S => S(4),
                           Co => CTMP_5_port);
   FAI_6 : FA_571 port map( A => A(5), B => B(5), Ci => CTMP_5_port, S => S(5),
                           Co => CTMP_6_port);
   FAI_7 : FA_570 port map( A => A(6), B => B(6), Ci => CTMP_6_port, S => S(6),
                           Co => CTMP_7_port);
   FAI_8 : FA_569 port map( A => A(7), B => B(7), Ci => CTMP_7_port, S => S(7),
                           Co => CTMP_8_port);
   FAI_9 : FA_568 port map( A => A(8), B => B(8), Ci => CTMP_8_port, S => S(8),
                           Co => CTMP_9_port);
   FAI_10 : FA_567 port map( A => A(9), B => B(9), Ci => CTMP_9_port, S => S(9)
                           , Co => CTMP_10_port);
   FAI_11 : FA_566 port map( A => A(10), B => B(10), Ci => CTMP_10_port, S => 
                           S(10), Co => CTMP_11_port);
   FAI_12 : FA_565 port map( A => A(11), B => B(11), Ci => CTMP_11_port, S => 
                           S(11), Co => CTMP_12_port);
   FAI_13 : FA_564 port map( A => A(12), B => B(12), Ci => CTMP_12_port, S => 
                           S(12), Co => CTMP_13_port);
   FAI_14 : FA_563 port map( A => A(13), B => B(13), Ci => CTMP_13_port, S => 
                           S(13), Co => CTMP_14_port);
   FAI_15 : FA_562 port map( A => A(14), B => B(14), Ci => CTMP_14_port, S => 
                           S(14), Co => CTMP_15_port);
   FAI_16 : FA_561 port map( A => A(15), B => B(15), Ci => CTMP_15_port, S => 
                           S(15), Co => CTMP_16_port);
   FAI_17 : FA_560 port map( A => A(16), B => B(16), Ci => CTMP_16_port, S => 
                           S(16), Co => CTMP_17_port);
   FAI_18 : FA_559 port map( A => A(17), B => B(17), Ci => CTMP_17_port, S => 
                           S(17), Co => CTMP_18_port);
   FAI_19 : FA_558 port map( A => A(18), B => B(18), Ci => CTMP_18_port, S => 
                           S(18), Co => CTMP_19_port);
   FAI_20 : FA_557 port map( A => A(19), B => B(19), Ci => CTMP_19_port, S => 
                           S(19), Co => CTMP_20_port);
   FAI_21 : FA_556 port map( A => A(20), B => B(20), Ci => CTMP_20_port, S => 
                           S(20), Co => CTMP_21_port);
   FAI_22 : FA_555 port map( A => A(21), B => B(21), Ci => CTMP_21_port, S => 
                           S(21), Co => CTMP_22_port);
   FAI_23 : FA_554 port map( A => A(22), B => B(22), Ci => CTMP_22_port, S => 
                           S(22), Co => CTMP_23_port);
   FAI_24 : FA_553 port map( A => A(23), B => B(23), Ci => CTMP_23_port, S => 
                           S(23), Co => CTMP_24_port);
   FAI_25 : FA_552 port map( A => A(24), B => B(24), Ci => CTMP_24_port, S => 
                           S(24), Co => CTMP_25_port);
   FAI_26 : FA_551 port map( A => A(25), B => B(25), Ci => CTMP_25_port, S => 
                           S(25), Co => CTMP_26_port);
   FAI_27 : FA_550 port map( A => A(26), B => B(26), Ci => CTMP_26_port, S => 
                           S(26), Co => CTMP_27_port);
   FAI_28 : FA_549 port map( A => A(27), B => B(27), Ci => CTMP_27_port, S => 
                           S(27), Co => CTMP_28_port);
   FAI_29 : FA_548 port map( A => A(28), B => B(28), Ci => CTMP_28_port, S => 
                           S(28), Co => CTMP_29_port);
   FAI_30 : FA_547 port map( A => A(29), B => B(29), Ci => CTMP_29_port, S => 
                           S(29), Co => CTMP_30_port);
   FAI_31 : FA_546 port map( A => A(30), B => B(30), Ci => CTMP_30_port, S => 
                           S(30), Co => CTMP_31_port);
   FAI_32 : FA_545 port map( A => A(31), B => B(31), Ci => CTMP_31_port, S => 
                           S(31), Co => CTMP_32_port);
   FAI_33 : FA_544 port map( A => A(32), B => B(32), Ci => CTMP_32_port, S => 
                           S(32), Co => CTMP_33_port);
   FAI_34 : FA_543 port map( A => A(33), B => B(33), Ci => CTMP_33_port, S => 
                           S(33), Co => CTMP_34_port);
   FAI_35 : FA_542 port map( A => A(34), B => B(34), Ci => CTMP_34_port, S => 
                           S(34), Co => CTMP_35_port);
   FAI_36 : FA_541 port map( A => A(35), B => B(35), Ci => CTMP_35_port, S => 
                           S(35), Co => CTMP_36_port);
   FAI_37 : FA_540 port map( A => A(36), B => B(36), Ci => CTMP_36_port, S => 
                           S(36), Co => CTMP_37_port);
   FAI_38 : FA_539 port map( A => A(37), B => B(37), Ci => CTMP_37_port, S => 
                           S(37), Co => CTMP_38_port);
   FAI_39 : FA_538 port map( A => A(38), B => B(38), Ci => CTMP_38_port, S => 
                           S(38), Co => CTMP_39_port);
   FAI_40 : FA_537 port map( A => A(39), B => B(39), Ci => CTMP_39_port, S => 
                           S(39), Co => CTMP_40_port);
   FAI_41 : FA_536 port map( A => A(40), B => B(40), Ci => CTMP_40_port, S => 
                           S(40), Co => CTMP_41_port);
   FAI_42 : FA_535 port map( A => A(41), B => B(41), Ci => CTMP_41_port, S => 
                           S(41), Co => CTMP_42_port);
   FAI_43 : FA_534 port map( A => A(42), B => B(42), Ci => CTMP_42_port, S => 
                           S(42), Co => CTMP_43_port);
   FAI_44 : FA_533 port map( A => A(43), B => B(43), Ci => CTMP_43_port, S => 
                           S(43), Co => CTMP_44_port);
   FAI_45 : FA_532 port map( A => A(44), B => B(44), Ci => CTMP_44_port, S => 
                           S(44), Co => CTMP_45_port);
   FAI_46 : FA_531 port map( A => A(45), B => B(45), Ci => CTMP_45_port, S => 
                           S(45), Co => CTMP_46_port);
   FAI_47 : FA_530 port map( A => A(46), B => B(46), Ci => CTMP_46_port, S => 
                           S(46), Co => CTMP_47_port);
   FAI_48 : FA_529 port map( A => A(47), B => B(47), Ci => CTMP_47_port, S => 
                           S(47), Co => CTMP_48_port);
   FAI_49 : FA_528 port map( A => A(48), B => B(48), Ci => CTMP_48_port, S => 
                           S(48), Co => CTMP_49_port);
   FAI_50 : FA_527 port map( A => A(49), B => B(49), Ci => CTMP_49_port, S => 
                           S(49), Co => CTMP_50_port);
   FAI_51 : FA_526 port map( A => A(50), B => B(50), Ci => CTMP_50_port, S => 
                           S(50), Co => CTMP_51_port);
   FAI_52 : FA_525 port map( A => A(51), B => B(51), Ci => CTMP_51_port, S => 
                           S(51), Co => CTMP_52_port);
   FAI_53 : FA_524 port map( A => A(52), B => B(52), Ci => CTMP_52_port, S => 
                           S(52), Co => CTMP_53_port);
   FAI_54 : FA_523 port map( A => A(53), B => B(53), Ci => CTMP_53_port, S => 
                           S(53), Co => CTMP_54_port);
   FAI_55 : FA_522 port map( A => A(54), B => B(54), Ci => CTMP_54_port, S => 
                           S(54), Co => CTMP_55_port);
   FAI_56 : FA_521 port map( A => A(55), B => B(55), Ci => CTMP_55_port, S => 
                           S(55), Co => CTMP_56_port);
   FAI_57 : FA_520 port map( A => A(56), B => B(56), Ci => CTMP_56_port, S => 
                           S(56), Co => CTMP_57_port);
   FAI_58 : FA_519 port map( A => A(57), B => B(57), Ci => CTMP_57_port, S => 
                           S(57), Co => CTMP_58_port);
   FAI_59 : FA_518 port map( A => A(58), B => B(58), Ci => CTMP_58_port, S => 
                           S(58), Co => CTMP_59_port);
   FAI_60 : FA_517 port map( A => A(59), B => B(59), Ci => CTMP_59_port, S => 
                           S(59), Co => CTMP_60_port);
   FAI_61 : FA_516 port map( A => A(60), B => B(60), Ci => CTMP_60_port, S => 
                           S(60), Co => CTMP_61_port);
   FAI_62 : FA_515 port map( A => A(61), B => B(61), Ci => CTMP_61_port, S => 
                           S(61), Co => CTMP_62_port);
   FAI_63 : FA_514 port map( A => A(62), B => B(62), Ci => CTMP_62_port, S => 
                           S(62), Co => CTMP_63_port);
   FAI_64 : FA_513 port map( A => A(63), B => B(63), Ci => CTMP_63_port, S => 
                           S(63), Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity RCA_NbitRca64_8 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_NbitRca64_8;

architecture SYN_STRUCTURAL of RCA_NbitRca64_8 is

   component FA_449
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_450
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_451
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_452
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_453
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_454
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_455
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_456
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_457
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_458
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_459
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_460
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_461
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_462
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_463
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_464
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_465
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_466
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_467
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_468
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_469
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_470
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_471
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_472
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_473
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_474
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_475
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_476
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_477
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_478
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_479
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_480
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_481
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_482
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_483
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_484
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_485
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_486
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_487
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_488
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_489
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_490
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_491
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_492
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_493
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_494
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_495
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_496
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_497
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_498
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_499
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_500
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_501
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_502
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_503
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_504
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_505
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_506
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_507
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_508
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_509
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_510
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_511
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_512
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_63_port, CTMP_62_port, CTMP_61_port, CTMP_60_port, CTMP_59_port,
      CTMP_58_port, CTMP_57_port, CTMP_56_port, CTMP_55_port, CTMP_54_port, 
      CTMP_53_port, CTMP_52_port, CTMP_51_port, CTMP_50_port, CTMP_49_port, 
      CTMP_48_port, CTMP_47_port, CTMP_46_port, CTMP_45_port, CTMP_44_port, 
      CTMP_43_port, CTMP_42_port, CTMP_41_port, CTMP_40_port, CTMP_39_port, 
      CTMP_38_port, CTMP_37_port, CTMP_36_port, CTMP_35_port, CTMP_34_port, 
      CTMP_33_port, CTMP_32_port, CTMP_31_port, CTMP_30_port, CTMP_29_port, 
      CTMP_28_port, CTMP_27_port, CTMP_26_port, CTMP_25_port, CTMP_24_port, 
      CTMP_23_port, CTMP_22_port, CTMP_21_port, CTMP_20_port, CTMP_19_port, 
      CTMP_18_port, CTMP_17_port, CTMP_16_port, CTMP_15_port, CTMP_14_port, 
      CTMP_13_port, CTMP_12_port, CTMP_11_port, CTMP_10_port, CTMP_9_port, 
      CTMP_8_port, CTMP_7_port, CTMP_6_port, CTMP_5_port, CTMP_4_port, 
      CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_512 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_511 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_510 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_509 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => CTMP_4_port);
   FAI_5 : FA_508 port map( A => A(4), B => B(4), Ci => CTMP_4_port, S => S(4),
                           Co => CTMP_5_port);
   FAI_6 : FA_507 port map( A => A(5), B => B(5), Ci => CTMP_5_port, S => S(5),
                           Co => CTMP_6_port);
   FAI_7 : FA_506 port map( A => A(6), B => B(6), Ci => CTMP_6_port, S => S(6),
                           Co => CTMP_7_port);
   FAI_8 : FA_505 port map( A => A(7), B => B(7), Ci => CTMP_7_port, S => S(7),
                           Co => CTMP_8_port);
   FAI_9 : FA_504 port map( A => A(8), B => B(8), Ci => CTMP_8_port, S => S(8),
                           Co => CTMP_9_port);
   FAI_10 : FA_503 port map( A => A(9), B => B(9), Ci => CTMP_9_port, S => S(9)
                           , Co => CTMP_10_port);
   FAI_11 : FA_502 port map( A => A(10), B => B(10), Ci => CTMP_10_port, S => 
                           S(10), Co => CTMP_11_port);
   FAI_12 : FA_501 port map( A => A(11), B => B(11), Ci => CTMP_11_port, S => 
                           S(11), Co => CTMP_12_port);
   FAI_13 : FA_500 port map( A => A(12), B => B(12), Ci => CTMP_12_port, S => 
                           S(12), Co => CTMP_13_port);
   FAI_14 : FA_499 port map( A => A(13), B => B(13), Ci => CTMP_13_port, S => 
                           S(13), Co => CTMP_14_port);
   FAI_15 : FA_498 port map( A => A(14), B => B(14), Ci => CTMP_14_port, S => 
                           S(14), Co => CTMP_15_port);
   FAI_16 : FA_497 port map( A => A(15), B => B(15), Ci => CTMP_15_port, S => 
                           S(15), Co => CTMP_16_port);
   FAI_17 : FA_496 port map( A => A(16), B => B(16), Ci => CTMP_16_port, S => 
                           S(16), Co => CTMP_17_port);
   FAI_18 : FA_495 port map( A => A(17), B => B(17), Ci => CTMP_17_port, S => 
                           S(17), Co => CTMP_18_port);
   FAI_19 : FA_494 port map( A => A(18), B => B(18), Ci => CTMP_18_port, S => 
                           S(18), Co => CTMP_19_port);
   FAI_20 : FA_493 port map( A => A(19), B => B(19), Ci => CTMP_19_port, S => 
                           S(19), Co => CTMP_20_port);
   FAI_21 : FA_492 port map( A => A(20), B => B(20), Ci => CTMP_20_port, S => 
                           S(20), Co => CTMP_21_port);
   FAI_22 : FA_491 port map( A => A(21), B => B(21), Ci => CTMP_21_port, S => 
                           S(21), Co => CTMP_22_port);
   FAI_23 : FA_490 port map( A => A(22), B => B(22), Ci => CTMP_22_port, S => 
                           S(22), Co => CTMP_23_port);
   FAI_24 : FA_489 port map( A => A(23), B => B(23), Ci => CTMP_23_port, S => 
                           S(23), Co => CTMP_24_port);
   FAI_25 : FA_488 port map( A => A(24), B => B(24), Ci => CTMP_24_port, S => 
                           S(24), Co => CTMP_25_port);
   FAI_26 : FA_487 port map( A => A(25), B => B(25), Ci => CTMP_25_port, S => 
                           S(25), Co => CTMP_26_port);
   FAI_27 : FA_486 port map( A => A(26), B => B(26), Ci => CTMP_26_port, S => 
                           S(26), Co => CTMP_27_port);
   FAI_28 : FA_485 port map( A => A(27), B => B(27), Ci => CTMP_27_port, S => 
                           S(27), Co => CTMP_28_port);
   FAI_29 : FA_484 port map( A => A(28), B => B(28), Ci => CTMP_28_port, S => 
                           S(28), Co => CTMP_29_port);
   FAI_30 : FA_483 port map( A => A(29), B => B(29), Ci => CTMP_29_port, S => 
                           S(29), Co => CTMP_30_port);
   FAI_31 : FA_482 port map( A => A(30), B => B(30), Ci => CTMP_30_port, S => 
                           S(30), Co => CTMP_31_port);
   FAI_32 : FA_481 port map( A => A(31), B => B(31), Ci => CTMP_31_port, S => 
                           S(31), Co => CTMP_32_port);
   FAI_33 : FA_480 port map( A => A(32), B => B(32), Ci => CTMP_32_port, S => 
                           S(32), Co => CTMP_33_port);
   FAI_34 : FA_479 port map( A => A(33), B => B(33), Ci => CTMP_33_port, S => 
                           S(33), Co => CTMP_34_port);
   FAI_35 : FA_478 port map( A => A(34), B => B(34), Ci => CTMP_34_port, S => 
                           S(34), Co => CTMP_35_port);
   FAI_36 : FA_477 port map( A => A(35), B => B(35), Ci => CTMP_35_port, S => 
                           S(35), Co => CTMP_36_port);
   FAI_37 : FA_476 port map( A => A(36), B => B(36), Ci => CTMP_36_port, S => 
                           S(36), Co => CTMP_37_port);
   FAI_38 : FA_475 port map( A => A(37), B => B(37), Ci => CTMP_37_port, S => 
                           S(37), Co => CTMP_38_port);
   FAI_39 : FA_474 port map( A => A(38), B => B(38), Ci => CTMP_38_port, S => 
                           S(38), Co => CTMP_39_port);
   FAI_40 : FA_473 port map( A => A(39), B => B(39), Ci => CTMP_39_port, S => 
                           S(39), Co => CTMP_40_port);
   FAI_41 : FA_472 port map( A => A(40), B => B(40), Ci => CTMP_40_port, S => 
                           S(40), Co => CTMP_41_port);
   FAI_42 : FA_471 port map( A => A(41), B => B(41), Ci => CTMP_41_port, S => 
                           S(41), Co => CTMP_42_port);
   FAI_43 : FA_470 port map( A => A(42), B => B(42), Ci => CTMP_42_port, S => 
                           S(42), Co => CTMP_43_port);
   FAI_44 : FA_469 port map( A => A(43), B => B(43), Ci => CTMP_43_port, S => 
                           S(43), Co => CTMP_44_port);
   FAI_45 : FA_468 port map( A => A(44), B => B(44), Ci => CTMP_44_port, S => 
                           S(44), Co => CTMP_45_port);
   FAI_46 : FA_467 port map( A => A(45), B => B(45), Ci => CTMP_45_port, S => 
                           S(45), Co => CTMP_46_port);
   FAI_47 : FA_466 port map( A => A(46), B => B(46), Ci => CTMP_46_port, S => 
                           S(46), Co => CTMP_47_port);
   FAI_48 : FA_465 port map( A => A(47), B => B(47), Ci => CTMP_47_port, S => 
                           S(47), Co => CTMP_48_port);
   FAI_49 : FA_464 port map( A => A(48), B => B(48), Ci => CTMP_48_port, S => 
                           S(48), Co => CTMP_49_port);
   FAI_50 : FA_463 port map( A => A(49), B => B(49), Ci => CTMP_49_port, S => 
                           S(49), Co => CTMP_50_port);
   FAI_51 : FA_462 port map( A => A(50), B => B(50), Ci => CTMP_50_port, S => 
                           S(50), Co => CTMP_51_port);
   FAI_52 : FA_461 port map( A => A(51), B => B(51), Ci => CTMP_51_port, S => 
                           S(51), Co => CTMP_52_port);
   FAI_53 : FA_460 port map( A => A(52), B => B(52), Ci => CTMP_52_port, S => 
                           S(52), Co => CTMP_53_port);
   FAI_54 : FA_459 port map( A => A(53), B => B(53), Ci => CTMP_53_port, S => 
                           S(53), Co => CTMP_54_port);
   FAI_55 : FA_458 port map( A => A(54), B => B(54), Ci => CTMP_54_port, S => 
                           S(54), Co => CTMP_55_port);
   FAI_56 : FA_457 port map( A => A(55), B => B(55), Ci => CTMP_55_port, S => 
                           S(55), Co => CTMP_56_port);
   FAI_57 : FA_456 port map( A => A(56), B => B(56), Ci => CTMP_56_port, S => 
                           S(56), Co => CTMP_57_port);
   FAI_58 : FA_455 port map( A => A(57), B => B(57), Ci => CTMP_57_port, S => 
                           S(57), Co => CTMP_58_port);
   FAI_59 : FA_454 port map( A => A(58), B => B(58), Ci => CTMP_58_port, S => 
                           S(58), Co => CTMP_59_port);
   FAI_60 : FA_453 port map( A => A(59), B => B(59), Ci => CTMP_59_port, S => 
                           S(59), Co => CTMP_60_port);
   FAI_61 : FA_452 port map( A => A(60), B => B(60), Ci => CTMP_60_port, S => 
                           S(60), Co => CTMP_61_port);
   FAI_62 : FA_451 port map( A => A(61), B => B(61), Ci => CTMP_61_port, S => 
                           S(61), Co => CTMP_62_port);
   FAI_63 : FA_450 port map( A => A(62), B => B(62), Ci => CTMP_62_port, S => 
                           S(62), Co => CTMP_63_port);
   FAI_64 : FA_449 port map( A => A(63), B => B(63), Ci => CTMP_63_port, S => 
                           S(63), Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity RCA_NbitRca64_7 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_NbitRca64_7;

architecture SYN_STRUCTURAL of RCA_NbitRca64_7 is

   component FA_385
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_386
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_387
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_388
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_389
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_390
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_391
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_392
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_393
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_394
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_395
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_396
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_397
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_398
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_399
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_400
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_401
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_402
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_403
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_404
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_405
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_406
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_407
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_408
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_409
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_410
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_411
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_412
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_413
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_414
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_415
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_416
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_417
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_418
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_419
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_420
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_421
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_422
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_423
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_424
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_425
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_426
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_427
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_428
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_429
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_430
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_431
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_432
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_433
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_434
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_435
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_436
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_437
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_438
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_439
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_440
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_441
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_442
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_443
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_444
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_445
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_446
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_447
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_448
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_63_port, CTMP_62_port, CTMP_61_port, CTMP_60_port, CTMP_59_port,
      CTMP_58_port, CTMP_57_port, CTMP_56_port, CTMP_55_port, CTMP_54_port, 
      CTMP_53_port, CTMP_52_port, CTMP_51_port, CTMP_50_port, CTMP_49_port, 
      CTMP_48_port, CTMP_47_port, CTMP_46_port, CTMP_45_port, CTMP_44_port, 
      CTMP_43_port, CTMP_42_port, CTMP_41_port, CTMP_40_port, CTMP_39_port, 
      CTMP_38_port, CTMP_37_port, CTMP_36_port, CTMP_35_port, CTMP_34_port, 
      CTMP_33_port, CTMP_32_port, CTMP_31_port, CTMP_30_port, CTMP_29_port, 
      CTMP_28_port, CTMP_27_port, CTMP_26_port, CTMP_25_port, CTMP_24_port, 
      CTMP_23_port, CTMP_22_port, CTMP_21_port, CTMP_20_port, CTMP_19_port, 
      CTMP_18_port, CTMP_17_port, CTMP_16_port, CTMP_15_port, CTMP_14_port, 
      CTMP_13_port, CTMP_12_port, CTMP_11_port, CTMP_10_port, CTMP_9_port, 
      CTMP_8_port, CTMP_7_port, CTMP_6_port, CTMP_5_port, CTMP_4_port, 
      CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_448 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_447 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_446 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_445 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => CTMP_4_port);
   FAI_5 : FA_444 port map( A => A(4), B => B(4), Ci => CTMP_4_port, S => S(4),
                           Co => CTMP_5_port);
   FAI_6 : FA_443 port map( A => A(5), B => B(5), Ci => CTMP_5_port, S => S(5),
                           Co => CTMP_6_port);
   FAI_7 : FA_442 port map( A => A(6), B => B(6), Ci => CTMP_6_port, S => S(6),
                           Co => CTMP_7_port);
   FAI_8 : FA_441 port map( A => A(7), B => B(7), Ci => CTMP_7_port, S => S(7),
                           Co => CTMP_8_port);
   FAI_9 : FA_440 port map( A => A(8), B => B(8), Ci => CTMP_8_port, S => S(8),
                           Co => CTMP_9_port);
   FAI_10 : FA_439 port map( A => A(9), B => B(9), Ci => CTMP_9_port, S => S(9)
                           , Co => CTMP_10_port);
   FAI_11 : FA_438 port map( A => A(10), B => B(10), Ci => CTMP_10_port, S => 
                           S(10), Co => CTMP_11_port);
   FAI_12 : FA_437 port map( A => A(11), B => B(11), Ci => CTMP_11_port, S => 
                           S(11), Co => CTMP_12_port);
   FAI_13 : FA_436 port map( A => A(12), B => B(12), Ci => CTMP_12_port, S => 
                           S(12), Co => CTMP_13_port);
   FAI_14 : FA_435 port map( A => A(13), B => B(13), Ci => CTMP_13_port, S => 
                           S(13), Co => CTMP_14_port);
   FAI_15 : FA_434 port map( A => A(14), B => B(14), Ci => CTMP_14_port, S => 
                           S(14), Co => CTMP_15_port);
   FAI_16 : FA_433 port map( A => A(15), B => B(15), Ci => CTMP_15_port, S => 
                           S(15), Co => CTMP_16_port);
   FAI_17 : FA_432 port map( A => A(16), B => B(16), Ci => CTMP_16_port, S => 
                           S(16), Co => CTMP_17_port);
   FAI_18 : FA_431 port map( A => A(17), B => B(17), Ci => CTMP_17_port, S => 
                           S(17), Co => CTMP_18_port);
   FAI_19 : FA_430 port map( A => A(18), B => B(18), Ci => CTMP_18_port, S => 
                           S(18), Co => CTMP_19_port);
   FAI_20 : FA_429 port map( A => A(19), B => B(19), Ci => CTMP_19_port, S => 
                           S(19), Co => CTMP_20_port);
   FAI_21 : FA_428 port map( A => A(20), B => B(20), Ci => CTMP_20_port, S => 
                           S(20), Co => CTMP_21_port);
   FAI_22 : FA_427 port map( A => A(21), B => B(21), Ci => CTMP_21_port, S => 
                           S(21), Co => CTMP_22_port);
   FAI_23 : FA_426 port map( A => A(22), B => B(22), Ci => CTMP_22_port, S => 
                           S(22), Co => CTMP_23_port);
   FAI_24 : FA_425 port map( A => A(23), B => B(23), Ci => CTMP_23_port, S => 
                           S(23), Co => CTMP_24_port);
   FAI_25 : FA_424 port map( A => A(24), B => B(24), Ci => CTMP_24_port, S => 
                           S(24), Co => CTMP_25_port);
   FAI_26 : FA_423 port map( A => A(25), B => B(25), Ci => CTMP_25_port, S => 
                           S(25), Co => CTMP_26_port);
   FAI_27 : FA_422 port map( A => A(26), B => B(26), Ci => CTMP_26_port, S => 
                           S(26), Co => CTMP_27_port);
   FAI_28 : FA_421 port map( A => A(27), B => B(27), Ci => CTMP_27_port, S => 
                           S(27), Co => CTMP_28_port);
   FAI_29 : FA_420 port map( A => A(28), B => B(28), Ci => CTMP_28_port, S => 
                           S(28), Co => CTMP_29_port);
   FAI_30 : FA_419 port map( A => A(29), B => B(29), Ci => CTMP_29_port, S => 
                           S(29), Co => CTMP_30_port);
   FAI_31 : FA_418 port map( A => A(30), B => B(30), Ci => CTMP_30_port, S => 
                           S(30), Co => CTMP_31_port);
   FAI_32 : FA_417 port map( A => A(31), B => B(31), Ci => CTMP_31_port, S => 
                           S(31), Co => CTMP_32_port);
   FAI_33 : FA_416 port map( A => A(32), B => B(32), Ci => CTMP_32_port, S => 
                           S(32), Co => CTMP_33_port);
   FAI_34 : FA_415 port map( A => A(33), B => B(33), Ci => CTMP_33_port, S => 
                           S(33), Co => CTMP_34_port);
   FAI_35 : FA_414 port map( A => A(34), B => B(34), Ci => CTMP_34_port, S => 
                           S(34), Co => CTMP_35_port);
   FAI_36 : FA_413 port map( A => A(35), B => B(35), Ci => CTMP_35_port, S => 
                           S(35), Co => CTMP_36_port);
   FAI_37 : FA_412 port map( A => A(36), B => B(36), Ci => CTMP_36_port, S => 
                           S(36), Co => CTMP_37_port);
   FAI_38 : FA_411 port map( A => A(37), B => B(37), Ci => CTMP_37_port, S => 
                           S(37), Co => CTMP_38_port);
   FAI_39 : FA_410 port map( A => A(38), B => B(38), Ci => CTMP_38_port, S => 
                           S(38), Co => CTMP_39_port);
   FAI_40 : FA_409 port map( A => A(39), B => B(39), Ci => CTMP_39_port, S => 
                           S(39), Co => CTMP_40_port);
   FAI_41 : FA_408 port map( A => A(40), B => B(40), Ci => CTMP_40_port, S => 
                           S(40), Co => CTMP_41_port);
   FAI_42 : FA_407 port map( A => A(41), B => B(41), Ci => CTMP_41_port, S => 
                           S(41), Co => CTMP_42_port);
   FAI_43 : FA_406 port map( A => A(42), B => B(42), Ci => CTMP_42_port, S => 
                           S(42), Co => CTMP_43_port);
   FAI_44 : FA_405 port map( A => A(43), B => B(43), Ci => CTMP_43_port, S => 
                           S(43), Co => CTMP_44_port);
   FAI_45 : FA_404 port map( A => A(44), B => B(44), Ci => CTMP_44_port, S => 
                           S(44), Co => CTMP_45_port);
   FAI_46 : FA_403 port map( A => A(45), B => B(45), Ci => CTMP_45_port, S => 
                           S(45), Co => CTMP_46_port);
   FAI_47 : FA_402 port map( A => A(46), B => B(46), Ci => CTMP_46_port, S => 
                           S(46), Co => CTMP_47_port);
   FAI_48 : FA_401 port map( A => A(47), B => B(47), Ci => CTMP_47_port, S => 
                           S(47), Co => CTMP_48_port);
   FAI_49 : FA_400 port map( A => A(48), B => B(48), Ci => CTMP_48_port, S => 
                           S(48), Co => CTMP_49_port);
   FAI_50 : FA_399 port map( A => A(49), B => B(49), Ci => CTMP_49_port, S => 
                           S(49), Co => CTMP_50_port);
   FAI_51 : FA_398 port map( A => A(50), B => B(50), Ci => CTMP_50_port, S => 
                           S(50), Co => CTMP_51_port);
   FAI_52 : FA_397 port map( A => A(51), B => B(51), Ci => CTMP_51_port, S => 
                           S(51), Co => CTMP_52_port);
   FAI_53 : FA_396 port map( A => A(52), B => B(52), Ci => CTMP_52_port, S => 
                           S(52), Co => CTMP_53_port);
   FAI_54 : FA_395 port map( A => A(53), B => B(53), Ci => CTMP_53_port, S => 
                           S(53), Co => CTMP_54_port);
   FAI_55 : FA_394 port map( A => A(54), B => B(54), Ci => CTMP_54_port, S => 
                           S(54), Co => CTMP_55_port);
   FAI_56 : FA_393 port map( A => A(55), B => B(55), Ci => CTMP_55_port, S => 
                           S(55), Co => CTMP_56_port);
   FAI_57 : FA_392 port map( A => A(56), B => B(56), Ci => CTMP_56_port, S => 
                           S(56), Co => CTMP_57_port);
   FAI_58 : FA_391 port map( A => A(57), B => B(57), Ci => CTMP_57_port, S => 
                           S(57), Co => CTMP_58_port);
   FAI_59 : FA_390 port map( A => A(58), B => B(58), Ci => CTMP_58_port, S => 
                           S(58), Co => CTMP_59_port);
   FAI_60 : FA_389 port map( A => A(59), B => B(59), Ci => CTMP_59_port, S => 
                           S(59), Co => CTMP_60_port);
   FAI_61 : FA_388 port map( A => A(60), B => B(60), Ci => CTMP_60_port, S => 
                           S(60), Co => CTMP_61_port);
   FAI_62 : FA_387 port map( A => A(61), B => B(61), Ci => CTMP_61_port, S => 
                           S(61), Co => CTMP_62_port);
   FAI_63 : FA_386 port map( A => A(62), B => B(62), Ci => CTMP_62_port, S => 
                           S(62), Co => CTMP_63_port);
   FAI_64 : FA_385 port map( A => A(63), B => B(63), Ci => CTMP_63_port, S => 
                           S(63), Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity RCA_NbitRca64_6 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_NbitRca64_6;

architecture SYN_STRUCTURAL of RCA_NbitRca64_6 is

   component FA_321
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_322
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_323
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_324
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_325
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_326
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_327
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_328
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_329
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_330
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_331
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_332
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_333
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_334
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_335
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_336
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_337
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_338
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_339
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_340
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_341
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_342
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_343
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_344
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_345
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_346
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_347
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_348
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_349
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_350
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_351
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_352
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_353
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_354
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_355
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_356
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_357
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_358
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_359
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_360
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_361
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_362
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_363
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_364
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_365
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_366
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_367
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_368
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_369
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_370
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_371
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_372
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_373
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_374
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_375
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_376
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_377
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_378
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_379
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_380
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_381
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_382
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_383
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_384
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_63_port, CTMP_62_port, CTMP_61_port, CTMP_60_port, CTMP_59_port,
      CTMP_58_port, CTMP_57_port, CTMP_56_port, CTMP_55_port, CTMP_54_port, 
      CTMP_53_port, CTMP_52_port, CTMP_51_port, CTMP_50_port, CTMP_49_port, 
      CTMP_48_port, CTMP_47_port, CTMP_46_port, CTMP_45_port, CTMP_44_port, 
      CTMP_43_port, CTMP_42_port, CTMP_41_port, CTMP_40_port, CTMP_39_port, 
      CTMP_38_port, CTMP_37_port, CTMP_36_port, CTMP_35_port, CTMP_34_port, 
      CTMP_33_port, CTMP_32_port, CTMP_31_port, CTMP_30_port, CTMP_29_port, 
      CTMP_28_port, CTMP_27_port, CTMP_26_port, CTMP_25_port, CTMP_24_port, 
      CTMP_23_port, CTMP_22_port, CTMP_21_port, CTMP_20_port, CTMP_19_port, 
      CTMP_18_port, CTMP_17_port, CTMP_16_port, CTMP_15_port, CTMP_14_port, 
      CTMP_13_port, CTMP_12_port, CTMP_11_port, CTMP_10_port, CTMP_9_port, 
      CTMP_8_port, CTMP_7_port, CTMP_6_port, CTMP_5_port, CTMP_4_port, 
      CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_384 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_383 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_382 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_381 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => CTMP_4_port);
   FAI_5 : FA_380 port map( A => A(4), B => B(4), Ci => CTMP_4_port, S => S(4),
                           Co => CTMP_5_port);
   FAI_6 : FA_379 port map( A => A(5), B => B(5), Ci => CTMP_5_port, S => S(5),
                           Co => CTMP_6_port);
   FAI_7 : FA_378 port map( A => A(6), B => B(6), Ci => CTMP_6_port, S => S(6),
                           Co => CTMP_7_port);
   FAI_8 : FA_377 port map( A => A(7), B => B(7), Ci => CTMP_7_port, S => S(7),
                           Co => CTMP_8_port);
   FAI_9 : FA_376 port map( A => A(8), B => B(8), Ci => CTMP_8_port, S => S(8),
                           Co => CTMP_9_port);
   FAI_10 : FA_375 port map( A => A(9), B => B(9), Ci => CTMP_9_port, S => S(9)
                           , Co => CTMP_10_port);
   FAI_11 : FA_374 port map( A => A(10), B => B(10), Ci => CTMP_10_port, S => 
                           S(10), Co => CTMP_11_port);
   FAI_12 : FA_373 port map( A => A(11), B => B(11), Ci => CTMP_11_port, S => 
                           S(11), Co => CTMP_12_port);
   FAI_13 : FA_372 port map( A => A(12), B => B(12), Ci => CTMP_12_port, S => 
                           S(12), Co => CTMP_13_port);
   FAI_14 : FA_371 port map( A => A(13), B => B(13), Ci => CTMP_13_port, S => 
                           S(13), Co => CTMP_14_port);
   FAI_15 : FA_370 port map( A => A(14), B => B(14), Ci => CTMP_14_port, S => 
                           S(14), Co => CTMP_15_port);
   FAI_16 : FA_369 port map( A => A(15), B => B(15), Ci => CTMP_15_port, S => 
                           S(15), Co => CTMP_16_port);
   FAI_17 : FA_368 port map( A => A(16), B => B(16), Ci => CTMP_16_port, S => 
                           S(16), Co => CTMP_17_port);
   FAI_18 : FA_367 port map( A => A(17), B => B(17), Ci => CTMP_17_port, S => 
                           S(17), Co => CTMP_18_port);
   FAI_19 : FA_366 port map( A => A(18), B => B(18), Ci => CTMP_18_port, S => 
                           S(18), Co => CTMP_19_port);
   FAI_20 : FA_365 port map( A => A(19), B => B(19), Ci => CTMP_19_port, S => 
                           S(19), Co => CTMP_20_port);
   FAI_21 : FA_364 port map( A => A(20), B => B(20), Ci => CTMP_20_port, S => 
                           S(20), Co => CTMP_21_port);
   FAI_22 : FA_363 port map( A => A(21), B => B(21), Ci => CTMP_21_port, S => 
                           S(21), Co => CTMP_22_port);
   FAI_23 : FA_362 port map( A => A(22), B => B(22), Ci => CTMP_22_port, S => 
                           S(22), Co => CTMP_23_port);
   FAI_24 : FA_361 port map( A => A(23), B => B(23), Ci => CTMP_23_port, S => 
                           S(23), Co => CTMP_24_port);
   FAI_25 : FA_360 port map( A => A(24), B => B(24), Ci => CTMP_24_port, S => 
                           S(24), Co => CTMP_25_port);
   FAI_26 : FA_359 port map( A => A(25), B => B(25), Ci => CTMP_25_port, S => 
                           S(25), Co => CTMP_26_port);
   FAI_27 : FA_358 port map( A => A(26), B => B(26), Ci => CTMP_26_port, S => 
                           S(26), Co => CTMP_27_port);
   FAI_28 : FA_357 port map( A => A(27), B => B(27), Ci => CTMP_27_port, S => 
                           S(27), Co => CTMP_28_port);
   FAI_29 : FA_356 port map( A => A(28), B => B(28), Ci => CTMP_28_port, S => 
                           S(28), Co => CTMP_29_port);
   FAI_30 : FA_355 port map( A => A(29), B => B(29), Ci => CTMP_29_port, S => 
                           S(29), Co => CTMP_30_port);
   FAI_31 : FA_354 port map( A => A(30), B => B(30), Ci => CTMP_30_port, S => 
                           S(30), Co => CTMP_31_port);
   FAI_32 : FA_353 port map( A => A(31), B => B(31), Ci => CTMP_31_port, S => 
                           S(31), Co => CTMP_32_port);
   FAI_33 : FA_352 port map( A => A(32), B => B(32), Ci => CTMP_32_port, S => 
                           S(32), Co => CTMP_33_port);
   FAI_34 : FA_351 port map( A => A(33), B => B(33), Ci => CTMP_33_port, S => 
                           S(33), Co => CTMP_34_port);
   FAI_35 : FA_350 port map( A => A(34), B => B(34), Ci => CTMP_34_port, S => 
                           S(34), Co => CTMP_35_port);
   FAI_36 : FA_349 port map( A => A(35), B => B(35), Ci => CTMP_35_port, S => 
                           S(35), Co => CTMP_36_port);
   FAI_37 : FA_348 port map( A => A(36), B => B(36), Ci => CTMP_36_port, S => 
                           S(36), Co => CTMP_37_port);
   FAI_38 : FA_347 port map( A => A(37), B => B(37), Ci => CTMP_37_port, S => 
                           S(37), Co => CTMP_38_port);
   FAI_39 : FA_346 port map( A => A(38), B => B(38), Ci => CTMP_38_port, S => 
                           S(38), Co => CTMP_39_port);
   FAI_40 : FA_345 port map( A => A(39), B => B(39), Ci => CTMP_39_port, S => 
                           S(39), Co => CTMP_40_port);
   FAI_41 : FA_344 port map( A => A(40), B => B(40), Ci => CTMP_40_port, S => 
                           S(40), Co => CTMP_41_port);
   FAI_42 : FA_343 port map( A => A(41), B => B(41), Ci => CTMP_41_port, S => 
                           S(41), Co => CTMP_42_port);
   FAI_43 : FA_342 port map( A => A(42), B => B(42), Ci => CTMP_42_port, S => 
                           S(42), Co => CTMP_43_port);
   FAI_44 : FA_341 port map( A => A(43), B => B(43), Ci => CTMP_43_port, S => 
                           S(43), Co => CTMP_44_port);
   FAI_45 : FA_340 port map( A => A(44), B => B(44), Ci => CTMP_44_port, S => 
                           S(44), Co => CTMP_45_port);
   FAI_46 : FA_339 port map( A => A(45), B => B(45), Ci => CTMP_45_port, S => 
                           S(45), Co => CTMP_46_port);
   FAI_47 : FA_338 port map( A => A(46), B => B(46), Ci => CTMP_46_port, S => 
                           S(46), Co => CTMP_47_port);
   FAI_48 : FA_337 port map( A => A(47), B => B(47), Ci => CTMP_47_port, S => 
                           S(47), Co => CTMP_48_port);
   FAI_49 : FA_336 port map( A => A(48), B => B(48), Ci => CTMP_48_port, S => 
                           S(48), Co => CTMP_49_port);
   FAI_50 : FA_335 port map( A => A(49), B => B(49), Ci => CTMP_49_port, S => 
                           S(49), Co => CTMP_50_port);
   FAI_51 : FA_334 port map( A => A(50), B => B(50), Ci => CTMP_50_port, S => 
                           S(50), Co => CTMP_51_port);
   FAI_52 : FA_333 port map( A => A(51), B => B(51), Ci => CTMP_51_port, S => 
                           S(51), Co => CTMP_52_port);
   FAI_53 : FA_332 port map( A => A(52), B => B(52), Ci => CTMP_52_port, S => 
                           S(52), Co => CTMP_53_port);
   FAI_54 : FA_331 port map( A => A(53), B => B(53), Ci => CTMP_53_port, S => 
                           S(53), Co => CTMP_54_port);
   FAI_55 : FA_330 port map( A => A(54), B => B(54), Ci => CTMP_54_port, S => 
                           S(54), Co => CTMP_55_port);
   FAI_56 : FA_329 port map( A => A(55), B => B(55), Ci => CTMP_55_port, S => 
                           S(55), Co => CTMP_56_port);
   FAI_57 : FA_328 port map( A => A(56), B => B(56), Ci => CTMP_56_port, S => 
                           S(56), Co => CTMP_57_port);
   FAI_58 : FA_327 port map( A => A(57), B => B(57), Ci => CTMP_57_port, S => 
                           S(57), Co => CTMP_58_port);
   FAI_59 : FA_326 port map( A => A(58), B => B(58), Ci => CTMP_58_port, S => 
                           S(58), Co => CTMP_59_port);
   FAI_60 : FA_325 port map( A => A(59), B => B(59), Ci => CTMP_59_port, S => 
                           S(59), Co => CTMP_60_port);
   FAI_61 : FA_324 port map( A => A(60), B => B(60), Ci => CTMP_60_port, S => 
                           S(60), Co => CTMP_61_port);
   FAI_62 : FA_323 port map( A => A(61), B => B(61), Ci => CTMP_61_port, S => 
                           S(61), Co => CTMP_62_port);
   FAI_63 : FA_322 port map( A => A(62), B => B(62), Ci => CTMP_62_port, S => 
                           S(62), Co => CTMP_63_port);
   FAI_64 : FA_321 port map( A => A(63), B => B(63), Ci => CTMP_63_port, S => 
                           S(63), Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity RCA_NbitRca64_5 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_NbitRca64_5;

architecture SYN_STRUCTURAL of RCA_NbitRca64_5 is

   component FA_257
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_258
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_259
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_260
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_261
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_262
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_263
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_264
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_265
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_266
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_267
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_268
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_269
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_270
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_271
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_272
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_273
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_274
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_275
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_276
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_277
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_278
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_279
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_280
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_281
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_282
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_283
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_284
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_285
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_286
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_287
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_288
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_289
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_290
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_291
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_292
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_293
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_294
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_295
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_296
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_297
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_298
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_299
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_300
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_301
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_302
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_303
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_304
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_305
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_306
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_307
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_308
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_309
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_310
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_311
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_312
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_313
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_314
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_315
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_316
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_317
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_318
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_319
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_320
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_63_port, CTMP_62_port, CTMP_61_port, CTMP_60_port, CTMP_59_port,
      CTMP_58_port, CTMP_57_port, CTMP_56_port, CTMP_55_port, CTMP_54_port, 
      CTMP_53_port, CTMP_52_port, CTMP_51_port, CTMP_50_port, CTMP_49_port, 
      CTMP_48_port, CTMP_47_port, CTMP_46_port, CTMP_45_port, CTMP_44_port, 
      CTMP_43_port, CTMP_42_port, CTMP_41_port, CTMP_40_port, CTMP_39_port, 
      CTMP_38_port, CTMP_37_port, CTMP_36_port, CTMP_35_port, CTMP_34_port, 
      CTMP_33_port, CTMP_32_port, CTMP_31_port, CTMP_30_port, CTMP_29_port, 
      CTMP_28_port, CTMP_27_port, CTMP_26_port, CTMP_25_port, CTMP_24_port, 
      CTMP_23_port, CTMP_22_port, CTMP_21_port, CTMP_20_port, CTMP_19_port, 
      CTMP_18_port, CTMP_17_port, CTMP_16_port, CTMP_15_port, CTMP_14_port, 
      CTMP_13_port, CTMP_12_port, CTMP_11_port, CTMP_10_port, CTMP_9_port, 
      CTMP_8_port, CTMP_7_port, CTMP_6_port, CTMP_5_port, CTMP_4_port, 
      CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_320 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_319 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_318 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_317 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => CTMP_4_port);
   FAI_5 : FA_316 port map( A => A(4), B => B(4), Ci => CTMP_4_port, S => S(4),
                           Co => CTMP_5_port);
   FAI_6 : FA_315 port map( A => A(5), B => B(5), Ci => CTMP_5_port, S => S(5),
                           Co => CTMP_6_port);
   FAI_7 : FA_314 port map( A => A(6), B => B(6), Ci => CTMP_6_port, S => S(6),
                           Co => CTMP_7_port);
   FAI_8 : FA_313 port map( A => A(7), B => B(7), Ci => CTMP_7_port, S => S(7),
                           Co => CTMP_8_port);
   FAI_9 : FA_312 port map( A => A(8), B => B(8), Ci => CTMP_8_port, S => S(8),
                           Co => CTMP_9_port);
   FAI_10 : FA_311 port map( A => A(9), B => B(9), Ci => CTMP_9_port, S => S(9)
                           , Co => CTMP_10_port);
   FAI_11 : FA_310 port map( A => A(10), B => B(10), Ci => CTMP_10_port, S => 
                           S(10), Co => CTMP_11_port);
   FAI_12 : FA_309 port map( A => A(11), B => B(11), Ci => CTMP_11_port, S => 
                           S(11), Co => CTMP_12_port);
   FAI_13 : FA_308 port map( A => A(12), B => B(12), Ci => CTMP_12_port, S => 
                           S(12), Co => CTMP_13_port);
   FAI_14 : FA_307 port map( A => A(13), B => B(13), Ci => CTMP_13_port, S => 
                           S(13), Co => CTMP_14_port);
   FAI_15 : FA_306 port map( A => A(14), B => B(14), Ci => CTMP_14_port, S => 
                           S(14), Co => CTMP_15_port);
   FAI_16 : FA_305 port map( A => A(15), B => B(15), Ci => CTMP_15_port, S => 
                           S(15), Co => CTMP_16_port);
   FAI_17 : FA_304 port map( A => A(16), B => B(16), Ci => CTMP_16_port, S => 
                           S(16), Co => CTMP_17_port);
   FAI_18 : FA_303 port map( A => A(17), B => B(17), Ci => CTMP_17_port, S => 
                           S(17), Co => CTMP_18_port);
   FAI_19 : FA_302 port map( A => A(18), B => B(18), Ci => CTMP_18_port, S => 
                           S(18), Co => CTMP_19_port);
   FAI_20 : FA_301 port map( A => A(19), B => B(19), Ci => CTMP_19_port, S => 
                           S(19), Co => CTMP_20_port);
   FAI_21 : FA_300 port map( A => A(20), B => B(20), Ci => CTMP_20_port, S => 
                           S(20), Co => CTMP_21_port);
   FAI_22 : FA_299 port map( A => A(21), B => B(21), Ci => CTMP_21_port, S => 
                           S(21), Co => CTMP_22_port);
   FAI_23 : FA_298 port map( A => A(22), B => B(22), Ci => CTMP_22_port, S => 
                           S(22), Co => CTMP_23_port);
   FAI_24 : FA_297 port map( A => A(23), B => B(23), Ci => CTMP_23_port, S => 
                           S(23), Co => CTMP_24_port);
   FAI_25 : FA_296 port map( A => A(24), B => B(24), Ci => CTMP_24_port, S => 
                           S(24), Co => CTMP_25_port);
   FAI_26 : FA_295 port map( A => A(25), B => B(25), Ci => CTMP_25_port, S => 
                           S(25), Co => CTMP_26_port);
   FAI_27 : FA_294 port map( A => A(26), B => B(26), Ci => CTMP_26_port, S => 
                           S(26), Co => CTMP_27_port);
   FAI_28 : FA_293 port map( A => A(27), B => B(27), Ci => CTMP_27_port, S => 
                           S(27), Co => CTMP_28_port);
   FAI_29 : FA_292 port map( A => A(28), B => B(28), Ci => CTMP_28_port, S => 
                           S(28), Co => CTMP_29_port);
   FAI_30 : FA_291 port map( A => A(29), B => B(29), Ci => CTMP_29_port, S => 
                           S(29), Co => CTMP_30_port);
   FAI_31 : FA_290 port map( A => A(30), B => B(30), Ci => CTMP_30_port, S => 
                           S(30), Co => CTMP_31_port);
   FAI_32 : FA_289 port map( A => A(31), B => B(31), Ci => CTMP_31_port, S => 
                           S(31), Co => CTMP_32_port);
   FAI_33 : FA_288 port map( A => A(32), B => B(32), Ci => CTMP_32_port, S => 
                           S(32), Co => CTMP_33_port);
   FAI_34 : FA_287 port map( A => A(33), B => B(33), Ci => CTMP_33_port, S => 
                           S(33), Co => CTMP_34_port);
   FAI_35 : FA_286 port map( A => A(34), B => B(34), Ci => CTMP_34_port, S => 
                           S(34), Co => CTMP_35_port);
   FAI_36 : FA_285 port map( A => A(35), B => B(35), Ci => CTMP_35_port, S => 
                           S(35), Co => CTMP_36_port);
   FAI_37 : FA_284 port map( A => A(36), B => B(36), Ci => CTMP_36_port, S => 
                           S(36), Co => CTMP_37_port);
   FAI_38 : FA_283 port map( A => A(37), B => B(37), Ci => CTMP_37_port, S => 
                           S(37), Co => CTMP_38_port);
   FAI_39 : FA_282 port map( A => A(38), B => B(38), Ci => CTMP_38_port, S => 
                           S(38), Co => CTMP_39_port);
   FAI_40 : FA_281 port map( A => A(39), B => B(39), Ci => CTMP_39_port, S => 
                           S(39), Co => CTMP_40_port);
   FAI_41 : FA_280 port map( A => A(40), B => B(40), Ci => CTMP_40_port, S => 
                           S(40), Co => CTMP_41_port);
   FAI_42 : FA_279 port map( A => A(41), B => B(41), Ci => CTMP_41_port, S => 
                           S(41), Co => CTMP_42_port);
   FAI_43 : FA_278 port map( A => A(42), B => B(42), Ci => CTMP_42_port, S => 
                           S(42), Co => CTMP_43_port);
   FAI_44 : FA_277 port map( A => A(43), B => B(43), Ci => CTMP_43_port, S => 
                           S(43), Co => CTMP_44_port);
   FAI_45 : FA_276 port map( A => A(44), B => B(44), Ci => CTMP_44_port, S => 
                           S(44), Co => CTMP_45_port);
   FAI_46 : FA_275 port map( A => A(45), B => B(45), Ci => CTMP_45_port, S => 
                           S(45), Co => CTMP_46_port);
   FAI_47 : FA_274 port map( A => A(46), B => B(46), Ci => CTMP_46_port, S => 
                           S(46), Co => CTMP_47_port);
   FAI_48 : FA_273 port map( A => A(47), B => B(47), Ci => CTMP_47_port, S => 
                           S(47), Co => CTMP_48_port);
   FAI_49 : FA_272 port map( A => A(48), B => B(48), Ci => CTMP_48_port, S => 
                           S(48), Co => CTMP_49_port);
   FAI_50 : FA_271 port map( A => A(49), B => B(49), Ci => CTMP_49_port, S => 
                           S(49), Co => CTMP_50_port);
   FAI_51 : FA_270 port map( A => A(50), B => B(50), Ci => CTMP_50_port, S => 
                           S(50), Co => CTMP_51_port);
   FAI_52 : FA_269 port map( A => A(51), B => B(51), Ci => CTMP_51_port, S => 
                           S(51), Co => CTMP_52_port);
   FAI_53 : FA_268 port map( A => A(52), B => B(52), Ci => CTMP_52_port, S => 
                           S(52), Co => CTMP_53_port);
   FAI_54 : FA_267 port map( A => A(53), B => B(53), Ci => CTMP_53_port, S => 
                           S(53), Co => CTMP_54_port);
   FAI_55 : FA_266 port map( A => A(54), B => B(54), Ci => CTMP_54_port, S => 
                           S(54), Co => CTMP_55_port);
   FAI_56 : FA_265 port map( A => A(55), B => B(55), Ci => CTMP_55_port, S => 
                           S(55), Co => CTMP_56_port);
   FAI_57 : FA_264 port map( A => A(56), B => B(56), Ci => CTMP_56_port, S => 
                           S(56), Co => CTMP_57_port);
   FAI_58 : FA_263 port map( A => A(57), B => B(57), Ci => CTMP_57_port, S => 
                           S(57), Co => CTMP_58_port);
   FAI_59 : FA_262 port map( A => A(58), B => B(58), Ci => CTMP_58_port, S => 
                           S(58), Co => CTMP_59_port);
   FAI_60 : FA_261 port map( A => A(59), B => B(59), Ci => CTMP_59_port, S => 
                           S(59), Co => CTMP_60_port);
   FAI_61 : FA_260 port map( A => A(60), B => B(60), Ci => CTMP_60_port, S => 
                           S(60), Co => CTMP_61_port);
   FAI_62 : FA_259 port map( A => A(61), B => B(61), Ci => CTMP_61_port, S => 
                           S(61), Co => CTMP_62_port);
   FAI_63 : FA_258 port map( A => A(62), B => B(62), Ci => CTMP_62_port, S => 
                           S(62), Co => CTMP_63_port);
   FAI_64 : FA_257 port map( A => A(63), B => B(63), Ci => CTMP_63_port, S => 
                           S(63), Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity RCA_NbitRca64_4 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_NbitRca64_4;

architecture SYN_STRUCTURAL of RCA_NbitRca64_4 is

   component FA_193
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_194
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_195
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_196
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_197
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_198
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_199
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_200
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_201
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_202
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_203
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_204
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_205
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_206
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_207
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_208
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_209
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_210
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_211
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_212
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_213
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_214
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_215
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_216
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_217
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_218
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_219
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_220
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_221
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_222
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_223
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_224
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_225
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_226
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_227
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_228
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_229
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_230
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_231
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_232
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_233
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_234
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_235
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_236
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_237
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_238
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_239
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_240
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_241
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_242
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_243
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_244
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_245
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_246
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_247
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_248
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_249
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_250
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_251
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_252
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_253
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_254
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_255
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_256
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_63_port, CTMP_62_port, CTMP_61_port, CTMP_60_port, CTMP_59_port,
      CTMP_58_port, CTMP_57_port, CTMP_56_port, CTMP_55_port, CTMP_54_port, 
      CTMP_53_port, CTMP_52_port, CTMP_51_port, CTMP_50_port, CTMP_49_port, 
      CTMP_48_port, CTMP_47_port, CTMP_46_port, CTMP_45_port, CTMP_44_port, 
      CTMP_43_port, CTMP_42_port, CTMP_41_port, CTMP_40_port, CTMP_39_port, 
      CTMP_38_port, CTMP_37_port, CTMP_36_port, CTMP_35_port, CTMP_34_port, 
      CTMP_33_port, CTMP_32_port, CTMP_31_port, CTMP_30_port, CTMP_29_port, 
      CTMP_28_port, CTMP_27_port, CTMP_26_port, CTMP_25_port, CTMP_24_port, 
      CTMP_23_port, CTMP_22_port, CTMP_21_port, CTMP_20_port, CTMP_19_port, 
      CTMP_18_port, CTMP_17_port, CTMP_16_port, CTMP_15_port, CTMP_14_port, 
      CTMP_13_port, CTMP_12_port, CTMP_11_port, CTMP_10_port, CTMP_9_port, 
      CTMP_8_port, CTMP_7_port, CTMP_6_port, CTMP_5_port, CTMP_4_port, 
      CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_256 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_255 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_254 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_253 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => CTMP_4_port);
   FAI_5 : FA_252 port map( A => A(4), B => B(4), Ci => CTMP_4_port, S => S(4),
                           Co => CTMP_5_port);
   FAI_6 : FA_251 port map( A => A(5), B => B(5), Ci => CTMP_5_port, S => S(5),
                           Co => CTMP_6_port);
   FAI_7 : FA_250 port map( A => A(6), B => B(6), Ci => CTMP_6_port, S => S(6),
                           Co => CTMP_7_port);
   FAI_8 : FA_249 port map( A => A(7), B => B(7), Ci => CTMP_7_port, S => S(7),
                           Co => CTMP_8_port);
   FAI_9 : FA_248 port map( A => A(8), B => B(8), Ci => CTMP_8_port, S => S(8),
                           Co => CTMP_9_port);
   FAI_10 : FA_247 port map( A => A(9), B => B(9), Ci => CTMP_9_port, S => S(9)
                           , Co => CTMP_10_port);
   FAI_11 : FA_246 port map( A => A(10), B => B(10), Ci => CTMP_10_port, S => 
                           S(10), Co => CTMP_11_port);
   FAI_12 : FA_245 port map( A => A(11), B => B(11), Ci => CTMP_11_port, S => 
                           S(11), Co => CTMP_12_port);
   FAI_13 : FA_244 port map( A => A(12), B => B(12), Ci => CTMP_12_port, S => 
                           S(12), Co => CTMP_13_port);
   FAI_14 : FA_243 port map( A => A(13), B => B(13), Ci => CTMP_13_port, S => 
                           S(13), Co => CTMP_14_port);
   FAI_15 : FA_242 port map( A => A(14), B => B(14), Ci => CTMP_14_port, S => 
                           S(14), Co => CTMP_15_port);
   FAI_16 : FA_241 port map( A => A(15), B => B(15), Ci => CTMP_15_port, S => 
                           S(15), Co => CTMP_16_port);
   FAI_17 : FA_240 port map( A => A(16), B => B(16), Ci => CTMP_16_port, S => 
                           S(16), Co => CTMP_17_port);
   FAI_18 : FA_239 port map( A => A(17), B => B(17), Ci => CTMP_17_port, S => 
                           S(17), Co => CTMP_18_port);
   FAI_19 : FA_238 port map( A => A(18), B => B(18), Ci => CTMP_18_port, S => 
                           S(18), Co => CTMP_19_port);
   FAI_20 : FA_237 port map( A => A(19), B => B(19), Ci => CTMP_19_port, S => 
                           S(19), Co => CTMP_20_port);
   FAI_21 : FA_236 port map( A => A(20), B => B(20), Ci => CTMP_20_port, S => 
                           S(20), Co => CTMP_21_port);
   FAI_22 : FA_235 port map( A => A(21), B => B(21), Ci => CTMP_21_port, S => 
                           S(21), Co => CTMP_22_port);
   FAI_23 : FA_234 port map( A => A(22), B => B(22), Ci => CTMP_22_port, S => 
                           S(22), Co => CTMP_23_port);
   FAI_24 : FA_233 port map( A => A(23), B => B(23), Ci => CTMP_23_port, S => 
                           S(23), Co => CTMP_24_port);
   FAI_25 : FA_232 port map( A => A(24), B => B(24), Ci => CTMP_24_port, S => 
                           S(24), Co => CTMP_25_port);
   FAI_26 : FA_231 port map( A => A(25), B => B(25), Ci => CTMP_25_port, S => 
                           S(25), Co => CTMP_26_port);
   FAI_27 : FA_230 port map( A => A(26), B => B(26), Ci => CTMP_26_port, S => 
                           S(26), Co => CTMP_27_port);
   FAI_28 : FA_229 port map( A => A(27), B => B(27), Ci => CTMP_27_port, S => 
                           S(27), Co => CTMP_28_port);
   FAI_29 : FA_228 port map( A => A(28), B => B(28), Ci => CTMP_28_port, S => 
                           S(28), Co => CTMP_29_port);
   FAI_30 : FA_227 port map( A => A(29), B => B(29), Ci => CTMP_29_port, S => 
                           S(29), Co => CTMP_30_port);
   FAI_31 : FA_226 port map( A => A(30), B => B(30), Ci => CTMP_30_port, S => 
                           S(30), Co => CTMP_31_port);
   FAI_32 : FA_225 port map( A => A(31), B => B(31), Ci => CTMP_31_port, S => 
                           S(31), Co => CTMP_32_port);
   FAI_33 : FA_224 port map( A => A(32), B => B(32), Ci => CTMP_32_port, S => 
                           S(32), Co => CTMP_33_port);
   FAI_34 : FA_223 port map( A => A(33), B => B(33), Ci => CTMP_33_port, S => 
                           S(33), Co => CTMP_34_port);
   FAI_35 : FA_222 port map( A => A(34), B => B(34), Ci => CTMP_34_port, S => 
                           S(34), Co => CTMP_35_port);
   FAI_36 : FA_221 port map( A => A(35), B => B(35), Ci => CTMP_35_port, S => 
                           S(35), Co => CTMP_36_port);
   FAI_37 : FA_220 port map( A => A(36), B => B(36), Ci => CTMP_36_port, S => 
                           S(36), Co => CTMP_37_port);
   FAI_38 : FA_219 port map( A => A(37), B => B(37), Ci => CTMP_37_port, S => 
                           S(37), Co => CTMP_38_port);
   FAI_39 : FA_218 port map( A => A(38), B => B(38), Ci => CTMP_38_port, S => 
                           S(38), Co => CTMP_39_port);
   FAI_40 : FA_217 port map( A => A(39), B => B(39), Ci => CTMP_39_port, S => 
                           S(39), Co => CTMP_40_port);
   FAI_41 : FA_216 port map( A => A(40), B => B(40), Ci => CTMP_40_port, S => 
                           S(40), Co => CTMP_41_port);
   FAI_42 : FA_215 port map( A => A(41), B => B(41), Ci => CTMP_41_port, S => 
                           S(41), Co => CTMP_42_port);
   FAI_43 : FA_214 port map( A => A(42), B => B(42), Ci => CTMP_42_port, S => 
                           S(42), Co => CTMP_43_port);
   FAI_44 : FA_213 port map( A => A(43), B => B(43), Ci => CTMP_43_port, S => 
                           S(43), Co => CTMP_44_port);
   FAI_45 : FA_212 port map( A => A(44), B => B(44), Ci => CTMP_44_port, S => 
                           S(44), Co => CTMP_45_port);
   FAI_46 : FA_211 port map( A => A(45), B => B(45), Ci => CTMP_45_port, S => 
                           S(45), Co => CTMP_46_port);
   FAI_47 : FA_210 port map( A => A(46), B => B(46), Ci => CTMP_46_port, S => 
                           S(46), Co => CTMP_47_port);
   FAI_48 : FA_209 port map( A => A(47), B => B(47), Ci => CTMP_47_port, S => 
                           S(47), Co => CTMP_48_port);
   FAI_49 : FA_208 port map( A => A(48), B => B(48), Ci => CTMP_48_port, S => 
                           S(48), Co => CTMP_49_port);
   FAI_50 : FA_207 port map( A => A(49), B => B(49), Ci => CTMP_49_port, S => 
                           S(49), Co => CTMP_50_port);
   FAI_51 : FA_206 port map( A => A(50), B => B(50), Ci => CTMP_50_port, S => 
                           S(50), Co => CTMP_51_port);
   FAI_52 : FA_205 port map( A => A(51), B => B(51), Ci => CTMP_51_port, S => 
                           S(51), Co => CTMP_52_port);
   FAI_53 : FA_204 port map( A => A(52), B => B(52), Ci => CTMP_52_port, S => 
                           S(52), Co => CTMP_53_port);
   FAI_54 : FA_203 port map( A => A(53), B => B(53), Ci => CTMP_53_port, S => 
                           S(53), Co => CTMP_54_port);
   FAI_55 : FA_202 port map( A => A(54), B => B(54), Ci => CTMP_54_port, S => 
                           S(54), Co => CTMP_55_port);
   FAI_56 : FA_201 port map( A => A(55), B => B(55), Ci => CTMP_55_port, S => 
                           S(55), Co => CTMP_56_port);
   FAI_57 : FA_200 port map( A => A(56), B => B(56), Ci => CTMP_56_port, S => 
                           S(56), Co => CTMP_57_port);
   FAI_58 : FA_199 port map( A => A(57), B => B(57), Ci => CTMP_57_port, S => 
                           S(57), Co => CTMP_58_port);
   FAI_59 : FA_198 port map( A => A(58), B => B(58), Ci => CTMP_58_port, S => 
                           S(58), Co => CTMP_59_port);
   FAI_60 : FA_197 port map( A => A(59), B => B(59), Ci => CTMP_59_port, S => 
                           S(59), Co => CTMP_60_port);
   FAI_61 : FA_196 port map( A => A(60), B => B(60), Ci => CTMP_60_port, S => 
                           S(60), Co => CTMP_61_port);
   FAI_62 : FA_195 port map( A => A(61), B => B(61), Ci => CTMP_61_port, S => 
                           S(61), Co => CTMP_62_port);
   FAI_63 : FA_194 port map( A => A(62), B => B(62), Ci => CTMP_62_port, S => 
                           S(62), Co => CTMP_63_port);
   FAI_64 : FA_193 port map( A => A(63), B => B(63), Ci => CTMP_63_port, S => 
                           S(63), Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity RCA_NbitRca64_3 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_NbitRca64_3;

architecture SYN_STRUCTURAL of RCA_NbitRca64_3 is

   component FA_129
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_130
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_131
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_132
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_133
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_134
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_135
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_136
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_137
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_138
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_139
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_140
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_141
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_142
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_143
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_144
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_145
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_146
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_147
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_148
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_149
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_150
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_151
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_152
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_153
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_154
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_155
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_156
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_157
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_158
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_159
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_160
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_161
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_162
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_163
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_164
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_165
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_166
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_167
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_168
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_169
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_170
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_171
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_172
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_173
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_174
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_175
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_176
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_177
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_178
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_179
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_180
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_181
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_182
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_183
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_184
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_185
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_186
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_187
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_188
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_189
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_190
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_191
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_192
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_63_port, CTMP_62_port, CTMP_61_port, CTMP_60_port, CTMP_59_port,
      CTMP_58_port, CTMP_57_port, CTMP_56_port, CTMP_55_port, CTMP_54_port, 
      CTMP_53_port, CTMP_52_port, CTMP_51_port, CTMP_50_port, CTMP_49_port, 
      CTMP_48_port, CTMP_47_port, CTMP_46_port, CTMP_45_port, CTMP_44_port, 
      CTMP_43_port, CTMP_42_port, CTMP_41_port, CTMP_40_port, CTMP_39_port, 
      CTMP_38_port, CTMP_37_port, CTMP_36_port, CTMP_35_port, CTMP_34_port, 
      CTMP_33_port, CTMP_32_port, CTMP_31_port, CTMP_30_port, CTMP_29_port, 
      CTMP_28_port, CTMP_27_port, CTMP_26_port, CTMP_25_port, CTMP_24_port, 
      CTMP_23_port, CTMP_22_port, CTMP_21_port, CTMP_20_port, CTMP_19_port, 
      CTMP_18_port, CTMP_17_port, CTMP_16_port, CTMP_15_port, CTMP_14_port, 
      CTMP_13_port, CTMP_12_port, CTMP_11_port, CTMP_10_port, CTMP_9_port, 
      CTMP_8_port, CTMP_7_port, CTMP_6_port, CTMP_5_port, CTMP_4_port, 
      CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_192 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_191 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_190 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_189 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => CTMP_4_port);
   FAI_5 : FA_188 port map( A => A(4), B => B(4), Ci => CTMP_4_port, S => S(4),
                           Co => CTMP_5_port);
   FAI_6 : FA_187 port map( A => A(5), B => B(5), Ci => CTMP_5_port, S => S(5),
                           Co => CTMP_6_port);
   FAI_7 : FA_186 port map( A => A(6), B => B(6), Ci => CTMP_6_port, S => S(6),
                           Co => CTMP_7_port);
   FAI_8 : FA_185 port map( A => A(7), B => B(7), Ci => CTMP_7_port, S => S(7),
                           Co => CTMP_8_port);
   FAI_9 : FA_184 port map( A => A(8), B => B(8), Ci => CTMP_8_port, S => S(8),
                           Co => CTMP_9_port);
   FAI_10 : FA_183 port map( A => A(9), B => B(9), Ci => CTMP_9_port, S => S(9)
                           , Co => CTMP_10_port);
   FAI_11 : FA_182 port map( A => A(10), B => B(10), Ci => CTMP_10_port, S => 
                           S(10), Co => CTMP_11_port);
   FAI_12 : FA_181 port map( A => A(11), B => B(11), Ci => CTMP_11_port, S => 
                           S(11), Co => CTMP_12_port);
   FAI_13 : FA_180 port map( A => A(12), B => B(12), Ci => CTMP_12_port, S => 
                           S(12), Co => CTMP_13_port);
   FAI_14 : FA_179 port map( A => A(13), B => B(13), Ci => CTMP_13_port, S => 
                           S(13), Co => CTMP_14_port);
   FAI_15 : FA_178 port map( A => A(14), B => B(14), Ci => CTMP_14_port, S => 
                           S(14), Co => CTMP_15_port);
   FAI_16 : FA_177 port map( A => A(15), B => B(15), Ci => CTMP_15_port, S => 
                           S(15), Co => CTMP_16_port);
   FAI_17 : FA_176 port map( A => A(16), B => B(16), Ci => CTMP_16_port, S => 
                           S(16), Co => CTMP_17_port);
   FAI_18 : FA_175 port map( A => A(17), B => B(17), Ci => CTMP_17_port, S => 
                           S(17), Co => CTMP_18_port);
   FAI_19 : FA_174 port map( A => A(18), B => B(18), Ci => CTMP_18_port, S => 
                           S(18), Co => CTMP_19_port);
   FAI_20 : FA_173 port map( A => A(19), B => B(19), Ci => CTMP_19_port, S => 
                           S(19), Co => CTMP_20_port);
   FAI_21 : FA_172 port map( A => A(20), B => B(20), Ci => CTMP_20_port, S => 
                           S(20), Co => CTMP_21_port);
   FAI_22 : FA_171 port map( A => A(21), B => B(21), Ci => CTMP_21_port, S => 
                           S(21), Co => CTMP_22_port);
   FAI_23 : FA_170 port map( A => A(22), B => B(22), Ci => CTMP_22_port, S => 
                           S(22), Co => CTMP_23_port);
   FAI_24 : FA_169 port map( A => A(23), B => B(23), Ci => CTMP_23_port, S => 
                           S(23), Co => CTMP_24_port);
   FAI_25 : FA_168 port map( A => A(24), B => B(24), Ci => CTMP_24_port, S => 
                           S(24), Co => CTMP_25_port);
   FAI_26 : FA_167 port map( A => A(25), B => B(25), Ci => CTMP_25_port, S => 
                           S(25), Co => CTMP_26_port);
   FAI_27 : FA_166 port map( A => A(26), B => B(26), Ci => CTMP_26_port, S => 
                           S(26), Co => CTMP_27_port);
   FAI_28 : FA_165 port map( A => A(27), B => B(27), Ci => CTMP_27_port, S => 
                           S(27), Co => CTMP_28_port);
   FAI_29 : FA_164 port map( A => A(28), B => B(28), Ci => CTMP_28_port, S => 
                           S(28), Co => CTMP_29_port);
   FAI_30 : FA_163 port map( A => A(29), B => B(29), Ci => CTMP_29_port, S => 
                           S(29), Co => CTMP_30_port);
   FAI_31 : FA_162 port map( A => A(30), B => B(30), Ci => CTMP_30_port, S => 
                           S(30), Co => CTMP_31_port);
   FAI_32 : FA_161 port map( A => A(31), B => B(31), Ci => CTMP_31_port, S => 
                           S(31), Co => CTMP_32_port);
   FAI_33 : FA_160 port map( A => A(32), B => B(32), Ci => CTMP_32_port, S => 
                           S(32), Co => CTMP_33_port);
   FAI_34 : FA_159 port map( A => A(33), B => B(33), Ci => CTMP_33_port, S => 
                           S(33), Co => CTMP_34_port);
   FAI_35 : FA_158 port map( A => A(34), B => B(34), Ci => CTMP_34_port, S => 
                           S(34), Co => CTMP_35_port);
   FAI_36 : FA_157 port map( A => A(35), B => B(35), Ci => CTMP_35_port, S => 
                           S(35), Co => CTMP_36_port);
   FAI_37 : FA_156 port map( A => A(36), B => B(36), Ci => CTMP_36_port, S => 
                           S(36), Co => CTMP_37_port);
   FAI_38 : FA_155 port map( A => A(37), B => B(37), Ci => CTMP_37_port, S => 
                           S(37), Co => CTMP_38_port);
   FAI_39 : FA_154 port map( A => A(38), B => B(38), Ci => CTMP_38_port, S => 
                           S(38), Co => CTMP_39_port);
   FAI_40 : FA_153 port map( A => A(39), B => B(39), Ci => CTMP_39_port, S => 
                           S(39), Co => CTMP_40_port);
   FAI_41 : FA_152 port map( A => A(40), B => B(40), Ci => CTMP_40_port, S => 
                           S(40), Co => CTMP_41_port);
   FAI_42 : FA_151 port map( A => A(41), B => B(41), Ci => CTMP_41_port, S => 
                           S(41), Co => CTMP_42_port);
   FAI_43 : FA_150 port map( A => A(42), B => B(42), Ci => CTMP_42_port, S => 
                           S(42), Co => CTMP_43_port);
   FAI_44 : FA_149 port map( A => A(43), B => B(43), Ci => CTMP_43_port, S => 
                           S(43), Co => CTMP_44_port);
   FAI_45 : FA_148 port map( A => A(44), B => B(44), Ci => CTMP_44_port, S => 
                           S(44), Co => CTMP_45_port);
   FAI_46 : FA_147 port map( A => A(45), B => B(45), Ci => CTMP_45_port, S => 
                           S(45), Co => CTMP_46_port);
   FAI_47 : FA_146 port map( A => A(46), B => B(46), Ci => CTMP_46_port, S => 
                           S(46), Co => CTMP_47_port);
   FAI_48 : FA_145 port map( A => A(47), B => B(47), Ci => CTMP_47_port, S => 
                           S(47), Co => CTMP_48_port);
   FAI_49 : FA_144 port map( A => A(48), B => B(48), Ci => CTMP_48_port, S => 
                           S(48), Co => CTMP_49_port);
   FAI_50 : FA_143 port map( A => A(49), B => B(49), Ci => CTMP_49_port, S => 
                           S(49), Co => CTMP_50_port);
   FAI_51 : FA_142 port map( A => A(50), B => B(50), Ci => CTMP_50_port, S => 
                           S(50), Co => CTMP_51_port);
   FAI_52 : FA_141 port map( A => A(51), B => B(51), Ci => CTMP_51_port, S => 
                           S(51), Co => CTMP_52_port);
   FAI_53 : FA_140 port map( A => A(52), B => B(52), Ci => CTMP_52_port, S => 
                           S(52), Co => CTMP_53_port);
   FAI_54 : FA_139 port map( A => A(53), B => B(53), Ci => CTMP_53_port, S => 
                           S(53), Co => CTMP_54_port);
   FAI_55 : FA_138 port map( A => A(54), B => B(54), Ci => CTMP_54_port, S => 
                           S(54), Co => CTMP_55_port);
   FAI_56 : FA_137 port map( A => A(55), B => B(55), Ci => CTMP_55_port, S => 
                           S(55), Co => CTMP_56_port);
   FAI_57 : FA_136 port map( A => A(56), B => B(56), Ci => CTMP_56_port, S => 
                           S(56), Co => CTMP_57_port);
   FAI_58 : FA_135 port map( A => A(57), B => B(57), Ci => CTMP_57_port, S => 
                           S(57), Co => CTMP_58_port);
   FAI_59 : FA_134 port map( A => A(58), B => B(58), Ci => CTMP_58_port, S => 
                           S(58), Co => CTMP_59_port);
   FAI_60 : FA_133 port map( A => A(59), B => B(59), Ci => CTMP_59_port, S => 
                           S(59), Co => CTMP_60_port);
   FAI_61 : FA_132 port map( A => A(60), B => B(60), Ci => CTMP_60_port, S => 
                           S(60), Co => CTMP_61_port);
   FAI_62 : FA_131 port map( A => A(61), B => B(61), Ci => CTMP_61_port, S => 
                           S(61), Co => CTMP_62_port);
   FAI_63 : FA_130 port map( A => A(62), B => B(62), Ci => CTMP_62_port, S => 
                           S(62), Co => CTMP_63_port);
   FAI_64 : FA_129 port map( A => A(63), B => B(63), Ci => CTMP_63_port, S => 
                           S(63), Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity RCA_NbitRca64_2 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_NbitRca64_2;

architecture SYN_STRUCTURAL of RCA_NbitRca64_2 is

   component FA_65
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_66
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_67
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_68
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_69
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_70
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_71
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_72
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_73
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_74
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_75
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_76
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_77
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_78
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_79
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_80
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_81
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_82
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_83
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_84
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_85
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_86
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_87
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_88
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_89
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_90
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_91
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_92
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_93
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_94
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_95
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_96
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_97
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_98
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_99
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_100
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_101
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_102
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_103
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_104
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_105
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_106
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_107
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_108
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_109
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_110
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_111
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_112
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_113
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_114
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_115
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_116
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_117
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_118
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_119
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_120
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_121
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_122
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_123
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_124
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_125
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_126
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_127
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_128
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_63_port, CTMP_62_port, CTMP_61_port, CTMP_60_port, CTMP_59_port,
      CTMP_58_port, CTMP_57_port, CTMP_56_port, CTMP_55_port, CTMP_54_port, 
      CTMP_53_port, CTMP_52_port, CTMP_51_port, CTMP_50_port, CTMP_49_port, 
      CTMP_48_port, CTMP_47_port, CTMP_46_port, CTMP_45_port, CTMP_44_port, 
      CTMP_43_port, CTMP_42_port, CTMP_41_port, CTMP_40_port, CTMP_39_port, 
      CTMP_38_port, CTMP_37_port, CTMP_36_port, CTMP_35_port, CTMP_34_port, 
      CTMP_33_port, CTMP_32_port, CTMP_31_port, CTMP_30_port, CTMP_29_port, 
      CTMP_28_port, CTMP_27_port, CTMP_26_port, CTMP_25_port, CTMP_24_port, 
      CTMP_23_port, CTMP_22_port, CTMP_21_port, CTMP_20_port, CTMP_19_port, 
      CTMP_18_port, CTMP_17_port, CTMP_16_port, CTMP_15_port, CTMP_14_port, 
      CTMP_13_port, CTMP_12_port, CTMP_11_port, CTMP_10_port, CTMP_9_port, 
      CTMP_8_port, CTMP_7_port, CTMP_6_port, CTMP_5_port, CTMP_4_port, 
      CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_128 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_127 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_126 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_125 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => CTMP_4_port);
   FAI_5 : FA_124 port map( A => A(4), B => B(4), Ci => CTMP_4_port, S => S(4),
                           Co => CTMP_5_port);
   FAI_6 : FA_123 port map( A => A(5), B => B(5), Ci => CTMP_5_port, S => S(5),
                           Co => CTMP_6_port);
   FAI_7 : FA_122 port map( A => A(6), B => B(6), Ci => CTMP_6_port, S => S(6),
                           Co => CTMP_7_port);
   FAI_8 : FA_121 port map( A => A(7), B => B(7), Ci => CTMP_7_port, S => S(7),
                           Co => CTMP_8_port);
   FAI_9 : FA_120 port map( A => A(8), B => B(8), Ci => CTMP_8_port, S => S(8),
                           Co => CTMP_9_port);
   FAI_10 : FA_119 port map( A => A(9), B => B(9), Ci => CTMP_9_port, S => S(9)
                           , Co => CTMP_10_port);
   FAI_11 : FA_118 port map( A => A(10), B => B(10), Ci => CTMP_10_port, S => 
                           S(10), Co => CTMP_11_port);
   FAI_12 : FA_117 port map( A => A(11), B => B(11), Ci => CTMP_11_port, S => 
                           S(11), Co => CTMP_12_port);
   FAI_13 : FA_116 port map( A => A(12), B => B(12), Ci => CTMP_12_port, S => 
                           S(12), Co => CTMP_13_port);
   FAI_14 : FA_115 port map( A => A(13), B => B(13), Ci => CTMP_13_port, S => 
                           S(13), Co => CTMP_14_port);
   FAI_15 : FA_114 port map( A => A(14), B => B(14), Ci => CTMP_14_port, S => 
                           S(14), Co => CTMP_15_port);
   FAI_16 : FA_113 port map( A => A(15), B => B(15), Ci => CTMP_15_port, S => 
                           S(15), Co => CTMP_16_port);
   FAI_17 : FA_112 port map( A => A(16), B => B(16), Ci => CTMP_16_port, S => 
                           S(16), Co => CTMP_17_port);
   FAI_18 : FA_111 port map( A => A(17), B => B(17), Ci => CTMP_17_port, S => 
                           S(17), Co => CTMP_18_port);
   FAI_19 : FA_110 port map( A => A(18), B => B(18), Ci => CTMP_18_port, S => 
                           S(18), Co => CTMP_19_port);
   FAI_20 : FA_109 port map( A => A(19), B => B(19), Ci => CTMP_19_port, S => 
                           S(19), Co => CTMP_20_port);
   FAI_21 : FA_108 port map( A => A(20), B => B(20), Ci => CTMP_20_port, S => 
                           S(20), Co => CTMP_21_port);
   FAI_22 : FA_107 port map( A => A(21), B => B(21), Ci => CTMP_21_port, S => 
                           S(21), Co => CTMP_22_port);
   FAI_23 : FA_106 port map( A => A(22), B => B(22), Ci => CTMP_22_port, S => 
                           S(22), Co => CTMP_23_port);
   FAI_24 : FA_105 port map( A => A(23), B => B(23), Ci => CTMP_23_port, S => 
                           S(23), Co => CTMP_24_port);
   FAI_25 : FA_104 port map( A => A(24), B => B(24), Ci => CTMP_24_port, S => 
                           S(24), Co => CTMP_25_port);
   FAI_26 : FA_103 port map( A => A(25), B => B(25), Ci => CTMP_25_port, S => 
                           S(25), Co => CTMP_26_port);
   FAI_27 : FA_102 port map( A => A(26), B => B(26), Ci => CTMP_26_port, S => 
                           S(26), Co => CTMP_27_port);
   FAI_28 : FA_101 port map( A => A(27), B => B(27), Ci => CTMP_27_port, S => 
                           S(27), Co => CTMP_28_port);
   FAI_29 : FA_100 port map( A => A(28), B => B(28), Ci => CTMP_28_port, S => 
                           S(28), Co => CTMP_29_port);
   FAI_30 : FA_99 port map( A => A(29), B => B(29), Ci => CTMP_29_port, S => 
                           S(29), Co => CTMP_30_port);
   FAI_31 : FA_98 port map( A => A(30), B => B(30), Ci => CTMP_30_port, S => 
                           S(30), Co => CTMP_31_port);
   FAI_32 : FA_97 port map( A => A(31), B => B(31), Ci => CTMP_31_port, S => 
                           S(31), Co => CTMP_32_port);
   FAI_33 : FA_96 port map( A => A(32), B => B(32), Ci => CTMP_32_port, S => 
                           S(32), Co => CTMP_33_port);
   FAI_34 : FA_95 port map( A => A(33), B => B(33), Ci => CTMP_33_port, S => 
                           S(33), Co => CTMP_34_port);
   FAI_35 : FA_94 port map( A => A(34), B => B(34), Ci => CTMP_34_port, S => 
                           S(34), Co => CTMP_35_port);
   FAI_36 : FA_93 port map( A => A(35), B => B(35), Ci => CTMP_35_port, S => 
                           S(35), Co => CTMP_36_port);
   FAI_37 : FA_92 port map( A => A(36), B => B(36), Ci => CTMP_36_port, S => 
                           S(36), Co => CTMP_37_port);
   FAI_38 : FA_91 port map( A => A(37), B => B(37), Ci => CTMP_37_port, S => 
                           S(37), Co => CTMP_38_port);
   FAI_39 : FA_90 port map( A => A(38), B => B(38), Ci => CTMP_38_port, S => 
                           S(38), Co => CTMP_39_port);
   FAI_40 : FA_89 port map( A => A(39), B => B(39), Ci => CTMP_39_port, S => 
                           S(39), Co => CTMP_40_port);
   FAI_41 : FA_88 port map( A => A(40), B => B(40), Ci => CTMP_40_port, S => 
                           S(40), Co => CTMP_41_port);
   FAI_42 : FA_87 port map( A => A(41), B => B(41), Ci => CTMP_41_port, S => 
                           S(41), Co => CTMP_42_port);
   FAI_43 : FA_86 port map( A => A(42), B => B(42), Ci => CTMP_42_port, S => 
                           S(42), Co => CTMP_43_port);
   FAI_44 : FA_85 port map( A => A(43), B => B(43), Ci => CTMP_43_port, S => 
                           S(43), Co => CTMP_44_port);
   FAI_45 : FA_84 port map( A => A(44), B => B(44), Ci => CTMP_44_port, S => 
                           S(44), Co => CTMP_45_port);
   FAI_46 : FA_83 port map( A => A(45), B => B(45), Ci => CTMP_45_port, S => 
                           S(45), Co => CTMP_46_port);
   FAI_47 : FA_82 port map( A => A(46), B => B(46), Ci => CTMP_46_port, S => 
                           S(46), Co => CTMP_47_port);
   FAI_48 : FA_81 port map( A => A(47), B => B(47), Ci => CTMP_47_port, S => 
                           S(47), Co => CTMP_48_port);
   FAI_49 : FA_80 port map( A => A(48), B => B(48), Ci => CTMP_48_port, S => 
                           S(48), Co => CTMP_49_port);
   FAI_50 : FA_79 port map( A => A(49), B => B(49), Ci => CTMP_49_port, S => 
                           S(49), Co => CTMP_50_port);
   FAI_51 : FA_78 port map( A => A(50), B => B(50), Ci => CTMP_50_port, S => 
                           S(50), Co => CTMP_51_port);
   FAI_52 : FA_77 port map( A => A(51), B => B(51), Ci => CTMP_51_port, S => 
                           S(51), Co => CTMP_52_port);
   FAI_53 : FA_76 port map( A => A(52), B => B(52), Ci => CTMP_52_port, S => 
                           S(52), Co => CTMP_53_port);
   FAI_54 : FA_75 port map( A => A(53), B => B(53), Ci => CTMP_53_port, S => 
                           S(53), Co => CTMP_54_port);
   FAI_55 : FA_74 port map( A => A(54), B => B(54), Ci => CTMP_54_port, S => 
                           S(54), Co => CTMP_55_port);
   FAI_56 : FA_73 port map( A => A(55), B => B(55), Ci => CTMP_55_port, S => 
                           S(55), Co => CTMP_56_port);
   FAI_57 : FA_72 port map( A => A(56), B => B(56), Ci => CTMP_56_port, S => 
                           S(56), Co => CTMP_57_port);
   FAI_58 : FA_71 port map( A => A(57), B => B(57), Ci => CTMP_57_port, S => 
                           S(57), Co => CTMP_58_port);
   FAI_59 : FA_70 port map( A => A(58), B => B(58), Ci => CTMP_58_port, S => 
                           S(58), Co => CTMP_59_port);
   FAI_60 : FA_69 port map( A => A(59), B => B(59), Ci => CTMP_59_port, S => 
                           S(59), Co => CTMP_60_port);
   FAI_61 : FA_68 port map( A => A(60), B => B(60), Ci => CTMP_60_port, S => 
                           S(60), Co => CTMP_61_port);
   FAI_62 : FA_67 port map( A => A(61), B => B(61), Ci => CTMP_61_port, S => 
                           S(61), Co => CTMP_62_port);
   FAI_63 : FA_66 port map( A => A(62), B => B(62), Ci => CTMP_62_port, S => 
                           S(62), Co => CTMP_63_port);
   FAI_64 : FA_65 port map( A => A(63), B => B(63), Ci => CTMP_63_port, S => 
                           S(63), Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity RCA_NbitRca64_1 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_NbitRca64_1;

architecture SYN_STRUCTURAL of RCA_NbitRca64_1 is

   component FA_1
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_2
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_3
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_4
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_5
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_6
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_7
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_8
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_9
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_10
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_11
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_12
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_13
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_14
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_15
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_16
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_17
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_18
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_19
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_20
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_21
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_22
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_23
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_24
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_25
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_26
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_27
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_28
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_29
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_30
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_31
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_32
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_33
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_34
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_35
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_36
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_37
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_38
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_39
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_40
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_41
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_42
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_43
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_44
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_45
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_46
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_47
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_48
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_49
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_50
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_51
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_52
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_53
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_54
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_55
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_56
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_57
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_58
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_59
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_60
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_61
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_62
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_63
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_64
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_63_port, CTMP_62_port, CTMP_61_port, CTMP_60_port, CTMP_59_port,
      CTMP_58_port, CTMP_57_port, CTMP_56_port, CTMP_55_port, CTMP_54_port, 
      CTMP_53_port, CTMP_52_port, CTMP_51_port, CTMP_50_port, CTMP_49_port, 
      CTMP_48_port, CTMP_47_port, CTMP_46_port, CTMP_45_port, CTMP_44_port, 
      CTMP_43_port, CTMP_42_port, CTMP_41_port, CTMP_40_port, CTMP_39_port, 
      CTMP_38_port, CTMP_37_port, CTMP_36_port, CTMP_35_port, CTMP_34_port, 
      CTMP_33_port, CTMP_32_port, CTMP_31_port, CTMP_30_port, CTMP_29_port, 
      CTMP_28_port, CTMP_27_port, CTMP_26_port, CTMP_25_port, CTMP_24_port, 
      CTMP_23_port, CTMP_22_port, CTMP_21_port, CTMP_20_port, CTMP_19_port, 
      CTMP_18_port, CTMP_17_port, CTMP_16_port, CTMP_15_port, CTMP_14_port, 
      CTMP_13_port, CTMP_12_port, CTMP_11_port, CTMP_10_port, CTMP_9_port, 
      CTMP_8_port, CTMP_7_port, CTMP_6_port, CTMP_5_port, CTMP_4_port, 
      CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_64 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_63 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_62 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_61 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => CTMP_4_port);
   FAI_5 : FA_60 port map( A => A(4), B => B(4), Ci => CTMP_4_port, S => S(4), 
                           Co => CTMP_5_port);
   FAI_6 : FA_59 port map( A => A(5), B => B(5), Ci => CTMP_5_port, S => S(5), 
                           Co => CTMP_6_port);
   FAI_7 : FA_58 port map( A => A(6), B => B(6), Ci => CTMP_6_port, S => S(6), 
                           Co => CTMP_7_port);
   FAI_8 : FA_57 port map( A => A(7), B => B(7), Ci => CTMP_7_port, S => S(7), 
                           Co => CTMP_8_port);
   FAI_9 : FA_56 port map( A => A(8), B => B(8), Ci => CTMP_8_port, S => S(8), 
                           Co => CTMP_9_port);
   FAI_10 : FA_55 port map( A => A(9), B => B(9), Ci => CTMP_9_port, S => S(9),
                           Co => CTMP_10_port);
   FAI_11 : FA_54 port map( A => A(10), B => B(10), Ci => CTMP_10_port, S => 
                           S(10), Co => CTMP_11_port);
   FAI_12 : FA_53 port map( A => A(11), B => B(11), Ci => CTMP_11_port, S => 
                           S(11), Co => CTMP_12_port);
   FAI_13 : FA_52 port map( A => A(12), B => B(12), Ci => CTMP_12_port, S => 
                           S(12), Co => CTMP_13_port);
   FAI_14 : FA_51 port map( A => A(13), B => B(13), Ci => CTMP_13_port, S => 
                           S(13), Co => CTMP_14_port);
   FAI_15 : FA_50 port map( A => A(14), B => B(14), Ci => CTMP_14_port, S => 
                           S(14), Co => CTMP_15_port);
   FAI_16 : FA_49 port map( A => A(15), B => B(15), Ci => CTMP_15_port, S => 
                           S(15), Co => CTMP_16_port);
   FAI_17 : FA_48 port map( A => A(16), B => B(16), Ci => CTMP_16_port, S => 
                           S(16), Co => CTMP_17_port);
   FAI_18 : FA_47 port map( A => A(17), B => B(17), Ci => CTMP_17_port, S => 
                           S(17), Co => CTMP_18_port);
   FAI_19 : FA_46 port map( A => A(18), B => B(18), Ci => CTMP_18_port, S => 
                           S(18), Co => CTMP_19_port);
   FAI_20 : FA_45 port map( A => A(19), B => B(19), Ci => CTMP_19_port, S => 
                           S(19), Co => CTMP_20_port);
   FAI_21 : FA_44 port map( A => A(20), B => B(20), Ci => CTMP_20_port, S => 
                           S(20), Co => CTMP_21_port);
   FAI_22 : FA_43 port map( A => A(21), B => B(21), Ci => CTMP_21_port, S => 
                           S(21), Co => CTMP_22_port);
   FAI_23 : FA_42 port map( A => A(22), B => B(22), Ci => CTMP_22_port, S => 
                           S(22), Co => CTMP_23_port);
   FAI_24 : FA_41 port map( A => A(23), B => B(23), Ci => CTMP_23_port, S => 
                           S(23), Co => CTMP_24_port);
   FAI_25 : FA_40 port map( A => A(24), B => B(24), Ci => CTMP_24_port, S => 
                           S(24), Co => CTMP_25_port);
   FAI_26 : FA_39 port map( A => A(25), B => B(25), Ci => CTMP_25_port, S => 
                           S(25), Co => CTMP_26_port);
   FAI_27 : FA_38 port map( A => A(26), B => B(26), Ci => CTMP_26_port, S => 
                           S(26), Co => CTMP_27_port);
   FAI_28 : FA_37 port map( A => A(27), B => B(27), Ci => CTMP_27_port, S => 
                           S(27), Co => CTMP_28_port);
   FAI_29 : FA_36 port map( A => A(28), B => B(28), Ci => CTMP_28_port, S => 
                           S(28), Co => CTMP_29_port);
   FAI_30 : FA_35 port map( A => A(29), B => B(29), Ci => CTMP_29_port, S => 
                           S(29), Co => CTMP_30_port);
   FAI_31 : FA_34 port map( A => A(30), B => B(30), Ci => CTMP_30_port, S => 
                           S(30), Co => CTMP_31_port);
   FAI_32 : FA_33 port map( A => A(31), B => B(31), Ci => CTMP_31_port, S => 
                           S(31), Co => CTMP_32_port);
   FAI_33 : FA_32 port map( A => A(32), B => B(32), Ci => CTMP_32_port, S => 
                           S(32), Co => CTMP_33_port);
   FAI_34 : FA_31 port map( A => A(33), B => B(33), Ci => CTMP_33_port, S => 
                           S(33), Co => CTMP_34_port);
   FAI_35 : FA_30 port map( A => A(34), B => B(34), Ci => CTMP_34_port, S => 
                           S(34), Co => CTMP_35_port);
   FAI_36 : FA_29 port map( A => A(35), B => B(35), Ci => CTMP_35_port, S => 
                           S(35), Co => CTMP_36_port);
   FAI_37 : FA_28 port map( A => A(36), B => B(36), Ci => CTMP_36_port, S => 
                           S(36), Co => CTMP_37_port);
   FAI_38 : FA_27 port map( A => A(37), B => B(37), Ci => CTMP_37_port, S => 
                           S(37), Co => CTMP_38_port);
   FAI_39 : FA_26 port map( A => A(38), B => B(38), Ci => CTMP_38_port, S => 
                           S(38), Co => CTMP_39_port);
   FAI_40 : FA_25 port map( A => A(39), B => B(39), Ci => CTMP_39_port, S => 
                           S(39), Co => CTMP_40_port);
   FAI_41 : FA_24 port map( A => A(40), B => B(40), Ci => CTMP_40_port, S => 
                           S(40), Co => CTMP_41_port);
   FAI_42 : FA_23 port map( A => A(41), B => B(41), Ci => CTMP_41_port, S => 
                           S(41), Co => CTMP_42_port);
   FAI_43 : FA_22 port map( A => A(42), B => B(42), Ci => CTMP_42_port, S => 
                           S(42), Co => CTMP_43_port);
   FAI_44 : FA_21 port map( A => A(43), B => B(43), Ci => CTMP_43_port, S => 
                           S(43), Co => CTMP_44_port);
   FAI_45 : FA_20 port map( A => A(44), B => B(44), Ci => CTMP_44_port, S => 
                           S(44), Co => CTMP_45_port);
   FAI_46 : FA_19 port map( A => A(45), B => B(45), Ci => CTMP_45_port, S => 
                           S(45), Co => CTMP_46_port);
   FAI_47 : FA_18 port map( A => A(46), B => B(46), Ci => CTMP_46_port, S => 
                           S(46), Co => CTMP_47_port);
   FAI_48 : FA_17 port map( A => A(47), B => B(47), Ci => CTMP_47_port, S => 
                           S(47), Co => CTMP_48_port);
   FAI_49 : FA_16 port map( A => A(48), B => B(48), Ci => CTMP_48_port, S => 
                           S(48), Co => CTMP_49_port);
   FAI_50 : FA_15 port map( A => A(49), B => B(49), Ci => CTMP_49_port, S => 
                           S(49), Co => CTMP_50_port);
   FAI_51 : FA_14 port map( A => A(50), B => B(50), Ci => CTMP_50_port, S => 
                           S(50), Co => CTMP_51_port);
   FAI_52 : FA_13 port map( A => A(51), B => B(51), Ci => CTMP_51_port, S => 
                           S(51), Co => CTMP_52_port);
   FAI_53 : FA_12 port map( A => A(52), B => B(52), Ci => CTMP_52_port, S => 
                           S(52), Co => CTMP_53_port);
   FAI_54 : FA_11 port map( A => A(53), B => B(53), Ci => CTMP_53_port, S => 
                           S(53), Co => CTMP_54_port);
   FAI_55 : FA_10 port map( A => A(54), B => B(54), Ci => CTMP_54_port, S => 
                           S(54), Co => CTMP_55_port);
   FAI_56 : FA_9 port map( A => A(55), B => B(55), Ci => CTMP_55_port, S => 
                           S(55), Co => CTMP_56_port);
   FAI_57 : FA_8 port map( A => A(56), B => B(56), Ci => CTMP_56_port, S => 
                           S(56), Co => CTMP_57_port);
   FAI_58 : FA_7 port map( A => A(57), B => B(57), Ci => CTMP_57_port, S => 
                           S(57), Co => CTMP_58_port);
   FAI_59 : FA_6 port map( A => A(58), B => B(58), Ci => CTMP_58_port, S => 
                           S(58), Co => CTMP_59_port);
   FAI_60 : FA_5 port map( A => A(59), B => B(59), Ci => CTMP_59_port, S => 
                           S(59), Co => CTMP_60_port);
   FAI_61 : FA_4 port map( A => A(60), B => B(60), Ci => CTMP_60_port, S => 
                           S(60), Co => CTMP_61_port);
   FAI_62 : FA_3 port map( A => A(61), B => B(61), Ci => CTMP_61_port, S => 
                           S(61), Co => CTMP_62_port);
   FAI_63 : FA_2 port map( A => A(62), B => B(62), Ci => CTMP_62_port, S => 
                           S(62), Co => CTMP_63_port);
   FAI_64 : FA_1 port map( A => A(63), B => B(63), Ci => CTMP_63_port, S => 
                           S(63), Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity IV_63 is

   port( A : in std_logic;  Y : out std_logic);

end IV_63;

architecture SYN_BEHAVIORAL of IV_63 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity IV_62 is

   port( A : in std_logic;  Y : out std_logic);

end IV_62;

architecture SYN_BEHAVIORAL of IV_62 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity IV_61 is

   port( A : in std_logic;  Y : out std_logic);

end IV_61;

architecture SYN_BEHAVIORAL of IV_61 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity IV_60 is

   port( A : in std_logic;  Y : out std_logic);

end IV_60;

architecture SYN_BEHAVIORAL of IV_60 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity IV_59 is

   port( A : in std_logic;  Y : out std_logic);

end IV_59;

architecture SYN_BEHAVIORAL of IV_59 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity IV_58 is

   port( A : in std_logic;  Y : out std_logic);

end IV_58;

architecture SYN_BEHAVIORAL of IV_58 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity IV_57 is

   port( A : in std_logic;  Y : out std_logic);

end IV_57;

architecture SYN_BEHAVIORAL of IV_57 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity IV_56 is

   port( A : in std_logic;  Y : out std_logic);

end IV_56;

architecture SYN_BEHAVIORAL of IV_56 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity IV_55 is

   port( A : in std_logic;  Y : out std_logic);

end IV_55;

architecture SYN_BEHAVIORAL of IV_55 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity IV_54 is

   port( A : in std_logic;  Y : out std_logic);

end IV_54;

architecture SYN_BEHAVIORAL of IV_54 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity IV_53 is

   port( A : in std_logic;  Y : out std_logic);

end IV_53;

architecture SYN_BEHAVIORAL of IV_53 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity IV_52 is

   port( A : in std_logic;  Y : out std_logic);

end IV_52;

architecture SYN_BEHAVIORAL of IV_52 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity IV_51 is

   port( A : in std_logic;  Y : out std_logic);

end IV_51;

architecture SYN_BEHAVIORAL of IV_51 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity IV_50 is

   port( A : in std_logic;  Y : out std_logic);

end IV_50;

architecture SYN_BEHAVIORAL of IV_50 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity IV_49 is

   port( A : in std_logic;  Y : out std_logic);

end IV_49;

architecture SYN_BEHAVIORAL of IV_49 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity IV_48 is

   port( A : in std_logic;  Y : out std_logic);

end IV_48;

architecture SYN_BEHAVIORAL of IV_48 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity IV_47 is

   port( A : in std_logic;  Y : out std_logic);

end IV_47;

architecture SYN_BEHAVIORAL of IV_47 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity IV_46 is

   port( A : in std_logic;  Y : out std_logic);

end IV_46;

architecture SYN_BEHAVIORAL of IV_46 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity IV_45 is

   port( A : in std_logic;  Y : out std_logic);

end IV_45;

architecture SYN_BEHAVIORAL of IV_45 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity IV_44 is

   port( A : in std_logic;  Y : out std_logic);

end IV_44;

architecture SYN_BEHAVIORAL of IV_44 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity IV_43 is

   port( A : in std_logic;  Y : out std_logic);

end IV_43;

architecture SYN_BEHAVIORAL of IV_43 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity IV_42 is

   port( A : in std_logic;  Y : out std_logic);

end IV_42;

architecture SYN_BEHAVIORAL of IV_42 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity IV_41 is

   port( A : in std_logic;  Y : out std_logic);

end IV_41;

architecture SYN_BEHAVIORAL of IV_41 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity IV_40 is

   port( A : in std_logic;  Y : out std_logic);

end IV_40;

architecture SYN_BEHAVIORAL of IV_40 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity IV_39 is

   port( A : in std_logic;  Y : out std_logic);

end IV_39;

architecture SYN_BEHAVIORAL of IV_39 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity IV_38 is

   port( A : in std_logic;  Y : out std_logic);

end IV_38;

architecture SYN_BEHAVIORAL of IV_38 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity IV_37 is

   port( A : in std_logic;  Y : out std_logic);

end IV_37;

architecture SYN_BEHAVIORAL of IV_37 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity IV_36 is

   port( A : in std_logic;  Y : out std_logic);

end IV_36;

architecture SYN_BEHAVIORAL of IV_36 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity IV_35 is

   port( A : in std_logic;  Y : out std_logic);

end IV_35;

architecture SYN_BEHAVIORAL of IV_35 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity IV_34 is

   port( A : in std_logic;  Y : out std_logic);

end IV_34;

architecture SYN_BEHAVIORAL of IV_34 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity IV_33 is

   port( A : in std_logic;  Y : out std_logic);

end IV_33;

architecture SYN_BEHAVIORAL of IV_33 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity IV_32 is

   port( A : in std_logic;  Y : out std_logic);

end IV_32;

architecture SYN_BEHAVIORAL of IV_32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity IV_31 is

   port( A : in std_logic;  Y : out std_logic);

end IV_31;

architecture SYN_BEHAVIORAL of IV_31 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity IV_30 is

   port( A : in std_logic;  Y : out std_logic);

end IV_30;

architecture SYN_BEHAVIORAL of IV_30 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity IV_29 is

   port( A : in std_logic;  Y : out std_logic);

end IV_29;

architecture SYN_BEHAVIORAL of IV_29 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity IV_28 is

   port( A : in std_logic;  Y : out std_logic);

end IV_28;

architecture SYN_BEHAVIORAL of IV_28 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity IV_27 is

   port( A : in std_logic;  Y : out std_logic);

end IV_27;

architecture SYN_BEHAVIORAL of IV_27 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity IV_26 is

   port( A : in std_logic;  Y : out std_logic);

end IV_26;

architecture SYN_BEHAVIORAL of IV_26 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity IV_25 is

   port( A : in std_logic;  Y : out std_logic);

end IV_25;

architecture SYN_BEHAVIORAL of IV_25 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity IV_24 is

   port( A : in std_logic;  Y : out std_logic);

end IV_24;

architecture SYN_BEHAVIORAL of IV_24 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity IV_23 is

   port( A : in std_logic;  Y : out std_logic);

end IV_23;

architecture SYN_BEHAVIORAL of IV_23 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity IV_22 is

   port( A : in std_logic;  Y : out std_logic);

end IV_22;

architecture SYN_BEHAVIORAL of IV_22 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity IV_21 is

   port( A : in std_logic;  Y : out std_logic);

end IV_21;

architecture SYN_BEHAVIORAL of IV_21 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity IV_20 is

   port( A : in std_logic;  Y : out std_logic);

end IV_20;

architecture SYN_BEHAVIORAL of IV_20 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity IV_19 is

   port( A : in std_logic;  Y : out std_logic);

end IV_19;

architecture SYN_BEHAVIORAL of IV_19 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity IV_18 is

   port( A : in std_logic;  Y : out std_logic);

end IV_18;

architecture SYN_BEHAVIORAL of IV_18 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity IV_17 is

   port( A : in std_logic;  Y : out std_logic);

end IV_17;

architecture SYN_BEHAVIORAL of IV_17 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity IV_16 is

   port( A : in std_logic;  Y : out std_logic);

end IV_16;

architecture SYN_BEHAVIORAL of IV_16 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity IV_15 is

   port( A : in std_logic;  Y : out std_logic);

end IV_15;

architecture SYN_BEHAVIORAL of IV_15 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity IV_14 is

   port( A : in std_logic;  Y : out std_logic);

end IV_14;

architecture SYN_BEHAVIORAL of IV_14 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity IV_13 is

   port( A : in std_logic;  Y : out std_logic);

end IV_13;

architecture SYN_BEHAVIORAL of IV_13 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity IV_12 is

   port( A : in std_logic;  Y : out std_logic);

end IV_12;

architecture SYN_BEHAVIORAL of IV_12 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity IV_11 is

   port( A : in std_logic;  Y : out std_logic);

end IV_11;

architecture SYN_BEHAVIORAL of IV_11 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity IV_10 is

   port( A : in std_logic;  Y : out std_logic);

end IV_10;

architecture SYN_BEHAVIORAL of IV_10 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity IV_9 is

   port( A : in std_logic;  Y : out std_logic);

end IV_9;

architecture SYN_BEHAVIORAL of IV_9 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity IV_8 is

   port( A : in std_logic;  Y : out std_logic);

end IV_8;

architecture SYN_BEHAVIORAL of IV_8 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity IV_7 is

   port( A : in std_logic;  Y : out std_logic);

end IV_7;

architecture SYN_BEHAVIORAL of IV_7 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity IV_6 is

   port( A : in std_logic;  Y : out std_logic);

end IV_6;

architecture SYN_BEHAVIORAL of IV_6 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity IV_5 is

   port( A : in std_logic;  Y : out std_logic);

end IV_5;

architecture SYN_BEHAVIORAL of IV_5 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity IV_4 is

   port( A : in std_logic;  Y : out std_logic);

end IV_4;

architecture SYN_BEHAVIORAL of IV_4 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity IV_3 is

   port( A : in std_logic;  Y : out std_logic);

end IV_3;

architecture SYN_BEHAVIORAL of IV_3 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity IV_2 is

   port( A : in std_logic;  Y : out std_logic);

end IV_2;

architecture SYN_BEHAVIORAL of IV_2 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity IV_1 is

   port( A : in std_logic;  Y : out std_logic);

end IV_1;

architecture SYN_BEHAVIORAL of IV_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_971 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_971;

architecture SYN_BEHAVIORAL of FA_971 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X2
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U1 : XOR2_X2 port map( A => Ci, B => n3, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n3, B2 => Ci, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_981 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_981;

architecture SYN_BEHAVIORAL of FA_981 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n2, n3 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U1 : INV_X2 port map( A => n5, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => n3, ZN => n5);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n3, B2 => Ci, ZN => n2);
   U5 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_985 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_985;

architecture SYN_BEHAVIORAL of FA_985 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n3, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U1 : INV_X1 port map( A => n2, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n3, B2 => Ci, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_1023 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1023;

architecture SYN_BEHAVIORAL of FA_1023 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net152921, net180154, n3, n2, n6, n7 : std_logic;

begin
   
   U1 : AOI22_X1 port map( A1 => B, A2 => n7, B1 => Ci, B2 => n3, ZN => n2);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : XNOR2_X1 port map( A => A, B => n6, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n6);
   U5 : XNOR2_X1 port map( A => A, B => n6, ZN => net180154);
   U6 : CLKBUF_X1 port map( A => A, Z => n7);
   U7 : CLKBUF_X1 port map( A => Ci, Z => net152921);
   U8 : XOR2_X1 port map( A => net152921, B => net180154, Z => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity FA_0 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_0;

architecture SYN_BEHAVIORAL of FA_0 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net180091, net179960, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => B, ZN => net179960);
   U2 : AOI21_X1 port map( B1 => A, B2 => Ci, A => B, ZN => n6);
   U3 : NOR2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U4 : CLKBUF_X1 port map( A => A, Z => net180091);
   U5 : NOR2_X1 port map( A1 => net180091, A2 => Ci, ZN => n5);
   U6 : XNOR2_X1 port map( A => net180091, B => net179960, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity RCA_NbitRca64_15 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_NbitRca64_15;

architecture SYN_STRUCTURAL of RCA_NbitRca64_15 is

   component FA_897
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_898
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_899
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_900
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_901
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_902
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_903
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_904
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_905
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_906
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_907
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_908
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_909
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_910
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_911
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_912
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_913
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_914
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_915
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_916
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_917
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_918
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_919
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_920
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_921
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_922
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_923
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_924
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_925
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_926
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_927
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_928
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_929
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_930
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_931
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_932
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_933
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_934
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_935
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_936
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_937
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_938
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_939
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_940
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_941
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_942
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_943
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_944
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_945
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_946
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_947
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_948
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_949
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_950
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_951
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_952
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_953
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_954
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_955
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_956
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_957
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_958
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_959
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_960
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_63_port, CTMP_62_port, CTMP_61_port, CTMP_60_port, CTMP_59_port,
      CTMP_58_port, CTMP_57_port, CTMP_56_port, CTMP_55_port, CTMP_54_port, 
      CTMP_53_port, CTMP_52_port, CTMP_51_port, CTMP_50_port, CTMP_49_port, 
      CTMP_48_port, CTMP_47_port, CTMP_46_port, CTMP_45_port, CTMP_44_port, 
      CTMP_43_port, CTMP_42_port, CTMP_41_port, CTMP_40_port, CTMP_39_port, 
      CTMP_38_port, CTMP_37_port, CTMP_36_port, CTMP_35_port, CTMP_34_port, 
      CTMP_33_port, CTMP_32_port, CTMP_31_port, CTMP_30_port, CTMP_29_port, 
      CTMP_28_port, CTMP_27_port, CTMP_26_port, CTMP_25_port, CTMP_24_port, 
      CTMP_23_port, CTMP_22_port, CTMP_21_port, CTMP_20_port, CTMP_19_port, 
      CTMP_18_port, CTMP_17_port, CTMP_16_port, CTMP_15_port, CTMP_14_port, 
      CTMP_13_port, CTMP_12_port, CTMP_11_port, CTMP_10_port, CTMP_9_port, 
      CTMP_8_port, CTMP_7_port, CTMP_6_port, CTMP_5_port, CTMP_4_port, 
      CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_960 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_959 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_958 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_957 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => CTMP_4_port);
   FAI_5 : FA_956 port map( A => A(4), B => B(4), Ci => CTMP_4_port, S => S(4),
                           Co => CTMP_5_port);
   FAI_6 : FA_955 port map( A => A(5), B => B(5), Ci => CTMP_5_port, S => S(5),
                           Co => CTMP_6_port);
   FAI_7 : FA_954 port map( A => A(6), B => B(6), Ci => CTMP_6_port, S => S(6),
                           Co => CTMP_7_port);
   FAI_8 : FA_953 port map( A => A(7), B => B(7), Ci => CTMP_7_port, S => S(7),
                           Co => CTMP_8_port);
   FAI_9 : FA_952 port map( A => A(8), B => B(8), Ci => CTMP_8_port, S => S(8),
                           Co => CTMP_9_port);
   FAI_10 : FA_951 port map( A => A(9), B => B(9), Ci => CTMP_9_port, S => S(9)
                           , Co => CTMP_10_port);
   FAI_11 : FA_950 port map( A => A(10), B => B(10), Ci => CTMP_10_port, S => 
                           S(10), Co => CTMP_11_port);
   FAI_12 : FA_949 port map( A => A(11), B => B(11), Ci => CTMP_11_port, S => 
                           S(11), Co => CTMP_12_port);
   FAI_13 : FA_948 port map( A => A(12), B => B(12), Ci => CTMP_12_port, S => 
                           S(12), Co => CTMP_13_port);
   FAI_14 : FA_947 port map( A => A(13), B => B(13), Ci => CTMP_13_port, S => 
                           S(13), Co => CTMP_14_port);
   FAI_15 : FA_946 port map( A => A(14), B => B(14), Ci => CTMP_14_port, S => 
                           S(14), Co => CTMP_15_port);
   FAI_16 : FA_945 port map( A => A(15), B => B(15), Ci => CTMP_15_port, S => 
                           S(15), Co => CTMP_16_port);
   FAI_17 : FA_944 port map( A => A(16), B => B(16), Ci => CTMP_16_port, S => 
                           S(16), Co => CTMP_17_port);
   FAI_18 : FA_943 port map( A => A(17), B => B(17), Ci => CTMP_17_port, S => 
                           S(17), Co => CTMP_18_port);
   FAI_19 : FA_942 port map( A => A(18), B => B(18), Ci => CTMP_18_port, S => 
                           S(18), Co => CTMP_19_port);
   FAI_20 : FA_941 port map( A => A(19), B => B(19), Ci => CTMP_19_port, S => 
                           S(19), Co => CTMP_20_port);
   FAI_21 : FA_940 port map( A => A(20), B => B(20), Ci => CTMP_20_port, S => 
                           S(20), Co => CTMP_21_port);
   FAI_22 : FA_939 port map( A => A(21), B => B(21), Ci => CTMP_21_port, S => 
                           S(21), Co => CTMP_22_port);
   FAI_23 : FA_938 port map( A => A(22), B => B(22), Ci => CTMP_22_port, S => 
                           S(22), Co => CTMP_23_port);
   FAI_24 : FA_937 port map( A => A(23), B => B(23), Ci => CTMP_23_port, S => 
                           S(23), Co => CTMP_24_port);
   FAI_25 : FA_936 port map( A => A(24), B => B(24), Ci => CTMP_24_port, S => 
                           S(24), Co => CTMP_25_port);
   FAI_26 : FA_935 port map( A => A(25), B => B(25), Ci => CTMP_25_port, S => 
                           S(25), Co => CTMP_26_port);
   FAI_27 : FA_934 port map( A => A(26), B => B(26), Ci => CTMP_26_port, S => 
                           S(26), Co => CTMP_27_port);
   FAI_28 : FA_933 port map( A => A(27), B => B(27), Ci => CTMP_27_port, S => 
                           S(27), Co => CTMP_28_port);
   FAI_29 : FA_932 port map( A => A(28), B => B(28), Ci => CTMP_28_port, S => 
                           S(28), Co => CTMP_29_port);
   FAI_30 : FA_931 port map( A => A(29), B => B(29), Ci => CTMP_29_port, S => 
                           S(29), Co => CTMP_30_port);
   FAI_31 : FA_930 port map( A => A(30), B => B(30), Ci => CTMP_30_port, S => 
                           S(30), Co => CTMP_31_port);
   FAI_32 : FA_929 port map( A => A(31), B => B(31), Ci => CTMP_31_port, S => 
                           S(31), Co => CTMP_32_port);
   FAI_33 : FA_928 port map( A => A(32), B => B(32), Ci => CTMP_32_port, S => 
                           S(32), Co => CTMP_33_port);
   FAI_34 : FA_927 port map( A => A(33), B => B(33), Ci => CTMP_33_port, S => 
                           S(33), Co => CTMP_34_port);
   FAI_35 : FA_926 port map( A => A(34), B => B(34), Ci => CTMP_34_port, S => 
                           S(34), Co => CTMP_35_port);
   FAI_36 : FA_925 port map( A => A(35), B => B(35), Ci => CTMP_35_port, S => 
                           S(35), Co => CTMP_36_port);
   FAI_37 : FA_924 port map( A => A(36), B => B(36), Ci => CTMP_36_port, S => 
                           S(36), Co => CTMP_37_port);
   FAI_38 : FA_923 port map( A => A(37), B => B(37), Ci => CTMP_37_port, S => 
                           S(37), Co => CTMP_38_port);
   FAI_39 : FA_922 port map( A => A(38), B => B(38), Ci => CTMP_38_port, S => 
                           S(38), Co => CTMP_39_port);
   FAI_40 : FA_921 port map( A => A(39), B => B(39), Ci => CTMP_39_port, S => 
                           S(39), Co => CTMP_40_port);
   FAI_41 : FA_920 port map( A => A(40), B => B(40), Ci => CTMP_40_port, S => 
                           S(40), Co => CTMP_41_port);
   FAI_42 : FA_919 port map( A => A(41), B => B(41), Ci => CTMP_41_port, S => 
                           S(41), Co => CTMP_42_port);
   FAI_43 : FA_918 port map( A => A(42), B => B(42), Ci => CTMP_42_port, S => 
                           S(42), Co => CTMP_43_port);
   FAI_44 : FA_917 port map( A => A(43), B => B(43), Ci => CTMP_43_port, S => 
                           S(43), Co => CTMP_44_port);
   FAI_45 : FA_916 port map( A => A(44), B => B(44), Ci => CTMP_44_port, S => 
                           S(44), Co => CTMP_45_port);
   FAI_46 : FA_915 port map( A => A(45), B => B(45), Ci => CTMP_45_port, S => 
                           S(45), Co => CTMP_46_port);
   FAI_47 : FA_914 port map( A => A(46), B => B(46), Ci => CTMP_46_port, S => 
                           S(46), Co => CTMP_47_port);
   FAI_48 : FA_913 port map( A => A(47), B => B(47), Ci => CTMP_47_port, S => 
                           S(47), Co => CTMP_48_port);
   FAI_49 : FA_912 port map( A => A(48), B => B(48), Ci => CTMP_48_port, S => 
                           S(48), Co => CTMP_49_port);
   FAI_50 : FA_911 port map( A => A(49), B => B(49), Ci => CTMP_49_port, S => 
                           S(49), Co => CTMP_50_port);
   FAI_51 : FA_910 port map( A => A(50), B => B(50), Ci => CTMP_50_port, S => 
                           S(50), Co => CTMP_51_port);
   FAI_52 : FA_909 port map( A => A(51), B => B(51), Ci => CTMP_51_port, S => 
                           S(51), Co => CTMP_52_port);
   FAI_53 : FA_908 port map( A => A(52), B => B(52), Ci => CTMP_52_port, S => 
                           S(52), Co => CTMP_53_port);
   FAI_54 : FA_907 port map( A => A(53), B => B(53), Ci => CTMP_53_port, S => 
                           S(53), Co => CTMP_54_port);
   FAI_55 : FA_906 port map( A => A(54), B => B(54), Ci => CTMP_54_port, S => 
                           S(54), Co => CTMP_55_port);
   FAI_56 : FA_905 port map( A => A(55), B => B(55), Ci => CTMP_55_port, S => 
                           S(55), Co => CTMP_56_port);
   FAI_57 : FA_904 port map( A => A(56), B => B(56), Ci => CTMP_56_port, S => 
                           S(56), Co => CTMP_57_port);
   FAI_58 : FA_903 port map( A => A(57), B => B(57), Ci => CTMP_57_port, S => 
                           S(57), Co => CTMP_58_port);
   FAI_59 : FA_902 port map( A => A(58), B => B(58), Ci => CTMP_58_port, S => 
                           S(58), Co => CTMP_59_port);
   FAI_60 : FA_901 port map( A => A(59), B => B(59), Ci => CTMP_59_port, S => 
                           S(59), Co => CTMP_60_port);
   FAI_61 : FA_900 port map( A => A(60), B => B(60), Ci => CTMP_60_port, S => 
                           S(60), Co => CTMP_61_port);
   FAI_62 : FA_899 port map( A => A(61), B => B(61), Ci => CTMP_61_port, S => 
                           S(61), Co => CTMP_62_port);
   FAI_63 : FA_898 port map( A => A(62), B => B(62), Ci => CTMP_62_port, S => 
                           S(62), Co => CTMP_63_port);
   FAI_64 : FA_897 port map( A => A(63), B => B(63), Ci => CTMP_63_port, S => 
                           S(63), Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity MUX51_MuxNbit64_0 is

   port( zeroSignal, A_signal, A_neg, A_shifted, A_neg_shifted : in 
         std_logic_vector (63 downto 0);  Sel : in std_logic_vector (2 downto 
         0);  Y : out std_logic_vector (63 downto 0));

end MUX51_MuxNbit64_0;

architecture SYN_BEHAVIORAL_2 of MUX51_MuxNbit64_0 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, 
      n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36
      , n37, n38, n39, n40, n41, n42, n43, n44, n45, n48, n49, n50, n51, n52, 
      n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67
      , n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, 
      n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98
      , n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, 
      n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n122, n123, 
      n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, 
      net146356, net146352, net146350, net146348, net146380, net146370, 
      net146368, net146366, net146394, net146412, net146410, net146408, 
      net146406, net146404, net146402, net146430, net146428, net146426, 
      net146424, net146422, net146420, net155681, net155950, net156061, 
      net156060, net156054, net156011, net146414, n46, net166315, net180058, 
      net180057, net156052, net156007, net156006, net146384, net179994, 
      net156057, net156053, net156050, net146416, net146362, n69, n68, n141, 
      n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, 
      n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, 
      n166, n167, n168, n169, n170, n171, n172 : std_logic;

begin
   
   U1 : INV_X1 port map( A => zeroSignal(4), ZN => net156054);
   U2 : NAND2_X1 port map( A1 => net156057, A2 => net156052, ZN => n153);
   U3 : AND2_X1 port map( A1 => n149, A2 => n144, ZN => n141);
   U4 : AND2_X1 port map( A1 => n146, A2 => net156060, ZN => n142);
   U5 : AND2_X1 port map( A1 => A_shifted(9), A2 => net146356, ZN => n143);
   U6 : AND2_X1 port map( A1 => n147, A2 => n148, ZN => n144);
   U7 : INV_X1 port map( A => n155, ZN => net156052);
   U8 : AND2_X1 port map( A1 => zeroSignal(9), A2 => net146380, ZN => n145);
   U9 : OR2_X1 port map( A1 => net156054, A2 => n153, ZN => n146);
   U10 : BUF_X2 port map( A => net146414, Z => net146408);
   U11 : CLKBUF_X1 port map( A => net180057, Z => net146414);
   U12 : INV_X2 port map( A => net156006, ZN => net146356);
   U13 : CLKBUF_X1 port map( A => net146362, Z => net146352);
   U14 : NAND2_X1 port map( A1 => A_shifted(16), A2 => net146348, ZN => n147);
   U15 : NAND2_X1 port map( A1 => zeroSignal(16), A2 => net146366, ZN => n148);
   U16 : NAND2_X1 port map( A1 => A_neg_shifted(16), A2 => net146394, ZN => 
                           n149);
   U17 : AOI211_X1 port map( C1 => A_neg_shifted(9), C2 => n155, A => n145, B 
                           => n143, ZN => n4);
   U18 : AND3_X1 port map( A1 => Sel(0), A2 => n150, A3 => n151, ZN => 
                           net179994);
   U19 : INV_X1 port map( A => Sel(1), ZN => n150);
   U20 : INV_X1 port map( A => Sel(2), ZN => n151);
   U21 : OR2_X1 port map( A1 => net156011, A2 => net180058, ZN => n152);
   U22 : INV_X2 port map( A => n152, ZN => net146406);
   U23 : NAND2_X1 port map( A1 => A_neg_shifted(7), A2 => n155, ZN => n172);
   U24 : NAND2_X1 port map( A1 => n13, A2 => n12, ZN => Y(7));
   U25 : NAND2_X1 port map( A1 => n68, A2 => n69, ZN => Y(3));
   U26 : AOI222_X1 port map( A1 => A_shifted(3), A2 => net146362, B1 => 
                           zeroSignal(3), B2 => net146370, C1 => 
                           A_neg_shifted(3), C2 => n155, ZN => n69);
   U27 : BUF_X1 port map( A => net146380, Z => net146370);
   U28 : INV_X2 port map( A => n153, ZN => net146380);
   U29 : INV_X1 port map( A => net156006, ZN => net146362);
   U30 : NAND2_X1 port map( A1 => A_shifted(4), A2 => net146362, ZN => 
                           net156060);
   U31 : AOI22_X1 port map( A1 => A_neg(3), A2 => net146406, B1 => A_signal(3),
                           B2 => net146424, ZN => n68);
   U32 : BUF_X2 port map( A => net179994, Z => net146424);
   U33 : BUF_X2 port map( A => net179994, Z => net146426);
   U34 : CLKBUF_X1 port map( A => net179994, Z => net146422);
   U35 : INV_X1 port map( A => Sel(0), ZN => net156050);
   U36 : NOR2_X1 port map( A1 => Sel(2), A2 => net156050, ZN => net156007);
   U37 : BUF_X1 port map( A => net180057, Z => net146416);
   U38 : CLKBUF_X1 port map( A => net146416, Z => net146402);
   U39 : AND2_X2 port map( A1 => net156053, A2 => Sel(2), ZN => n155);
   U40 : NAND2_X1 port map( A1 => A_neg_shifted(4), A2 => n155, ZN => net156061
                           );
   U41 : AOI222_X1 port map( A1 => A_shifted(2), A2 => net146352, B1 => 
                           zeroSignal(2), B2 => net146368, C1 => 
                           A_neg_shifted(2), C2 => n155, ZN => n91);
   U42 : NOR2_X1 port map( A1 => Sel(1), A2 => n154, ZN => net156053);
   U43 : BUF_X1 port map( A => Sel(0), Z => n154);
   U44 : OAI21_X1 port map( B1 => Sel(1), B2 => n154, A => n151, ZN => 
                           net156057);
   U45 : INV_X1 port map( A => net156052, ZN => net146384);
   U46 : NAND2_X1 port map( A1 => A_neg_shifted(6), A2 => net146384, ZN => 
                           net166315);
   U47 : AOI222_X1 port map( A1 => A_shifted(5), A2 => net146356, B1 => 
                           zeroSignal(5), B2 => net146380, C1 => 
                           A_neg_shifted(5), C2 => net146384, ZN => n25);
   U48 : INV_X4 port map( A => net156052, ZN => net146394);
   U49 : NAND2_X1 port map( A1 => net156007, A2 => Sel(1), ZN => net156006);
   U50 : OR2_X1 port map( A1 => Sel(2), A2 => Sel(0), ZN => net180058);
   U51 : BUF_X2 port map( A => net146426, Z => net146420);
   U52 : NOR2_X1 port map( A1 => net180058, A2 => net156011, ZN => net180057);
   U53 : BUF_X2 port map( A => net180057, Z => net146404);
   U54 : INV_X1 port map( A => Sel(1), ZN => net156011);
   U55 : NAND2_X1 port map( A1 => A_shifted(14), A2 => net146348, ZN => n156);
   U56 : NAND2_X1 port map( A1 => zeroSignal(14), A2 => net146366, ZN => n157);
   U57 : NAND2_X1 port map( A1 => A_neg_shifted(14), A2 => net146394, ZN => 
                           n158);
   U58 : AND3_X1 port map( A1 => n156, A2 => n157, A3 => n158, ZN => n125);
   U59 : NAND2_X1 port map( A1 => A_shifted(6), A2 => net146356, ZN => n159);
   U60 : NAND2_X1 port map( A1 => zeroSignal(6), A2 => net146380, ZN => n160);
   U61 : AND3_X1 port map( A1 => n159, A2 => n160, A3 => net166315, ZN => n15);
   U62 : NAND3_X1 port map( A1 => n46, A2 => net156061, A3 => n142, ZN => Y(4))
                           ;
   U63 : NAND2_X1 port map( A1 => A_shifted(12), A2 => net146348, ZN => n161);
   U64 : NAND2_X1 port map( A1 => zeroSignal(12), A2 => net146366, ZN => n162);
   U65 : NAND2_X1 port map( A1 => A_neg_shifted(12), A2 => net146394, ZN => 
                           n163);
   U66 : AND3_X1 port map( A1 => n161, A2 => n162, A3 => n163, ZN => n129);
   U67 : NAND2_X1 port map( A1 => A_shifted(10), A2 => net146348, ZN => n164);
   U68 : NAND2_X1 port map( A1 => zeroSignal(10), A2 => net146366, ZN => n165);
   U69 : NAND2_X1 port map( A1 => A_neg_shifted(10), A2 => net146394, ZN => 
                           n166);
   U70 : AND3_X1 port map( A1 => n166, A2 => n165, A3 => n164, ZN => n133);
   U71 : NAND2_X1 port map( A1 => A_shifted(8), A2 => net146356, ZN => n167);
   U72 : NAND2_X1 port map( A1 => zeroSignal(8), A2 => net146380, ZN => n168);
   U73 : NAND2_X1 port map( A1 => A_neg_shifted(8), A2 => net146394, ZN => n169
                           );
   U74 : AND3_X1 port map( A1 => n167, A2 => n168, A3 => n169, ZN => n11);
   U75 : NAND2_X1 port map( A1 => A_shifted(7), A2 => net146356, ZN => n170);
   U76 : NAND2_X1 port map( A1 => zeroSignal(7), A2 => net146380, ZN => n171);
   U77 : AND3_X1 port map( A1 => n170, A2 => n171, A3 => n172, ZN => n13);
   U78 : AOI22_X1 port map( A1 => A_neg(4), A2 => net146408, B1 => A_signal(4),
                           B2 => net146426, ZN => n46);
   U79 : CLKBUF_X1 port map( A => net146420, Z => net146430);
   U80 : BUF_X2 port map( A => net146422, Z => net146428);
   U81 : CLKBUF_X1 port map( A => net146414, Z => net146412);
   U82 : BUF_X2 port map( A => net146414, Z => net146410);
   U83 : CLKBUF_X1 port map( A => net146352, Z => net155681);
   U84 : CLKBUF_X1 port map( A => net146422, Z => net155950);
   U85 : CLKBUF_X1 port map( A => net146356, Z => net146348);
   U86 : CLKBUF_X1 port map( A => net146356, Z => net146350);
   U87 : BUF_X1 port map( A => net146380, Z => net146368);
   U88 : BUF_X1 port map( A => net146380, Z => net146366);
   U89 : NAND2_X1 port map( A1 => n130, A2 => n131, ZN => Y(11));
   U90 : NAND2_X1 port map( A1 => n126, A2 => n127, ZN => Y(13));
   U91 : NAND2_X1 port map( A1 => n42, A2 => n43, ZN => Y(51));
   U92 : AOI222_X1 port map( A1 => A_shifted(51), A2 => net146356, B1 => 
                           zeroSignal(51), B2 => net146380, C1 => 
                           A_neg_shifted(51), C2 => net146394, ZN => n43);
   U93 : AOI22_X1 port map( A1 => A_neg(51), A2 => net146408, B1 => 
                           A_signal(51), B2 => net146426, ZN => n42);
   U94 : NAND2_X1 port map( A1 => n124, A2 => n125, ZN => Y(14));
   U95 : NAND2_X1 port map( A1 => n128, A2 => n129, ZN => Y(12));
   U96 : AOI222_X1 port map( A1 => A_shifted(41), A2 => net146356, B1 => 
                           zeroSignal(41), B2 => net146370, C1 => 
                           A_neg_shifted(41), C2 => net146394, ZN => n65);
   U97 : NAND2_X1 port map( A1 => n40, A2 => n41, ZN => Y(52));
   U98 : AOI222_X1 port map( A1 => A_shifted(52), A2 => net146356, B1 => 
                           zeroSignal(52), B2 => net146380, C1 => 
                           A_neg_shifted(52), C2 => net146394, ZN => n41);
   U99 : AOI22_X1 port map( A1 => A_neg(52), A2 => net146408, B1 => 
                           A_signal(52), B2 => net146426, ZN => n40);
   U100 : AOI222_X1 port map( A1 => A_shifted(15), A2 => net146348, B1 => 
                           zeroSignal(15), B2 => net146366, C1 => 
                           A_neg_shifted(15), C2 => net146394, ZN => n123);
   U101 : NAND2_X1 port map( A1 => n36, A2 => n37, ZN => Y(54));
   U102 : AOI222_X1 port map( A1 => A_shifted(54), A2 => net146356, B1 => 
                           zeroSignal(54), B2 => net146380, C1 => 
                           A_neg_shifted(54), C2 => net146394, ZN => n37);
   U103 : AOI22_X1 port map( A1 => A_neg(54), A2 => net146410, B1 => 
                           A_signal(54), B2 => net146428, ZN => n36);
   U104 : NAND2_X1 port map( A1 => n60, A2 => n61, ZN => Y(43));
   U105 : NAND2_X1 port map( A1 => n118, A2 => n119, ZN => Y(17));
   U106 : AOI222_X1 port map( A1 => A_shifted(17), A2 => net146348, B1 => 
                           zeroSignal(17), B2 => net146366, C1 => 
                           A_neg_shifted(17), C2 => net146394, ZN => n119);
   U107 : NAND2_X1 port map( A1 => n34, A2 => n35, ZN => Y(55));
   U108 : AOI222_X1 port map( A1 => A_shifted(55), A2 => net146356, B1 => 
                           zeroSignal(55), B2 => net146380, C1 => 
                           A_neg_shifted(55), C2 => net146394, ZN => n35);
   U109 : AOI22_X1 port map( A1 => A_neg(55), A2 => net146410, B1 => 
                           A_signal(55), B2 => net146428, ZN => n34);
   U110 : NAND2_X1 port map( A1 => n38, A2 => n39, ZN => Y(53));
   U111 : AOI222_X1 port map( A1 => A_shifted(53), A2 => net146356, B1 => 
                           zeroSignal(53), B2 => net146380, C1 => 
                           A_neg_shifted(53), C2 => net146394, ZN => n39);
   U112 : AOI22_X1 port map( A1 => A_neg(53), A2 => net146410, B1 => 
                           A_signal(53), B2 => net146428, ZN => n38);
   U113 : NAND2_X1 port map( A1 => n32, A2 => n33, ZN => Y(56));
   U114 : AOI222_X1 port map( A1 => A_shifted(56), A2 => net146356, B1 => 
                           zeroSignal(56), B2 => net146380, C1 => 
                           A_neg_shifted(56), C2 => net146394, ZN => n33);
   U115 : AOI22_X1 port map( A1 => A_neg(56), A2 => net146410, B1 => 
                           A_signal(56), B2 => net146428, ZN => n32);
   U116 : AOI222_X1 port map( A1 => A_shifted(45), A2 => net146356, B1 => 
                           zeroSignal(45), B2 => net146380, C1 => 
                           A_neg_shifted(45), C2 => net146394, ZN => n57);
   U117 : NAND2_X1 port map( A1 => n116, A2 => n117, ZN => Y(18));
   U118 : AOI222_X1 port map( A1 => A_shifted(18), A2 => net146348, B1 => 
                           zeroSignal(18), B2 => net146366, C1 => 
                           A_neg_shifted(18), C2 => net146394, ZN => n117);
   U119 : NAND2_X1 port map( A1 => n30, A2 => n31, ZN => Y(57));
   U120 : AOI222_X1 port map( A1 => A_shifted(57), A2 => net146356, B1 => 
                           zeroSignal(57), B2 => net146380, C1 => 
                           A_neg_shifted(57), C2 => net146394, ZN => n31);
   U121 : AOI22_X1 port map( A1 => A_neg(57), A2 => net146410, B1 => 
                           A_signal(57), B2 => net146428, ZN => n30);
   U122 : AOI222_X1 port map( A1 => A_shifted(44), A2 => net146356, B1 => 
                           zeroSignal(44), B2 => net146380, C1 => 
                           A_neg_shifted(44), C2 => net146394, ZN => n59);
   U123 : NAND2_X1 port map( A1 => n106, A2 => n107, ZN => Y(22));
   U124 : AOI222_X1 port map( A1 => A_shifted(22), A2 => net146350, B1 => 
                           zeroSignal(22), B2 => net146368, C1 => 
                           A_neg_shifted(22), C2 => net146394, ZN => n107);
   U125 : AOI222_X1 port map( A1 => A_shifted(20), A2 => net146350, B1 => 
                           zeroSignal(20), B2 => net146368, C1 => 
                           A_neg_shifted(20), C2 => net146394, ZN => n111);
   U126 : NAND2_X1 port map( A1 => n62, A2 => n63, ZN => Y(42));
   U127 : AOI222_X1 port map( A1 => A_shifted(42), A2 => net146356, B1 => 
                           zeroSignal(42), B2 => net146380, C1 => 
                           A_neg_shifted(42), C2 => net146394, ZN => n63);
   U128 : NAND2_X1 port map( A1 => n28, A2 => n29, ZN => Y(58));
   U129 : AOI222_X1 port map( A1 => A_shifted(58), A2 => net146356, B1 => 
                           zeroSignal(58), B2 => net146380, C1 => 
                           A_neg_shifted(58), C2 => net146394, ZN => n29);
   U130 : AOI22_X1 port map( A1 => A_neg(58), A2 => net146410, B1 => 
                           A_signal(58), B2 => net146428, ZN => n28);
   U131 : NAND2_X1 port map( A1 => n102, A2 => n103, ZN => Y(24));
   U132 : AOI222_X1 port map( A1 => A_shifted(24), A2 => net146350, B1 => 
                           zeroSignal(24), B2 => net146368, C1 => 
                           A_neg_shifted(24), C2 => net146394, ZN => n103);
   U133 : AOI22_X1 port map( A1 => A_neg(24), A2 => net146404, B1 => 
                           A_signal(24), B2 => net155950, ZN => n102);
   U134 : NAND2_X1 port map( A1 => n104, A2 => n105, ZN => Y(23));
   U135 : AOI222_X1 port map( A1 => A_shifted(23), A2 => net146350, B1 => 
                           zeroSignal(23), B2 => net146368, C1 => 
                           A_neg_shifted(23), C2 => net146394, ZN => n105);
   U136 : AOI222_X1 port map( A1 => A_shifted(21), A2 => net146350, B1 => 
                           zeroSignal(21), B2 => net146368, C1 => 
                           A_neg_shifted(21), C2 => net146394, ZN => n109);
   U137 : NAND2_X1 port map( A1 => n100, A2 => n101, ZN => Y(25));
   U138 : AOI222_X1 port map( A1 => A_shifted(25), A2 => net146350, B1 => 
                           zeroSignal(25), B2 => net146368, C1 => 
                           A_neg_shifted(25), C2 => net146394, ZN => n101);
   U139 : AOI22_X1 port map( A1 => A_neg(25), A2 => net146404, B1 => 
                           A_signal(25), B2 => net155950, ZN => n100);
   U140 : NAND2_X1 port map( A1 => n26, A2 => n27, ZN => Y(59));
   U141 : AOI222_X1 port map( A1 => A_shifted(59), A2 => net146356, B1 => 
                           zeroSignal(59), B2 => net146380, C1 => 
                           A_neg_shifted(59), C2 => net146394, ZN => n27);
   U142 : AOI22_X1 port map( A1 => A_neg(59), A2 => net146410, B1 => 
                           A_signal(59), B2 => net146428, ZN => n26);
   U143 : NAND2_X1 port map( A1 => n18, A2 => n19, ZN => Y(62));
   U144 : AOI222_X1 port map( A1 => A_shifted(62), A2 => net146356, B1 => 
                           zeroSignal(62), B2 => net146380, C1 => 
                           A_neg_shifted(62), C2 => net146394, ZN => n19);
   U145 : AOI22_X1 port map( A1 => A_neg(62), A2 => net146410, B1 => 
                           A_signal(62), B2 => net146428, ZN => n18);
   U146 : NAND2_X1 port map( A1 => n98, A2 => n99, ZN => Y(26));
   U147 : AOI222_X1 port map( A1 => A_shifted(26), A2 => net146350, B1 => 
                           zeroSignal(26), B2 => net146368, C1 => 
                           A_neg_shifted(26), C2 => net146394, ZN => n99);
   U148 : AOI22_X1 port map( A1 => A_neg(26), A2 => net146404, B1 => 
                           A_signal(26), B2 => net155950, ZN => n98);
   U149 : NAND2_X1 port map( A1 => n16, A2 => n17, ZN => Y(63));
   U150 : AOI222_X1 port map( A1 => A_shifted(63), A2 => net146356, B1 => 
                           zeroSignal(63), B2 => net146380, C1 => 
                           A_neg_shifted(63), C2 => net146394, ZN => n17);
   U151 : AOI22_X1 port map( A1 => A_neg(63), A2 => net146410, B1 => 
                           A_signal(63), B2 => net146428, ZN => n16);
   U152 : NAND2_X1 port map( A1 => n22, A2 => n23, ZN => Y(60));
   U153 : AOI222_X1 port map( A1 => A_shifted(60), A2 => net146356, B1 => 
                           zeroSignal(60), B2 => net146380, C1 => 
                           A_neg_shifted(60), C2 => net146394, ZN => n23);
   U154 : AOI22_X1 port map( A1 => A_neg(60), A2 => net146410, B1 => 
                           A_signal(60), B2 => net146428, ZN => n22);
   U155 : NAND2_X1 port map( A1 => n20, A2 => n21, ZN => Y(61));
   U156 : AOI222_X1 port map( A1 => A_shifted(61), A2 => net146356, B1 => 
                           zeroSignal(61), B2 => net146380, C1 => 
                           A_neg_shifted(61), C2 => net146394, ZN => n21);
   U157 : AOI22_X1 port map( A1 => A_neg(61), A2 => net146410, B1 => 
                           A_signal(61), B2 => net146428, ZN => n20);
   U158 : NAND2_X1 port map( A1 => n88, A2 => n89, ZN => Y(30));
   U159 : AOI22_X1 port map( A1 => A_neg(30), A2 => net146404, B1 => 
                           A_signal(30), B2 => net155950, ZN => n88);
   U160 : AOI222_X1 port map( A1 => A_shifted(28), A2 => net146350, B1 => 
                           zeroSignal(28), B2 => net146368, C1 => 
                           A_neg_shifted(28), C2 => net146394, ZN => n95);
   U161 : AOI22_X1 port map( A1 => A_neg(28), A2 => net146404, B1 => 
                           A_signal(28), B2 => net155950, ZN => n94);
   U162 : AOI222_X1 port map( A1 => A_shifted(31), A2 => net155681, B1 => 
                           zeroSignal(31), B2 => net146370, C1 => 
                           A_neg_shifted(31), C2 => net146394, ZN => n87);
   U163 : AOI22_X1 port map( A1 => A_neg(31), A2 => net146406, B1 => 
                           A_signal(31), B2 => net146424, ZN => n86);
   U164 : AOI222_X1 port map( A1 => A_shifted(27), A2 => net146350, B1 => 
                           zeroSignal(27), B2 => net146368, C1 => 
                           A_neg_shifted(27), C2 => net146394, ZN => n97);
   U165 : AOI222_X1 port map( A1 => A_shifted(32), A2 => net155681, B1 => 
                           zeroSignal(32), B2 => net146370, C1 => 
                           A_neg_shifted(32), C2 => net146394, ZN => n85);
   U166 : AOI22_X1 port map( A1 => A_neg(32), A2 => net146406, B1 => 
                           A_signal(32), B2 => net146424, ZN => n84);
   U167 : NAND2_X1 port map( A1 => n92, A2 => n93, ZN => Y(29));
   U168 : AOI222_X1 port map( A1 => A_shifted(29), A2 => net146350, B1 => 
                           zeroSignal(29), B2 => net146368, C1 => 
                           A_neg_shifted(29), C2 => net146394, ZN => n93);
   U169 : NAND2_X1 port map( A1 => n48, A2 => n49, ZN => Y(49));
   U170 : NAND2_X1 port map( A1 => n82, A2 => n83, ZN => Y(33));
   U171 : AOI222_X1 port map( A1 => A_shifted(33), A2 => net155681, B1 => 
                           zeroSignal(33), B2 => net146370, C1 => 
                           A_neg_shifted(33), C2 => net146394, ZN => n83);
   U172 : AOI22_X1 port map( A1 => A_neg(33), A2 => net146406, B1 => 
                           A_signal(33), B2 => net146424, ZN => n82);
   U173 : AOI222_X1 port map( A1 => A_shifted(34), A2 => net155681, B1 => 
                           zeroSignal(34), B2 => net146370, C1 => 
                           A_neg_shifted(34), C2 => net146394, ZN => n81);
   U174 : AOI22_X1 port map( A1 => A_neg(34), A2 => net146406, B1 => 
                           A_signal(34), B2 => net146424, ZN => n80);
   U175 : AOI222_X1 port map( A1 => A_shifted(48), A2 => net146356, B1 => 
                           zeroSignal(48), B2 => net146380, C1 => 
                           A_neg_shifted(48), C2 => net146394, ZN => n51);
   U176 : NAND2_X1 port map( A1 => n44, A2 => n45, ZN => Y(50));
   U177 : AOI222_X1 port map( A1 => A_shifted(50), A2 => net146356, B1 => 
                           zeroSignal(50), B2 => net146380, C1 => 
                           A_neg_shifted(50), C2 => net146394, ZN => n45);
   U178 : AOI22_X1 port map( A1 => A_neg(40), A2 => net146406, B1 => 
                           A_signal(40), B2 => net146424, ZN => n66);
   U179 : NAND2_X1 port map( A1 => n76, A2 => n77, ZN => Y(36));
   U180 : AOI222_X1 port map( A1 => A_shifted(36), A2 => net155681, B1 => 
                           zeroSignal(36), B2 => net146370, C1 => 
                           A_neg_shifted(36), C2 => net146394, ZN => n77);
   U181 : AOI22_X1 port map( A1 => A_neg(36), A2 => net146406, B1 => 
                           A_signal(36), B2 => net146424, ZN => n76);
   U182 : AOI222_X1 port map( A1 => A_shifted(35), A2 => net155681, B1 => 
                           zeroSignal(35), B2 => net146370, C1 => 
                           A_neg_shifted(35), C2 => net146394, ZN => n79);
   U183 : NAND2_X1 port map( A1 => n74, A2 => n75, ZN => Y(37));
   U184 : AOI222_X1 port map( A1 => A_shifted(37), A2 => net155681, B1 => 
                           zeroSignal(37), B2 => net146370, C1 => 
                           A_neg_shifted(37), C2 => net146394, ZN => n75);
   U185 : AOI22_X1 port map( A1 => A_neg(37), A2 => net146406, B1 => 
                           A_signal(37), B2 => net146424, ZN => n74);
   U186 : NAND2_X1 port map( A1 => n72, A2 => n73, ZN => Y(38));
   U187 : AOI222_X1 port map( A1 => A_shifted(38), A2 => net155681, B1 => 
                           zeroSignal(38), B2 => net146370, C1 => 
                           A_neg_shifted(38), C2 => net146394, ZN => n73);
   U188 : AOI22_X1 port map( A1 => A_neg(38), A2 => net146406, B1 => 
                           A_signal(38), B2 => net146424, ZN => n72);
   U189 : AOI22_X1 port map( A1 => A_neg(1), A2 => net146402, B1 => A_signal(1)
                           , B2 => net146420, ZN => n112);
   U190 : AOI222_X1 port map( A1 => A_shifted(0), A2 => net146348, B1 => 
                           zeroSignal(0), B2 => net146366, C1 => 
                           A_neg_shifted(0), C2 => net146394, ZN => n135);
   U191 : AOI222_X1 port map( A1 => A_shifted(11), A2 => net146348, B1 => 
                           zeroSignal(11), B2 => net146366, C1 => 
                           A_neg_shifted(11), C2 => net146394, ZN => n131);
   U192 : AOI22_X1 port map( A1 => A_neg(2), A2 => net146404, B1 => A_signal(2)
                           , B2 => net146422, ZN => n90);
   U193 : AOI222_X1 port map( A1 => A_shifted(13), A2 => net146348, B1 => 
                           zeroSignal(13), B2 => net146366, C1 => 
                           A_neg_shifted(13), C2 => net146394, ZN => n127);
   U194 : NAND2_X1 port map( A1 => n134, A2 => n135, ZN => Y(0));
   U195 : NAND2_X1 port map( A1 => n112, A2 => n113, ZN => Y(1));
   U196 : AOI222_X1 port map( A1 => A_shifted(49), A2 => net146356, B1 => 
                           zeroSignal(49), B2 => net146380, C1 => 
                           A_neg_shifted(49), C2 => net146394, ZN => n49);
   U197 : NAND2_X1 port map( A1 => n50, A2 => n51, ZN => Y(48));
   U198 : NAND2_X1 port map( A1 => n11, A2 => n10, ZN => Y(8));
   U199 : AOI22_X1 port map( A1 => A_neg(50), A2 => net146408, B1 => 
                           A_signal(50), B2 => net146426, ZN => n44);
   U200 : NAND2_X1 port map( A1 => n3, A2 => n4, ZN => Y(9));
   U201 : NAND2_X1 port map( A1 => n14, A2 => n15, ZN => Y(6));
   U202 : AOI222_X1 port map( A1 => A_shifted(1), A2 => net146350, B1 => 
                           zeroSignal(1), B2 => net146366, C1 => 
                           A_neg_shifted(1), C2 => net146394, ZN => n113);
   U203 : AOI22_X1 port map( A1 => A_neg(0), A2 => net146402, B1 => A_signal(0)
                           , B2 => net146420, ZN => n134);
   U204 : AOI22_X1 port map( A1 => A_neg(49), A2 => net146408, B1 => 
                           A_signal(49), B2 => net146426, ZN => n48);
   U205 : AOI22_X1 port map( A1 => A_neg(48), A2 => net146408, B1 => 
                           A_signal(48), B2 => net146426, ZN => n50);
   U206 : NAND2_X1 port map( A1 => n52, A2 => n53, ZN => Y(47));
   U207 : AOI22_X1 port map( A1 => A_neg(47), A2 => net146408, B1 => 
                           A_signal(47), B2 => net146426, ZN => n52);
   U208 : AOI22_X1 port map( A1 => A_neg(46), A2 => net146408, B1 => 
                           A_signal(46), B2 => net146426, ZN => n54);
   U209 : AOI222_X1 port map( A1 => A_shifted(47), A2 => net146356, B1 => 
                           zeroSignal(47), B2 => net146380, C1 => 
                           A_neg_shifted(47), C2 => net146394, ZN => n53);
   U210 : NAND2_X1 port map( A1 => n54, A2 => n55, ZN => Y(46));
   U211 : NAND2_X1 port map( A1 => n66, A2 => n67, ZN => Y(40));
   U212 : AOI22_X1 port map( A1 => A_neg(35), A2 => net146406, B1 => 
                           A_signal(35), B2 => net146424, ZN => n78);
   U213 : NAND2_X1 port map( A1 => n78, A2 => n79, ZN => Y(35));
   U214 : NAND2_X1 port map( A1 => n90, A2 => n91, ZN => Y(2));
   U215 : NAND2_X1 port map( A1 => n80, A2 => n81, ZN => Y(34));
   U216 : NAND2_X1 port map( A1 => n84, A2 => n85, ZN => Y(32));
   U217 : NAND2_X1 port map( A1 => n56, A2 => n57, ZN => Y(45));
   U218 : AOI222_X1 port map( A1 => A_shifted(46), A2 => net146356, B1 => 
                           zeroSignal(46), B2 => net146380, C1 => 
                           A_neg_shifted(46), C2 => net146394, ZN => n55);
   U219 : AOI22_X1 port map( A1 => A_neg(45), A2 => net146408, B1 => 
                           A_signal(45), B2 => net146426, ZN => n56);
   U220 : AOI222_X1 port map( A1 => A_shifted(43), A2 => net146356, B1 => 
                           zeroSignal(43), B2 => net146380, C1 => 
                           A_neg_shifted(43), C2 => net146394, ZN => n61);
   U221 : AOI22_X1 port map( A1 => A_neg(42), A2 => net146408, B1 => 
                           A_signal(42), B2 => net146426, ZN => n62);
   U222 : NAND2_X1 port map( A1 => n86, A2 => n87, ZN => Y(31));
   U223 : NAND2_X1 port map( A1 => n58, A2 => n59, ZN => Y(44));
   U224 : AOI22_X1 port map( A1 => A_neg(44), A2 => net146408, B1 => 
                           A_signal(44), B2 => net146426, ZN => n58);
   U225 : AOI22_X1 port map( A1 => A_neg(27), A2 => net146404, B1 => 
                           A_signal(27), B2 => net155950, ZN => n96);
   U226 : NAND2_X1 port map( A1 => n96, A2 => n97, ZN => Y(27));
   U227 : AOI222_X1 port map( A1 => A_shifted(30), A2 => net155681, B1 => 
                           zeroSignal(30), B2 => net146368, C1 => 
                           A_neg_shifted(30), C2 => net146394, ZN => n89);
   U228 : AOI22_X1 port map( A1 => A_neg(29), A2 => net146404, B1 => 
                           A_signal(29), B2 => net155950, ZN => n92);
   U229 : AOI22_X1 port map( A1 => A_neg(20), A2 => net146404, B1 => 
                           A_signal(20), B2 => net155950, ZN => n110);
   U230 : NAND2_X1 port map( A1 => n94, A2 => n95, ZN => Y(28));
   U231 : AOI22_X1 port map( A1 => A_neg(23), A2 => net146404, B1 => 
                           A_signal(23), B2 => net155950, ZN => n104);
   U232 : AOI222_X1 port map( A1 => A_shifted(40), A2 => net146356, B1 => 
                           zeroSignal(40), B2 => net146370, C1 => 
                           A_neg_shifted(40), C2 => net146394, ZN => n67);
   U233 : AOI22_X1 port map( A1 => A_neg(43), A2 => net146408, B1 => 
                           A_signal(43), B2 => net146426, ZN => n60);
   U234 : NAND2_X1 port map( A1 => n110, A2 => n111, ZN => Y(20));
   U235 : AOI22_X1 port map( A1 => A_neg(19), A2 => net146402, B1 => 
                           A_signal(19), B2 => net146420, ZN => n114);
   U236 : NAND2_X1 port map( A1 => n114, A2 => n115, ZN => Y(19));
   U237 : AOI22_X1 port map( A1 => A_neg(41), A2 => net146406, B1 => 
                           A_signal(41), B2 => net146424, ZN => n64);
   U238 : AOI222_X1 port map( A1 => A_shifted(19), A2 => net146348, B1 => 
                           zeroSignal(19), B2 => net146366, C1 => 
                           A_neg_shifted(19), C2 => net146394, ZN => n115);
   U239 : AOI22_X1 port map( A1 => A_neg(18), A2 => net146402, B1 => 
                           A_signal(18), B2 => net146420, ZN => n116);
   U240 : AOI22_X1 port map( A1 => A_neg(21), A2 => net146404, B1 => 
                           A_signal(21), B2 => net155950, ZN => n108);
   U241 : NAND2_X1 port map( A1 => n108, A2 => n109, ZN => Y(21));
   U242 : AOI22_X1 port map( A1 => A_neg(16), A2 => net146402, B1 => 
                           A_signal(16), B2 => net146420, ZN => n120);
   U243 : NAND2_X1 port map( A1 => n120, A2 => n141, ZN => Y(16));
   U244 : AOI22_X1 port map( A1 => A_neg(22), A2 => net146404, B1 => 
                           A_signal(22), B2 => net155950, ZN => n106);
   U245 : AOI222_X1 port map( A1 => A_shifted(39), A2 => net155681, B1 => 
                           zeroSignal(39), B2 => net146370, C1 => 
                           A_neg_shifted(39), C2 => net146394, ZN => n71);
   U246 : NAND2_X1 port map( A1 => n64, A2 => n65, ZN => Y(41));
   U247 : AOI22_X1 port map( A1 => A_neg(17), A2 => net146402, B1 => 
                           A_signal(17), B2 => net146420, ZN => n118);
   U248 : NAND2_X1 port map( A1 => n70, A2 => n71, ZN => Y(39));
   U249 : AOI22_X1 port map( A1 => A_neg(14), A2 => net146402, B1 => 
                           A_signal(14), B2 => net146420, ZN => n124);
   U250 : AOI22_X1 port map( A1 => A_neg(12), A2 => net146402, B1 => 
                           A_signal(12), B2 => net146420, ZN => n128);
   U251 : AOI22_X1 port map( A1 => A_neg(10), A2 => net146402, B1 => 
                           A_signal(10), B2 => net146420, ZN => n132);
   U252 : NAND2_X1 port map( A1 => n132, A2 => n133, ZN => Y(10));
   U253 : AOI22_X1 port map( A1 => A_neg(15), A2 => net146402, B1 => 
                           A_signal(15), B2 => net146420, ZN => n122);
   U254 : NAND2_X1 port map( A1 => n122, A2 => n123, ZN => Y(15));
   U255 : AOI22_X1 port map( A1 => A_neg(13), A2 => net146402, B1 => 
                           A_signal(13), B2 => net146420, ZN => n126);
   U256 : AOI22_X1 port map( A1 => A_neg(11), A2 => net146402, B1 => 
                           A_signal(11), B2 => net146420, ZN => n130);
   U257 : AOI22_X1 port map( A1 => A_neg(9), A2 => net146412, B1 => A_signal(9)
                           , B2 => net146430, ZN => n3);
   U258 : AOI22_X1 port map( A1 => A_neg(8), A2 => net146412, B1 => A_signal(8)
                           , B2 => net146430, ZN => n10);
   U259 : AOI22_X1 port map( A1 => A_neg(7), A2 => net146412, B1 => A_signal(7)
                           , B2 => net146430, ZN => n12);
   U260 : AOI22_X1 port map( A1 => A_neg(6), A2 => net146412, B1 => A_signal(6)
                           , B2 => net146430, ZN => n14);
   U261 : AOI22_X1 port map( A1 => A_neg(5), A2 => net146410, B1 => A_signal(5)
                           , B2 => net146428, ZN => n24);
   U262 : NAND2_X1 port map( A1 => n24, A2 => n25, ZN => Y(5));
   U263 : AOI22_X1 port map( A1 => A_neg(39), A2 => net146406, B1 => 
                           A_signal(39), B2 => net146424, ZN => n70);

end SYN_BEHAVIORAL_2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity encoder_0 is

   port( pieceofB : in std_logic_vector (2 downto 0);  sel : out 
         std_logic_vector (2 downto 0));

end encoder_0;

architecture SYN_behavioral of encoder_0 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => pieceofB(1), A2 => pieceofB(0), ZN => n2);
   U4 : AND2_X1 port map( A1 => n2, A2 => pieceofB(2), ZN => n4);
   U5 : AND2_X1 port map( A1 => n3, A2 => n4, ZN => sel(2));
   U6 : INV_X1 port map( A => pieceofB(2), ZN => n1);
   U7 : OAI21_X1 port map( B1 => pieceofB(1), B2 => pieceofB(0), A => n2, ZN =>
                           n3);
   U8 : AOI21_X1 port map( B1 => n3, B2 => n2, A => pieceofB(2), ZN => sel(0));
   U9 : OAI22_X1 port map( A1 => n1, A2 => n3, B1 => pieceofB(2), B2 => n2, ZN 
                           => sel(1));

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity leftshifter_NbitShifter64_0 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_0;

architecture SYN_behavioral of leftshifter_NbitShifter64_0 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity RCA_NbitRca64_0 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_NbitRca64_0;

architecture SYN_STRUCTURAL of RCA_NbitRca64_0 is

   component FA_961
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_962
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_963
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_964
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_965
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_966
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_967
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_968
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_969
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_970
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_971
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_972
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_973
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_974
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_975
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_976
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_977
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_978
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_979
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_980
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_981
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_982
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_983
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_984
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_985
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_986
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_987
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_988
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_989
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_990
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_991
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_992
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_993
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_994
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_995
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_996
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_997
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_998
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_999
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1000
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1001
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1002
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1003
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1004
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1005
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1006
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1007
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1008
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1009
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1010
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1011
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1012
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1013
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1014
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1015
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1016
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1017
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1018
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1019
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1020
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1021
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1022
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1023
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_0
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_63_port, CTMP_62_port, CTMP_61_port, CTMP_60_port, CTMP_59_port,
      CTMP_58_port, CTMP_57_port, CTMP_56_port, CTMP_55_port, CTMP_54_port, 
      CTMP_53_port, CTMP_52_port, CTMP_51_port, CTMP_50_port, CTMP_49_port, 
      CTMP_48_port, CTMP_47_port, CTMP_46_port, CTMP_45_port, CTMP_44_port, 
      CTMP_43_port, CTMP_42_port, CTMP_41_port, CTMP_40_port, CTMP_39_port, 
      CTMP_38_port, CTMP_37_port, CTMP_36_port, CTMP_35_port, CTMP_34_port, 
      CTMP_33_port, CTMP_32_port, CTMP_31_port, CTMP_30_port, CTMP_29_port, 
      CTMP_28_port, CTMP_27_port, CTMP_26_port, CTMP_25_port, CTMP_24_port, 
      CTMP_23_port, CTMP_22_port, CTMP_21_port, CTMP_20_port, CTMP_19_port, 
      CTMP_18_port, CTMP_17_port, CTMP_16_port, CTMP_15_port, CTMP_14_port, 
      CTMP_13_port, CTMP_12_port, CTMP_11_port, CTMP_10_port, CTMP_9_port, 
      CTMP_8_port, CTMP_7_port, CTMP_6_port, CTMP_5_port, CTMP_4_port, 
      CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_0 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_1023 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1)
                           , Co => CTMP_2_port);
   FAI_3 : FA_1022 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2)
                           , Co => CTMP_3_port);
   FAI_4 : FA_1021 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3)
                           , Co => CTMP_4_port);
   FAI_5 : FA_1020 port map( A => A(4), B => B(4), Ci => CTMP_4_port, S => S(4)
                           , Co => CTMP_5_port);
   FAI_6 : FA_1019 port map( A => A(5), B => B(5), Ci => CTMP_5_port, S => S(5)
                           , Co => CTMP_6_port);
   FAI_7 : FA_1018 port map( A => A(6), B => B(6), Ci => CTMP_6_port, S => S(6)
                           , Co => CTMP_7_port);
   FAI_8 : FA_1017 port map( A => A(7), B => B(7), Ci => CTMP_7_port, S => S(7)
                           , Co => CTMP_8_port);
   FAI_9 : FA_1016 port map( A => A(8), B => B(8), Ci => CTMP_8_port, S => S(8)
                           , Co => CTMP_9_port);
   FAI_10 : FA_1015 port map( A => A(9), B => B(9), Ci => CTMP_9_port, S => 
                           S(9), Co => CTMP_10_port);
   FAI_11 : FA_1014 port map( A => A(10), B => B(10), Ci => CTMP_10_port, S => 
                           S(10), Co => CTMP_11_port);
   FAI_12 : FA_1013 port map( A => A(11), B => B(11), Ci => CTMP_11_port, S => 
                           S(11), Co => CTMP_12_port);
   FAI_13 : FA_1012 port map( A => A(12), B => B(12), Ci => CTMP_12_port, S => 
                           S(12), Co => CTMP_13_port);
   FAI_14 : FA_1011 port map( A => A(13), B => B(13), Ci => CTMP_13_port, S => 
                           S(13), Co => CTMP_14_port);
   FAI_15 : FA_1010 port map( A => A(14), B => B(14), Ci => CTMP_14_port, S => 
                           S(14), Co => CTMP_15_port);
   FAI_16 : FA_1009 port map( A => A(15), B => B(15), Ci => CTMP_15_port, S => 
                           S(15), Co => CTMP_16_port);
   FAI_17 : FA_1008 port map( A => A(16), B => B(16), Ci => CTMP_16_port, S => 
                           S(16), Co => CTMP_17_port);
   FAI_18 : FA_1007 port map( A => A(17), B => B(17), Ci => CTMP_17_port, S => 
                           S(17), Co => CTMP_18_port);
   FAI_19 : FA_1006 port map( A => A(18), B => B(18), Ci => CTMP_18_port, S => 
                           S(18), Co => CTMP_19_port);
   FAI_20 : FA_1005 port map( A => A(19), B => B(19), Ci => CTMP_19_port, S => 
                           S(19), Co => CTMP_20_port);
   FAI_21 : FA_1004 port map( A => A(20), B => B(20), Ci => CTMP_20_port, S => 
                           S(20), Co => CTMP_21_port);
   FAI_22 : FA_1003 port map( A => A(21), B => B(21), Ci => CTMP_21_port, S => 
                           S(21), Co => CTMP_22_port);
   FAI_23 : FA_1002 port map( A => A(22), B => B(22), Ci => CTMP_22_port, S => 
                           S(22), Co => CTMP_23_port);
   FAI_24 : FA_1001 port map( A => A(23), B => B(23), Ci => CTMP_23_port, S => 
                           S(23), Co => CTMP_24_port);
   FAI_25 : FA_1000 port map( A => A(24), B => B(24), Ci => CTMP_24_port, S => 
                           S(24), Co => CTMP_25_port);
   FAI_26 : FA_999 port map( A => A(25), B => B(25), Ci => CTMP_25_port, S => 
                           S(25), Co => CTMP_26_port);
   FAI_27 : FA_998 port map( A => A(26), B => B(26), Ci => CTMP_26_port, S => 
                           S(26), Co => CTMP_27_port);
   FAI_28 : FA_997 port map( A => A(27), B => B(27), Ci => CTMP_27_port, S => 
                           S(27), Co => CTMP_28_port);
   FAI_29 : FA_996 port map( A => A(28), B => B(28), Ci => CTMP_28_port, S => 
                           S(28), Co => CTMP_29_port);
   FAI_30 : FA_995 port map( A => A(29), B => B(29), Ci => CTMP_29_port, S => 
                           S(29), Co => CTMP_30_port);
   FAI_31 : FA_994 port map( A => A(30), B => B(30), Ci => CTMP_30_port, S => 
                           S(30), Co => CTMP_31_port);
   FAI_32 : FA_993 port map( A => A(31), B => B(31), Ci => CTMP_31_port, S => 
                           S(31), Co => CTMP_32_port);
   FAI_33 : FA_992 port map( A => A(32), B => B(32), Ci => CTMP_32_port, S => 
                           S(32), Co => CTMP_33_port);
   FAI_34 : FA_991 port map( A => A(33), B => B(33), Ci => CTMP_33_port, S => 
                           S(33), Co => CTMP_34_port);
   FAI_35 : FA_990 port map( A => A(34), B => B(34), Ci => CTMP_34_port, S => 
                           S(34), Co => CTMP_35_port);
   FAI_36 : FA_989 port map( A => A(35), B => B(35), Ci => CTMP_35_port, S => 
                           S(35), Co => CTMP_36_port);
   FAI_37 : FA_988 port map( A => A(36), B => B(36), Ci => CTMP_36_port, S => 
                           S(36), Co => CTMP_37_port);
   FAI_38 : FA_987 port map( A => A(37), B => B(37), Ci => CTMP_37_port, S => 
                           S(37), Co => CTMP_38_port);
   FAI_39 : FA_986 port map( A => A(38), B => B(38), Ci => CTMP_38_port, S => 
                           S(38), Co => CTMP_39_port);
   FAI_40 : FA_985 port map( A => A(39), B => B(39), Ci => CTMP_39_port, S => 
                           S(39), Co => CTMP_40_port);
   FAI_41 : FA_984 port map( A => A(40), B => B(40), Ci => CTMP_40_port, S => 
                           S(40), Co => CTMP_41_port);
   FAI_42 : FA_983 port map( A => A(41), B => B(41), Ci => CTMP_41_port, S => 
                           S(41), Co => CTMP_42_port);
   FAI_43 : FA_982 port map( A => A(42), B => B(42), Ci => CTMP_42_port, S => 
                           S(42), Co => CTMP_43_port);
   FAI_44 : FA_981 port map( A => A(43), B => B(43), Ci => CTMP_43_port, S => 
                           S(43), Co => CTMP_44_port);
   FAI_45 : FA_980 port map( A => A(44), B => B(44), Ci => CTMP_44_port, S => 
                           S(44), Co => CTMP_45_port);
   FAI_46 : FA_979 port map( A => A(45), B => B(45), Ci => CTMP_45_port, S => 
                           S(45), Co => CTMP_46_port);
   FAI_47 : FA_978 port map( A => A(46), B => B(46), Ci => CTMP_46_port, S => 
                           S(46), Co => CTMP_47_port);
   FAI_48 : FA_977 port map( A => A(47), B => B(47), Ci => CTMP_47_port, S => 
                           S(47), Co => CTMP_48_port);
   FAI_49 : FA_976 port map( A => A(48), B => B(48), Ci => CTMP_48_port, S => 
                           S(48), Co => CTMP_49_port);
   FAI_50 : FA_975 port map( A => A(49), B => B(49), Ci => CTMP_49_port, S => 
                           S(49), Co => CTMP_50_port);
   FAI_51 : FA_974 port map( A => A(50), B => B(50), Ci => CTMP_50_port, S => 
                           S(50), Co => CTMP_51_port);
   FAI_52 : FA_973 port map( A => A(51), B => B(51), Ci => CTMP_51_port, S => 
                           S(51), Co => CTMP_52_port);
   FAI_53 : FA_972 port map( A => A(52), B => B(52), Ci => CTMP_52_port, S => 
                           S(52), Co => CTMP_53_port);
   FAI_54 : FA_971 port map( A => A(53), B => B(53), Ci => CTMP_53_port, S => 
                           S(53), Co => CTMP_54_port);
   FAI_55 : FA_970 port map( A => A(54), B => B(54), Ci => CTMP_54_port, S => 
                           S(54), Co => CTMP_55_port);
   FAI_56 : FA_969 port map( A => A(55), B => B(55), Ci => CTMP_55_port, S => 
                           S(55), Co => CTMP_56_port);
   FAI_57 : FA_968 port map( A => A(56), B => B(56), Ci => CTMP_56_port, S => 
                           S(56), Co => CTMP_57_port);
   FAI_58 : FA_967 port map( A => A(57), B => B(57), Ci => CTMP_57_port, S => 
                           S(57), Co => CTMP_58_port);
   FAI_59 : FA_966 port map( A => A(58), B => B(58), Ci => CTMP_58_port, S => 
                           S(58), Co => CTMP_59_port);
   FAI_60 : FA_965 port map( A => A(59), B => B(59), Ci => CTMP_59_port, S => 
                           S(59), Co => CTMP_60_port);
   FAI_61 : FA_964 port map( A => A(60), B => B(60), Ci => CTMP_60_port, S => 
                           S(60), Co => CTMP_61_port);
   FAI_62 : FA_963 port map( A => A(61), B => B(61), Ci => CTMP_61_port, S => 
                           S(61), Co => CTMP_62_port);
   FAI_63 : FA_962 port map( A => A(62), B => B(62), Ci => CTMP_62_port, S => 
                           S(62), Co => CTMP_63_port);
   FAI_64 : FA_961 port map( A => A(63), B => B(63), Ci => CTMP_63_port, S => 
                           S(63), Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity IV_0 is

   port( A : in std_logic;  Y : out std_logic);

end IV_0;

architecture SYN_BEHAVIORAL of IV_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL.all;

entity BOOTHMUL is

   port( A, B : in std_logic_vector (31 downto 0);  P : out std_logic_vector 
         (63 downto 0));

end BOOTHMUL;

architecture SYN_STRUCTURAL of BOOTHMUL is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component RCA_NbitRca64_1
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NbitRca64_2
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NbitRca64_3
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NbitRca64_4
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NbitRca64_5
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NbitRca64_6
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NbitRca64_7
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NbitRca64_8
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NbitRca64_9
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NbitRca64_10
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NbitRca64_11
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NbitRca64_12
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NbitRca64_13
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NbitRca64_14
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NbitRca64_15
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component MUX51_MuxNbit64_1
      port( zeroSignal, A_signal, A_neg, A_shifted, A_neg_shifted : in 
            std_logic_vector (63 downto 0);  Sel : in std_logic_vector (2 
            downto 0);  Y : out std_logic_vector (63 downto 0));
   end component;
   
   component encoder_1
      port( pieceofB : in std_logic_vector (2 downto 0);  sel : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component MUX51_MuxNbit64_2
      port( zeroSignal, A_signal, A_neg, A_shifted, A_neg_shifted : in 
            std_logic_vector (63 downto 0);  Sel : in std_logic_vector (2 
            downto 0);  Y : out std_logic_vector (63 downto 0));
   end component;
   
   component encoder_2
      port( pieceofB : in std_logic_vector (2 downto 0);  sel : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component MUX51_MuxNbit64_3
      port( zeroSignal, A_signal, A_neg, A_shifted, A_neg_shifted : in 
            std_logic_vector (63 downto 0);  Sel : in std_logic_vector (2 
            downto 0);  Y : out std_logic_vector (63 downto 0));
   end component;
   
   component encoder_3
      port( pieceofB : in std_logic_vector (2 downto 0);  sel : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component MUX51_MuxNbit64_4
      port( zeroSignal, A_signal, A_neg, A_shifted, A_neg_shifted : in 
            std_logic_vector (63 downto 0);  Sel : in std_logic_vector (2 
            downto 0);  Y : out std_logic_vector (63 downto 0));
   end component;
   
   component encoder_4
      port( pieceofB : in std_logic_vector (2 downto 0);  sel : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component MUX51_MuxNbit64_5
      port( zeroSignal, A_signal, A_neg, A_shifted, A_neg_shifted : in 
            std_logic_vector (63 downto 0);  Sel : in std_logic_vector (2 
            downto 0);  Y : out std_logic_vector (63 downto 0));
   end component;
   
   component encoder_5
      port( pieceofB : in std_logic_vector (2 downto 0);  sel : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component MUX51_MuxNbit64_6
      port( zeroSignal, A_signal, A_neg, A_shifted, A_neg_shifted : in 
            std_logic_vector (63 downto 0);  Sel : in std_logic_vector (2 
            downto 0);  Y : out std_logic_vector (63 downto 0));
   end component;
   
   component encoder_6
      port( pieceofB : in std_logic_vector (2 downto 0);  sel : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component MUX51_MuxNbit64_7
      port( zeroSignal, A_signal, A_neg, A_shifted, A_neg_shifted : in 
            std_logic_vector (63 downto 0);  Sel : in std_logic_vector (2 
            downto 0);  Y : out std_logic_vector (63 downto 0));
   end component;
   
   component encoder_7
      port( pieceofB : in std_logic_vector (2 downto 0);  sel : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component MUX51_MuxNbit64_8
      port( zeroSignal, A_signal, A_neg, A_shifted, A_neg_shifted : in 
            std_logic_vector (63 downto 0);  Sel : in std_logic_vector (2 
            downto 0);  Y : out std_logic_vector (63 downto 0));
   end component;
   
   component encoder_8
      port( pieceofB : in std_logic_vector (2 downto 0);  sel : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component MUX51_MuxNbit64_9
      port( zeroSignal, A_signal, A_neg, A_shifted, A_neg_shifted : in 
            std_logic_vector (63 downto 0);  Sel : in std_logic_vector (2 
            downto 0);  Y : out std_logic_vector (63 downto 0));
   end component;
   
   component encoder_9
      port( pieceofB : in std_logic_vector (2 downto 0);  sel : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component MUX51_MuxNbit64_10
      port( zeroSignal, A_signal, A_neg, A_shifted, A_neg_shifted : in 
            std_logic_vector (63 downto 0);  Sel : in std_logic_vector (2 
            downto 0);  Y : out std_logic_vector (63 downto 0));
   end component;
   
   component encoder_10
      port( pieceofB : in std_logic_vector (2 downto 0);  sel : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component MUX51_MuxNbit64_11
      port( zeroSignal, A_signal, A_neg, A_shifted, A_neg_shifted : in 
            std_logic_vector (63 downto 0);  Sel : in std_logic_vector (2 
            downto 0);  Y : out std_logic_vector (63 downto 0));
   end component;
   
   component encoder_11
      port( pieceofB : in std_logic_vector (2 downto 0);  sel : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component MUX51_MuxNbit64_12
      port( zeroSignal, A_signal, A_neg, A_shifted, A_neg_shifted : in 
            std_logic_vector (63 downto 0);  Sel : in std_logic_vector (2 
            downto 0);  Y : out std_logic_vector (63 downto 0));
   end component;
   
   component encoder_12
      port( pieceofB : in std_logic_vector (2 downto 0);  sel : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component MUX51_MuxNbit64_13
      port( zeroSignal, A_signal, A_neg, A_shifted, A_neg_shifted : in 
            std_logic_vector (63 downto 0);  Sel : in std_logic_vector (2 
            downto 0);  Y : out std_logic_vector (63 downto 0));
   end component;
   
   component encoder_13
      port( pieceofB : in std_logic_vector (2 downto 0);  sel : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component MUX51_MuxNbit64_14
      port( zeroSignal, A_signal, A_neg, A_shifted, A_neg_shifted : in 
            std_logic_vector (63 downto 0);  Sel : in std_logic_vector (2 
            downto 0);  Y : out std_logic_vector (63 downto 0));
   end component;
   
   component encoder_14
      port( pieceofB : in std_logic_vector (2 downto 0);  sel : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component MUX51_MuxNbit64_15
      port( zeroSignal, A_signal, A_neg, A_shifted, A_neg_shifted : in 
            std_logic_vector (63 downto 0);  Sel : in std_logic_vector (2 
            downto 0);  Y : out std_logic_vector (63 downto 0));
   end component;
   
   component encoder_15
      port( pieceofB : in std_logic_vector (2 downto 0);  sel : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component MUX51_MuxNbit64_0
      port( zeroSignal, A_signal, A_neg, A_shifted, A_neg_shifted : in 
            std_logic_vector (63 downto 0);  Sel : in std_logic_vector (2 
            downto 0);  Y : out std_logic_vector (63 downto 0));
   end component;
   
   component encoder_0
      port( pieceofB : in std_logic_vector (2 downto 0);  sel : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_1
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_2
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_3
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_4
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_5
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_6
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_7
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_8
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_9
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_10
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_11
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_12
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_13
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_14
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_15
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_16
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_17
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_18
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_19
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_20
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_21
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_22
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_23
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_24
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_25
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_26
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_27
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_28
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_29
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_30
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_31
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_32
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_33
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_34
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_35
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_36
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_37
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_38
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_39
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_40
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_41
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_42
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_43
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_44
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_45
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_46
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_47
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_48
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_49
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_50
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_51
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_52
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_53
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_54
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_55
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_56
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_57
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_58
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_59
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_60
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_61
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_62
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_0
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component RCA_NbitRca64_0
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component IV_1
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_3
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_4
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_5
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_6
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_7
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_8
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_9
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_10
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_11
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_12
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_13
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_14
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_15
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_16
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_17
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_18
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_19
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_20
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_21
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_22
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_23
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_24
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_25
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_26
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_27
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_28
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_29
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_30
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_31
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_32
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_33
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_34
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_35
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_36
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_37
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_38
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_39
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_40
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_41
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_42
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_43
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_44
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_45
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_46
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_47
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_48
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_49
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_50
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_51
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_52
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_53
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_54
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_55
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_56
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_57
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_58
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_59
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_60
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_61
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_62
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_63
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_0
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, A_complement_63_port, 
      A_complement_62_port, A_complement_61_port, A_complement_60_port, 
      A_complement_59_port, A_complement_58_port, A_complement_57_port, 
      A_complement_56_port, A_complement_55_port, A_complement_54_port, 
      A_complement_53_port, A_complement_52_port, A_complement_51_port, 
      A_complement_50_port, A_complement_49_port, A_complement_48_port, 
      A_complement_47_port, A_complement_46_port, A_complement_45_port, 
      A_complement_44_port, A_complement_43_port, A_complement_42_port, 
      A_complement_41_port, A_complement_40_port, A_complement_39_port, 
      A_complement_38_port, A_complement_37_port, A_complement_36_port, 
      A_complement_35_port, A_complement_34_port, A_complement_33_port, 
      A_complement_32_port, A_complement_31_port, A_complement_30_port, 
      A_complement_29_port, A_complement_28_port, A_complement_27_port, 
      A_complement_26_port, A_complement_25_port, A_complement_24_port, 
      A_complement_23_port, A_complement_22_port, A_complement_21_port, 
      A_complement_20_port, A_complement_19_port, A_complement_18_port, 
      A_complement_17_port, A_complement_16_port, A_complement_15_port, 
      A_complement_14_port, A_complement_13_port, A_complement_12_port, 
      A_complement_11_port, A_complement_10_port, A_complement_9_port, 
      A_complement_8_port, A_complement_7_port, A_complement_6_port, 
      A_complement_5_port, A_complement_4_port, A_complement_3_port, 
      A_complement_2_port, A_complement_1_port, A_complement_0_port, 
      negative_inputs_0_63_port, negative_inputs_0_62_port, 
      negative_inputs_0_61_port, negative_inputs_0_60_port, 
      negative_inputs_0_59_port, negative_inputs_0_58_port, 
      negative_inputs_0_57_port, negative_inputs_0_56_port, 
      negative_inputs_0_55_port, negative_inputs_0_54_port, 
      negative_inputs_0_53_port, negative_inputs_0_52_port, 
      negative_inputs_0_51_port, negative_inputs_0_50_port, 
      negative_inputs_0_49_port, negative_inputs_0_48_port, 
      negative_inputs_0_47_port, negative_inputs_0_46_port, 
      negative_inputs_0_45_port, negative_inputs_0_44_port, 
      negative_inputs_0_43_port, negative_inputs_0_42_port, 
      negative_inputs_0_41_port, negative_inputs_0_40_port, 
      negative_inputs_0_39_port, negative_inputs_0_38_port, 
      negative_inputs_0_37_port, negative_inputs_0_36_port, 
      negative_inputs_0_35_port, negative_inputs_0_34_port, 
      negative_inputs_0_33_port, negative_inputs_0_32_port, 
      negative_inputs_0_31_port, negative_inputs_0_30_port, 
      negative_inputs_0_29_port, negative_inputs_0_28_port, 
      negative_inputs_0_27_port, negative_inputs_0_26_port, 
      negative_inputs_0_25_port, negative_inputs_0_24_port, 
      negative_inputs_0_23_port, negative_inputs_0_22_port, 
      negative_inputs_0_21_port, negative_inputs_0_20_port, 
      negative_inputs_0_19_port, negative_inputs_0_18_port, 
      negative_inputs_0_17_port, negative_inputs_0_16_port, 
      negative_inputs_0_15_port, negative_inputs_0_14_port, 
      negative_inputs_0_13_port, negative_inputs_0_12_port, 
      negative_inputs_0_11_port, negative_inputs_0_10_port, 
      negative_inputs_0_9_port, negative_inputs_0_8_port, 
      negative_inputs_0_7_port, negative_inputs_0_6_port, 
      negative_inputs_0_5_port, negative_inputs_0_4_port, 
      negative_inputs_0_3_port, negative_inputs_0_2_port, 
      negative_inputs_0_1_port, negative_inputs_0_0_port, 
      positive_inputs_8_63_port, positive_inputs_8_62_port, 
      positive_inputs_8_61_port, positive_inputs_8_60_port, 
      positive_inputs_8_59_port, positive_inputs_8_58_port, 
      positive_inputs_8_57_port, positive_inputs_8_56_port, 
      positive_inputs_8_55_port, positive_inputs_8_54_port, 
      positive_inputs_8_53_port, positive_inputs_8_52_port, 
      positive_inputs_8_51_port, positive_inputs_8_50_port, 
      positive_inputs_8_49_port, positive_inputs_8_48_port, 
      positive_inputs_8_47_port, positive_inputs_8_46_port, 
      positive_inputs_8_45_port, positive_inputs_8_44_port, 
      positive_inputs_8_43_port, positive_inputs_8_42_port, 
      positive_inputs_8_41_port, positive_inputs_8_40_port, 
      positive_inputs_8_39_port, positive_inputs_8_38_port, 
      positive_inputs_8_37_port, positive_inputs_8_36_port, 
      positive_inputs_8_35_port, positive_inputs_8_34_port, 
      positive_inputs_8_33_port, positive_inputs_8_32_port, 
      positive_inputs_8_31_port, positive_inputs_8_30_port, 
      positive_inputs_8_29_port, positive_inputs_8_28_port, 
      positive_inputs_8_27_port, positive_inputs_8_26_port, 
      positive_inputs_8_25_port, positive_inputs_8_24_port, 
      positive_inputs_8_23_port, positive_inputs_8_22_port, 
      positive_inputs_8_21_port, positive_inputs_8_20_port, 
      positive_inputs_8_19_port, positive_inputs_8_18_port, 
      positive_inputs_8_17_port, positive_inputs_8_16_port, 
      positive_inputs_8_15_port, positive_inputs_8_14_port, 
      positive_inputs_8_13_port, positive_inputs_8_12_port, 
      positive_inputs_8_11_port, positive_inputs_8_10_port, 
      positive_inputs_8_9_port, positive_inputs_8_8_port, 
      positive_inputs_8_7_port, positive_inputs_8_6_port, 
      positive_inputs_8_5_port, positive_inputs_8_4_port, 
      positive_inputs_8_3_port, positive_inputs_8_2_port, 
      positive_inputs_8_1_port, positive_inputs_7_63_port, 
      positive_inputs_7_62_port, positive_inputs_7_61_port, 
      positive_inputs_7_60_port, positive_inputs_7_59_port, 
      positive_inputs_7_58_port, positive_inputs_7_57_port, 
      positive_inputs_7_56_port, positive_inputs_7_55_port, 
      positive_inputs_7_54_port, positive_inputs_7_53_port, 
      positive_inputs_7_52_port, positive_inputs_7_51_port, 
      positive_inputs_7_50_port, positive_inputs_7_49_port, 
      positive_inputs_7_48_port, positive_inputs_7_47_port, 
      positive_inputs_7_46_port, positive_inputs_7_45_port, 
      positive_inputs_7_44_port, positive_inputs_7_43_port, 
      positive_inputs_7_42_port, positive_inputs_7_41_port, 
      positive_inputs_7_40_port, positive_inputs_7_39_port, 
      positive_inputs_7_38_port, positive_inputs_7_37_port, 
      positive_inputs_7_36_port, positive_inputs_7_35_port, 
      positive_inputs_7_34_port, positive_inputs_7_33_port, 
      positive_inputs_7_32_port, positive_inputs_7_31_port, 
      positive_inputs_7_30_port, positive_inputs_7_29_port, 
      positive_inputs_7_28_port, positive_inputs_7_27_port, 
      positive_inputs_7_26_port, positive_inputs_7_25_port, 
      positive_inputs_7_24_port, positive_inputs_7_23_port, 
      positive_inputs_7_22_port, positive_inputs_7_21_port, 
      positive_inputs_7_20_port, positive_inputs_7_19_port, 
      positive_inputs_7_18_port, positive_inputs_7_17_port, 
      positive_inputs_7_16_port, positive_inputs_7_15_port, 
      positive_inputs_7_14_port, positive_inputs_7_13_port, 
      positive_inputs_7_12_port, positive_inputs_7_11_port, 
      positive_inputs_7_10_port, positive_inputs_7_9_port, 
      positive_inputs_7_8_port, positive_inputs_7_7_port, 
      positive_inputs_7_6_port, positive_inputs_7_5_port, 
      positive_inputs_7_4_port, positive_inputs_7_3_port, 
      positive_inputs_7_2_port, positive_inputs_7_1_port, 
      positive_inputs_6_63_port, positive_inputs_6_62_port, 
      positive_inputs_6_61_port, positive_inputs_6_60_port, 
      positive_inputs_6_59_port, positive_inputs_6_58_port, 
      positive_inputs_6_57_port, positive_inputs_6_56_port, 
      positive_inputs_6_55_port, positive_inputs_6_54_port, 
      positive_inputs_6_53_port, positive_inputs_6_52_port, 
      positive_inputs_6_51_port, positive_inputs_6_50_port, 
      positive_inputs_6_49_port, positive_inputs_6_48_port, 
      positive_inputs_6_47_port, positive_inputs_6_46_port, 
      positive_inputs_6_45_port, positive_inputs_6_44_port, 
      positive_inputs_6_43_port, positive_inputs_6_42_port, 
      positive_inputs_6_41_port, positive_inputs_6_40_port, 
      positive_inputs_6_39_port, positive_inputs_6_38_port, 
      positive_inputs_6_37_port, positive_inputs_6_36_port, 
      positive_inputs_6_35_port, positive_inputs_6_34_port, 
      positive_inputs_6_33_port, positive_inputs_6_32_port, 
      positive_inputs_6_31_port, positive_inputs_6_30_port, 
      positive_inputs_6_29_port, positive_inputs_6_28_port, 
      positive_inputs_6_27_port, positive_inputs_6_26_port, 
      positive_inputs_6_25_port, positive_inputs_6_24_port, 
      positive_inputs_6_23_port, positive_inputs_6_22_port, 
      positive_inputs_6_21_port, positive_inputs_6_20_port, 
      positive_inputs_6_19_port, positive_inputs_6_18_port, 
      positive_inputs_6_17_port, positive_inputs_6_16_port, 
      positive_inputs_6_15_port, positive_inputs_6_14_port, 
      positive_inputs_6_13_port, positive_inputs_6_12_port, 
      positive_inputs_6_11_port, positive_inputs_6_10_port, 
      positive_inputs_6_9_port, positive_inputs_6_8_port, 
      positive_inputs_6_7_port, positive_inputs_6_6_port, 
      positive_inputs_6_5_port, positive_inputs_6_4_port, 
      positive_inputs_6_3_port, positive_inputs_6_2_port, 
      positive_inputs_6_1_port, positive_inputs_5_63_port, 
      positive_inputs_5_62_port, positive_inputs_5_61_port, 
      positive_inputs_5_60_port, positive_inputs_5_59_port, 
      positive_inputs_5_58_port, positive_inputs_5_57_port, 
      positive_inputs_5_56_port, positive_inputs_5_55_port, 
      positive_inputs_5_54_port, positive_inputs_5_53_port, 
      positive_inputs_5_52_port, positive_inputs_5_51_port, 
      positive_inputs_5_50_port, positive_inputs_5_49_port, 
      positive_inputs_5_48_port, positive_inputs_5_47_port, 
      positive_inputs_5_46_port, positive_inputs_5_45_port, 
      positive_inputs_5_44_port, positive_inputs_5_43_port, 
      positive_inputs_5_42_port, positive_inputs_5_41_port, 
      positive_inputs_5_40_port, positive_inputs_5_39_port, 
      positive_inputs_5_38_port, positive_inputs_5_37_port, 
      positive_inputs_5_36_port, positive_inputs_5_35_port, 
      positive_inputs_5_34_port, positive_inputs_5_33_port, 
      positive_inputs_5_32_port, positive_inputs_5_31_port, 
      positive_inputs_5_30_port, positive_inputs_5_29_port, 
      positive_inputs_5_28_port, positive_inputs_5_27_port, 
      positive_inputs_5_26_port, positive_inputs_5_25_port, 
      positive_inputs_5_24_port, positive_inputs_5_23_port, 
      positive_inputs_5_22_port, positive_inputs_5_21_port, 
      positive_inputs_5_20_port, positive_inputs_5_19_port, 
      positive_inputs_5_18_port, positive_inputs_5_17_port, 
      positive_inputs_5_16_port, positive_inputs_5_15_port, 
      positive_inputs_5_14_port, positive_inputs_5_13_port, 
      positive_inputs_5_12_port, positive_inputs_5_11_port, 
      positive_inputs_5_10_port, positive_inputs_5_9_port, 
      positive_inputs_5_8_port, positive_inputs_5_7_port, 
      positive_inputs_5_6_port, positive_inputs_5_5_port, 
      positive_inputs_5_4_port, positive_inputs_5_3_port, 
      positive_inputs_5_2_port, positive_inputs_5_1_port, 
      positive_inputs_4_63_port, positive_inputs_4_62_port, 
      positive_inputs_4_61_port, positive_inputs_4_60_port, 
      positive_inputs_4_59_port, positive_inputs_4_58_port, 
      positive_inputs_4_57_port, positive_inputs_4_56_port, 
      positive_inputs_4_55_port, positive_inputs_4_54_port, 
      positive_inputs_4_53_port, positive_inputs_4_52_port, 
      positive_inputs_4_51_port, positive_inputs_4_50_port, 
      positive_inputs_4_49_port, positive_inputs_4_48_port, 
      positive_inputs_4_47_port, positive_inputs_4_46_port, 
      positive_inputs_4_45_port, positive_inputs_4_44_port, 
      positive_inputs_4_43_port, positive_inputs_4_42_port, 
      positive_inputs_4_41_port, positive_inputs_4_40_port, 
      positive_inputs_4_39_port, positive_inputs_4_38_port, 
      positive_inputs_4_37_port, positive_inputs_4_36_port, 
      positive_inputs_4_35_port, positive_inputs_4_34_port, 
      positive_inputs_4_33_port, positive_inputs_4_32_port, 
      positive_inputs_4_31_port, positive_inputs_4_30_port, 
      positive_inputs_4_29_port, positive_inputs_4_28_port, 
      positive_inputs_4_27_port, positive_inputs_4_26_port, 
      positive_inputs_4_25_port, positive_inputs_4_24_port, 
      positive_inputs_4_23_port, positive_inputs_4_22_port, 
      positive_inputs_4_21_port, positive_inputs_4_20_port, 
      positive_inputs_4_19_port, positive_inputs_4_18_port, 
      positive_inputs_4_17_port, positive_inputs_4_16_port, 
      positive_inputs_4_15_port, positive_inputs_4_14_port, 
      positive_inputs_4_13_port, positive_inputs_4_12_port, 
      positive_inputs_4_11_port, positive_inputs_4_10_port, 
      positive_inputs_4_9_port, positive_inputs_4_8_port, 
      positive_inputs_4_7_port, positive_inputs_4_6_port, 
      positive_inputs_4_5_port, positive_inputs_4_4_port, 
      positive_inputs_4_3_port, positive_inputs_4_2_port, 
      positive_inputs_4_1_port, positive_inputs_3_63_port, 
      positive_inputs_3_62_port, positive_inputs_3_61_port, 
      positive_inputs_3_60_port, positive_inputs_3_59_port, 
      positive_inputs_3_58_port, positive_inputs_3_57_port, 
      positive_inputs_3_56_port, positive_inputs_3_55_port, 
      positive_inputs_3_54_port, positive_inputs_3_53_port, 
      positive_inputs_3_52_port, positive_inputs_3_51_port, 
      positive_inputs_3_50_port, positive_inputs_3_49_port, 
      positive_inputs_3_48_port, positive_inputs_3_47_port, 
      positive_inputs_3_46_port, positive_inputs_3_45_port, 
      positive_inputs_3_44_port, positive_inputs_3_43_port, 
      positive_inputs_3_42_port, positive_inputs_3_41_port, 
      positive_inputs_3_40_port, positive_inputs_3_39_port, 
      positive_inputs_3_38_port, positive_inputs_3_37_port, 
      positive_inputs_3_36_port, positive_inputs_3_35_port, 
      positive_inputs_3_34_port, positive_inputs_3_33_port, 
      positive_inputs_3_32_port, positive_inputs_3_31_port, 
      positive_inputs_3_30_port, positive_inputs_3_29_port, 
      positive_inputs_3_28_port, positive_inputs_3_27_port, 
      positive_inputs_3_26_port, positive_inputs_3_25_port, 
      positive_inputs_3_24_port, positive_inputs_3_23_port, 
      positive_inputs_3_22_port, positive_inputs_3_21_port, 
      positive_inputs_3_20_port, positive_inputs_3_19_port, 
      positive_inputs_3_18_port, positive_inputs_3_17_port, 
      positive_inputs_3_16_port, positive_inputs_3_15_port, 
      positive_inputs_3_14_port, positive_inputs_3_13_port, 
      positive_inputs_3_12_port, positive_inputs_3_11_port, 
      positive_inputs_3_10_port, positive_inputs_3_9_port, 
      positive_inputs_3_8_port, positive_inputs_3_7_port, 
      positive_inputs_3_6_port, positive_inputs_3_5_port, 
      positive_inputs_3_4_port, positive_inputs_3_3_port, 
      positive_inputs_3_2_port, positive_inputs_3_1_port, 
      positive_inputs_2_63_port, positive_inputs_2_62_port, 
      positive_inputs_2_61_port, positive_inputs_2_60_port, 
      positive_inputs_2_59_port, positive_inputs_2_58_port, 
      positive_inputs_2_57_port, positive_inputs_2_56_port, 
      positive_inputs_2_55_port, positive_inputs_2_54_port, 
      positive_inputs_2_53_port, positive_inputs_2_52_port, 
      positive_inputs_2_51_port, positive_inputs_2_50_port, 
      positive_inputs_2_49_port, positive_inputs_2_48_port, 
      positive_inputs_2_47_port, positive_inputs_2_46_port, 
      positive_inputs_2_45_port, positive_inputs_2_44_port, 
      positive_inputs_2_43_port, positive_inputs_2_42_port, 
      positive_inputs_2_41_port, positive_inputs_2_40_port, 
      positive_inputs_2_39_port, positive_inputs_2_38_port, 
      positive_inputs_2_37_port, positive_inputs_2_36_port, 
      positive_inputs_2_35_port, positive_inputs_2_34_port, 
      positive_inputs_2_33_port, positive_inputs_2_32_port, 
      positive_inputs_2_31_port, positive_inputs_2_30_port, 
      positive_inputs_2_29_port, positive_inputs_2_28_port, 
      positive_inputs_2_27_port, positive_inputs_2_26_port, 
      positive_inputs_2_25_port, positive_inputs_2_24_port, 
      positive_inputs_2_23_port, positive_inputs_2_22_port, 
      positive_inputs_2_21_port, positive_inputs_2_20_port, 
      positive_inputs_2_19_port, positive_inputs_2_18_port, 
      positive_inputs_2_17_port, positive_inputs_2_16_port, 
      positive_inputs_2_15_port, positive_inputs_2_14_port, 
      positive_inputs_2_13_port, positive_inputs_2_12_port, 
      positive_inputs_2_11_port, positive_inputs_2_10_port, 
      positive_inputs_2_9_port, positive_inputs_2_8_port, 
      positive_inputs_2_7_port, positive_inputs_2_6_port, 
      positive_inputs_2_5_port, positive_inputs_2_4_port, 
      positive_inputs_2_3_port, positive_inputs_2_2_port, 
      positive_inputs_2_1_port, positive_inputs_1_63_port, 
      positive_inputs_1_62_port, positive_inputs_1_61_port, 
      positive_inputs_1_60_port, positive_inputs_1_59_port, 
      positive_inputs_1_58_port, positive_inputs_1_57_port, 
      positive_inputs_1_56_port, positive_inputs_1_55_port, 
      positive_inputs_1_54_port, positive_inputs_1_53_port, 
      positive_inputs_1_52_port, positive_inputs_1_51_port, 
      positive_inputs_1_50_port, positive_inputs_1_49_port, 
      positive_inputs_1_48_port, positive_inputs_1_47_port, 
      positive_inputs_1_46_port, positive_inputs_1_45_port, 
      positive_inputs_1_44_port, positive_inputs_1_43_port, 
      positive_inputs_1_42_port, positive_inputs_1_41_port, 
      positive_inputs_1_40_port, positive_inputs_1_39_port, 
      positive_inputs_1_38_port, positive_inputs_1_37_port, 
      positive_inputs_1_36_port, positive_inputs_1_35_port, 
      positive_inputs_1_34_port, positive_inputs_1_33_port, 
      positive_inputs_1_32_port, positive_inputs_1_31_port, 
      positive_inputs_1_30_port, positive_inputs_1_29_port, 
      positive_inputs_1_28_port, positive_inputs_1_27_port, 
      positive_inputs_1_26_port, positive_inputs_1_25_port, 
      positive_inputs_1_24_port, positive_inputs_1_23_port, 
      positive_inputs_1_22_port, positive_inputs_1_21_port, 
      positive_inputs_1_20_port, positive_inputs_1_19_port, 
      positive_inputs_1_18_port, positive_inputs_1_17_port, 
      positive_inputs_1_16_port, positive_inputs_1_15_port, 
      positive_inputs_1_14_port, positive_inputs_1_13_port, 
      positive_inputs_1_12_port, positive_inputs_1_11_port, 
      positive_inputs_1_10_port, positive_inputs_1_9_port, 
      positive_inputs_1_8_port, positive_inputs_1_7_port, 
      positive_inputs_1_6_port, positive_inputs_1_5_port, 
      positive_inputs_1_4_port, positive_inputs_1_3_port, 
      positive_inputs_1_2_port, positive_inputs_1_1_port, 
      positive_inputs_16_63_port, positive_inputs_16_62_port, 
      positive_inputs_16_61_port, positive_inputs_16_60_port, 
      positive_inputs_16_59_port, positive_inputs_16_58_port, 
      positive_inputs_16_57_port, positive_inputs_16_56_port, 
      positive_inputs_16_55_port, positive_inputs_16_54_port, 
      positive_inputs_16_53_port, positive_inputs_16_52_port, 
      positive_inputs_16_51_port, positive_inputs_16_50_port, 
      positive_inputs_16_49_port, positive_inputs_16_48_port, 
      positive_inputs_16_47_port, positive_inputs_16_46_port, 
      positive_inputs_16_45_port, positive_inputs_16_44_port, 
      positive_inputs_16_43_port, positive_inputs_16_42_port, 
      positive_inputs_16_41_port, positive_inputs_16_40_port, 
      positive_inputs_16_39_port, positive_inputs_16_38_port, 
      positive_inputs_16_37_port, positive_inputs_16_36_port, 
      positive_inputs_16_35_port, positive_inputs_16_34_port, 
      positive_inputs_16_33_port, positive_inputs_16_32_port, 
      positive_inputs_16_31_port, positive_inputs_16_30_port, 
      positive_inputs_16_29_port, positive_inputs_16_28_port, 
      positive_inputs_16_27_port, positive_inputs_16_26_port, 
      positive_inputs_16_25_port, positive_inputs_16_24_port, 
      positive_inputs_16_23_port, positive_inputs_16_22_port, 
      positive_inputs_16_21_port, positive_inputs_16_20_port, 
      positive_inputs_16_19_port, positive_inputs_16_18_port, 
      positive_inputs_16_17_port, positive_inputs_16_16_port, 
      positive_inputs_16_15_port, positive_inputs_16_14_port, 
      positive_inputs_16_13_port, positive_inputs_16_12_port, 
      positive_inputs_16_11_port, positive_inputs_16_10_port, 
      positive_inputs_16_9_port, positive_inputs_16_8_port, 
      positive_inputs_16_7_port, positive_inputs_16_6_port, 
      positive_inputs_16_5_port, positive_inputs_16_4_port, 
      positive_inputs_16_3_port, positive_inputs_16_2_port, 
      positive_inputs_16_1_port, positive_inputs_15_63_port, 
      positive_inputs_15_62_port, positive_inputs_15_61_port, 
      positive_inputs_15_60_port, positive_inputs_15_59_port, 
      positive_inputs_15_58_port, positive_inputs_15_57_port, 
      positive_inputs_15_56_port, positive_inputs_15_55_port, 
      positive_inputs_15_54_port, positive_inputs_15_53_port, 
      positive_inputs_15_52_port, positive_inputs_15_51_port, 
      positive_inputs_15_50_port, positive_inputs_15_49_port, 
      positive_inputs_15_48_port, positive_inputs_15_47_port, 
      positive_inputs_15_46_port, positive_inputs_15_45_port, 
      positive_inputs_15_44_port, positive_inputs_15_43_port, 
      positive_inputs_15_42_port, positive_inputs_15_41_port, 
      positive_inputs_15_40_port, positive_inputs_15_39_port, 
      positive_inputs_15_38_port, positive_inputs_15_37_port, 
      positive_inputs_15_36_port, positive_inputs_15_35_port, 
      positive_inputs_15_34_port, positive_inputs_15_33_port, 
      positive_inputs_15_32_port, positive_inputs_15_31_port, 
      positive_inputs_15_30_port, positive_inputs_15_29_port, 
      positive_inputs_15_28_port, positive_inputs_15_27_port, 
      positive_inputs_15_26_port, positive_inputs_15_25_port, 
      positive_inputs_15_24_port, positive_inputs_15_23_port, 
      positive_inputs_15_22_port, positive_inputs_15_21_port, 
      positive_inputs_15_20_port, positive_inputs_15_19_port, 
      positive_inputs_15_18_port, positive_inputs_15_17_port, 
      positive_inputs_15_16_port, positive_inputs_15_15_port, 
      positive_inputs_15_14_port, positive_inputs_15_13_port, 
      positive_inputs_15_12_port, positive_inputs_15_11_port, 
      positive_inputs_15_10_port, positive_inputs_15_9_port, 
      positive_inputs_15_8_port, positive_inputs_15_7_port, 
      positive_inputs_15_6_port, positive_inputs_15_5_port, 
      positive_inputs_15_4_port, positive_inputs_15_3_port, 
      positive_inputs_15_2_port, positive_inputs_15_1_port, 
      positive_inputs_14_63_port, positive_inputs_14_62_port, 
      positive_inputs_14_61_port, positive_inputs_14_60_port, 
      positive_inputs_14_59_port, positive_inputs_14_58_port, 
      positive_inputs_14_57_port, positive_inputs_14_56_port, 
      positive_inputs_14_55_port, positive_inputs_14_54_port, 
      positive_inputs_14_53_port, positive_inputs_14_52_port, 
      positive_inputs_14_51_port, positive_inputs_14_50_port, 
      positive_inputs_14_49_port, positive_inputs_14_48_port, 
      positive_inputs_14_47_port, positive_inputs_14_46_port, 
      positive_inputs_14_45_port, positive_inputs_14_44_port, 
      positive_inputs_14_43_port, positive_inputs_14_42_port, 
      positive_inputs_14_41_port, positive_inputs_14_40_port, 
      positive_inputs_14_39_port, positive_inputs_14_38_port, 
      positive_inputs_14_37_port, positive_inputs_14_36_port, 
      positive_inputs_14_35_port, positive_inputs_14_34_port, 
      positive_inputs_14_33_port, positive_inputs_14_32_port, 
      positive_inputs_14_31_port, positive_inputs_14_30_port, 
      positive_inputs_14_29_port, positive_inputs_14_28_port, 
      positive_inputs_14_27_port, positive_inputs_14_26_port, 
      positive_inputs_14_25_port, positive_inputs_14_24_port, 
      positive_inputs_14_23_port, positive_inputs_14_22_port, 
      positive_inputs_14_21_port, positive_inputs_14_20_port, 
      positive_inputs_14_19_port, positive_inputs_14_18_port, 
      positive_inputs_14_17_port, positive_inputs_14_16_port, 
      positive_inputs_14_15_port, positive_inputs_14_14_port, 
      positive_inputs_14_13_port, positive_inputs_14_12_port, 
      positive_inputs_14_11_port, positive_inputs_14_10_port, 
      positive_inputs_14_9_port, positive_inputs_14_8_port, 
      positive_inputs_14_7_port, positive_inputs_14_6_port, 
      positive_inputs_14_5_port, positive_inputs_14_4_port, 
      positive_inputs_14_3_port, positive_inputs_14_2_port, 
      positive_inputs_14_1_port, positive_inputs_13_63_port, 
      positive_inputs_13_62_port, positive_inputs_13_61_port, 
      positive_inputs_13_60_port, positive_inputs_13_59_port, 
      positive_inputs_13_58_port, positive_inputs_13_57_port, 
      positive_inputs_13_56_port, positive_inputs_13_55_port, 
      positive_inputs_13_54_port, positive_inputs_13_53_port, 
      positive_inputs_13_52_port, positive_inputs_13_51_port, 
      positive_inputs_13_50_port, positive_inputs_13_49_port, 
      positive_inputs_13_48_port, positive_inputs_13_47_port, 
      positive_inputs_13_46_port, positive_inputs_13_45_port, 
      positive_inputs_13_44_port, positive_inputs_13_43_port, 
      positive_inputs_13_42_port, positive_inputs_13_41_port, 
      positive_inputs_13_40_port, positive_inputs_13_39_port, 
      positive_inputs_13_38_port, positive_inputs_13_37_port, 
      positive_inputs_13_36_port, positive_inputs_13_35_port, 
      positive_inputs_13_34_port, positive_inputs_13_33_port, 
      positive_inputs_13_32_port, positive_inputs_13_31_port, 
      positive_inputs_13_30_port, positive_inputs_13_29_port, 
      positive_inputs_13_28_port, positive_inputs_13_27_port, 
      positive_inputs_13_26_port, positive_inputs_13_25_port, 
      positive_inputs_13_24_port, positive_inputs_13_23_port, 
      positive_inputs_13_22_port, positive_inputs_13_21_port, 
      positive_inputs_13_20_port, positive_inputs_13_19_port, 
      positive_inputs_13_18_port, positive_inputs_13_17_port, 
      positive_inputs_13_16_port, positive_inputs_13_15_port, 
      positive_inputs_13_14_port, positive_inputs_13_13_port, 
      positive_inputs_13_12_port, positive_inputs_13_11_port, 
      positive_inputs_13_10_port, positive_inputs_13_9_port, 
      positive_inputs_13_8_port, positive_inputs_13_7_port, 
      positive_inputs_13_6_port, positive_inputs_13_5_port, 
      positive_inputs_13_4_port, positive_inputs_13_3_port, 
      positive_inputs_13_2_port, positive_inputs_13_1_port, 
      positive_inputs_12_63_port, positive_inputs_12_62_port, 
      positive_inputs_12_61_port, positive_inputs_12_60_port, 
      positive_inputs_12_59_port, positive_inputs_12_58_port, 
      positive_inputs_12_57_port, positive_inputs_12_56_port, 
      positive_inputs_12_55_port, positive_inputs_12_54_port, 
      positive_inputs_12_53_port, positive_inputs_12_52_port, 
      positive_inputs_12_51_port, positive_inputs_12_50_port, 
      positive_inputs_12_49_port, positive_inputs_12_48_port, 
      positive_inputs_12_47_port, positive_inputs_12_46_port, 
      positive_inputs_12_45_port, positive_inputs_12_44_port, 
      positive_inputs_12_43_port, positive_inputs_12_42_port, 
      positive_inputs_12_41_port, positive_inputs_12_40_port, 
      positive_inputs_12_39_port, positive_inputs_12_38_port, 
      positive_inputs_12_37_port, positive_inputs_12_36_port, 
      positive_inputs_12_35_port, positive_inputs_12_34_port, 
      positive_inputs_12_33_port, positive_inputs_12_32_port, 
      positive_inputs_12_31_port, positive_inputs_12_30_port, 
      positive_inputs_12_29_port, positive_inputs_12_28_port, 
      positive_inputs_12_27_port, positive_inputs_12_26_port, 
      positive_inputs_12_25_port, positive_inputs_12_24_port, 
      positive_inputs_12_23_port, positive_inputs_12_22_port, 
      positive_inputs_12_21_port, positive_inputs_12_20_port, 
      positive_inputs_12_19_port, positive_inputs_12_18_port, 
      positive_inputs_12_17_port, positive_inputs_12_16_port, 
      positive_inputs_12_15_port, positive_inputs_12_14_port, 
      positive_inputs_12_13_port, positive_inputs_12_12_port, 
      positive_inputs_12_11_port, positive_inputs_12_10_port, 
      positive_inputs_12_9_port, positive_inputs_12_8_port, 
      positive_inputs_12_7_port, positive_inputs_12_6_port, 
      positive_inputs_12_5_port, positive_inputs_12_4_port, 
      positive_inputs_12_3_port, positive_inputs_12_2_port, 
      positive_inputs_12_1_port, positive_inputs_11_63_port, 
      positive_inputs_11_62_port, positive_inputs_11_61_port, 
      positive_inputs_11_60_port, positive_inputs_11_59_port, 
      positive_inputs_11_58_port, positive_inputs_11_57_port, 
      positive_inputs_11_56_port, positive_inputs_11_55_port, 
      positive_inputs_11_54_port, positive_inputs_11_53_port, 
      positive_inputs_11_52_port, positive_inputs_11_51_port, 
      positive_inputs_11_50_port, positive_inputs_11_49_port, 
      positive_inputs_11_48_port, positive_inputs_11_47_port, 
      positive_inputs_11_46_port, positive_inputs_11_45_port, 
      positive_inputs_11_44_port, positive_inputs_11_43_port, 
      positive_inputs_11_42_port, positive_inputs_11_41_port, 
      positive_inputs_11_40_port, positive_inputs_11_39_port, 
      positive_inputs_11_38_port, positive_inputs_11_37_port, 
      positive_inputs_11_36_port, positive_inputs_11_35_port, 
      positive_inputs_11_34_port, positive_inputs_11_33_port, 
      positive_inputs_11_32_port, positive_inputs_11_31_port, 
      positive_inputs_11_30_port, positive_inputs_11_29_port, 
      positive_inputs_11_28_port, positive_inputs_11_27_port, 
      positive_inputs_11_26_port, positive_inputs_11_25_port, 
      positive_inputs_11_24_port, positive_inputs_11_23_port, 
      positive_inputs_11_22_port, positive_inputs_11_21_port, 
      positive_inputs_11_20_port, positive_inputs_11_19_port, 
      positive_inputs_11_18_port, positive_inputs_11_17_port, 
      positive_inputs_11_16_port, positive_inputs_11_15_port, 
      positive_inputs_11_14_port, positive_inputs_11_13_port, 
      positive_inputs_11_12_port, positive_inputs_11_11_port, 
      positive_inputs_11_10_port, positive_inputs_11_9_port, 
      positive_inputs_11_8_port, positive_inputs_11_7_port, 
      positive_inputs_11_6_port, positive_inputs_11_5_port, 
      positive_inputs_11_4_port, positive_inputs_11_3_port, 
      positive_inputs_11_2_port, positive_inputs_11_1_port, 
      positive_inputs_10_63_port, positive_inputs_10_62_port, 
      positive_inputs_10_61_port, positive_inputs_10_60_port, 
      positive_inputs_10_59_port, positive_inputs_10_58_port, 
      positive_inputs_10_57_port, positive_inputs_10_56_port, 
      positive_inputs_10_55_port, positive_inputs_10_54_port, 
      positive_inputs_10_53_port, positive_inputs_10_52_port, 
      positive_inputs_10_51_port, positive_inputs_10_50_port, 
      positive_inputs_10_49_port, positive_inputs_10_48_port, 
      positive_inputs_10_47_port, positive_inputs_10_46_port, 
      positive_inputs_10_45_port, positive_inputs_10_44_port, 
      positive_inputs_10_43_port, positive_inputs_10_42_port, 
      positive_inputs_10_41_port, positive_inputs_10_40_port, 
      positive_inputs_10_39_port, positive_inputs_10_38_port, 
      positive_inputs_10_37_port, positive_inputs_10_36_port, 
      positive_inputs_10_35_port, positive_inputs_10_34_port, 
      positive_inputs_10_33_port, positive_inputs_10_32_port, 
      positive_inputs_10_31_port, positive_inputs_10_30_port, 
      positive_inputs_10_29_port, positive_inputs_10_28_port, 
      positive_inputs_10_27_port, positive_inputs_10_26_port, 
      positive_inputs_10_25_port, positive_inputs_10_24_port, 
      positive_inputs_10_23_port, positive_inputs_10_22_port, 
      positive_inputs_10_21_port, positive_inputs_10_20_port, 
      positive_inputs_10_19_port, positive_inputs_10_18_port, 
      positive_inputs_10_17_port, positive_inputs_10_16_port, 
      positive_inputs_10_15_port, positive_inputs_10_14_port, 
      positive_inputs_10_13_port, positive_inputs_10_12_port, 
      positive_inputs_10_11_port, positive_inputs_10_10_port, 
      positive_inputs_10_9_port, positive_inputs_10_8_port, 
      positive_inputs_10_7_port, positive_inputs_10_6_port, 
      positive_inputs_10_5_port, positive_inputs_10_4_port, 
      positive_inputs_10_3_port, positive_inputs_10_2_port, 
      positive_inputs_10_1_port, positive_inputs_9_63_port, 
      positive_inputs_9_62_port, positive_inputs_9_61_port, 
      positive_inputs_9_60_port, positive_inputs_9_59_port, 
      positive_inputs_9_58_port, positive_inputs_9_57_port, 
      positive_inputs_9_56_port, positive_inputs_9_55_port, 
      positive_inputs_9_54_port, positive_inputs_9_53_port, 
      positive_inputs_9_52_port, positive_inputs_9_51_port, 
      positive_inputs_9_50_port, positive_inputs_9_49_port, 
      positive_inputs_9_48_port, positive_inputs_9_47_port, 
      positive_inputs_9_46_port, positive_inputs_9_45_port, 
      positive_inputs_9_44_port, positive_inputs_9_43_port, 
      positive_inputs_9_42_port, positive_inputs_9_41_port, 
      positive_inputs_9_40_port, positive_inputs_9_39_port, 
      positive_inputs_9_38_port, positive_inputs_9_37_port, 
      positive_inputs_9_36_port, positive_inputs_9_35_port, 
      positive_inputs_9_34_port, positive_inputs_9_33_port, 
      positive_inputs_9_32_port, positive_inputs_9_31_port, 
      positive_inputs_9_30_port, positive_inputs_9_29_port, 
      positive_inputs_9_28_port, positive_inputs_9_27_port, 
      positive_inputs_9_26_port, positive_inputs_9_25_port, 
      positive_inputs_9_24_port, positive_inputs_9_23_port, 
      positive_inputs_9_22_port, positive_inputs_9_21_port, 
      positive_inputs_9_20_port, positive_inputs_9_19_port, 
      positive_inputs_9_18_port, positive_inputs_9_17_port, 
      positive_inputs_9_16_port, positive_inputs_9_15_port, 
      positive_inputs_9_14_port, positive_inputs_9_13_port, 
      positive_inputs_9_12_port, positive_inputs_9_11_port, 
      positive_inputs_9_10_port, positive_inputs_9_9_port, 
      positive_inputs_9_8_port, positive_inputs_9_7_port, 
      positive_inputs_9_6_port, positive_inputs_9_5_port, 
      positive_inputs_9_4_port, positive_inputs_9_3_port, 
      positive_inputs_9_2_port, positive_inputs_9_1_port, 
      positive_inputs_24_63_port, positive_inputs_24_62_port, 
      positive_inputs_24_61_port, positive_inputs_24_60_port, 
      positive_inputs_24_59_port, positive_inputs_24_58_port, 
      positive_inputs_24_57_port, positive_inputs_24_56_port, 
      positive_inputs_24_55_port, positive_inputs_24_54_port, 
      positive_inputs_24_53_port, positive_inputs_24_52_port, 
      positive_inputs_24_51_port, positive_inputs_24_50_port, 
      positive_inputs_24_49_port, positive_inputs_24_48_port, 
      positive_inputs_24_47_port, positive_inputs_24_46_port, 
      positive_inputs_24_45_port, positive_inputs_24_44_port, 
      positive_inputs_24_43_port, positive_inputs_24_42_port, 
      positive_inputs_24_41_port, positive_inputs_24_40_port, 
      positive_inputs_24_39_port, positive_inputs_24_38_port, 
      positive_inputs_24_37_port, positive_inputs_24_36_port, 
      positive_inputs_24_35_port, positive_inputs_24_34_port, 
      positive_inputs_24_33_port, positive_inputs_24_32_port, 
      positive_inputs_24_31_port, positive_inputs_24_30_port, 
      positive_inputs_24_29_port, positive_inputs_24_28_port, 
      positive_inputs_24_27_port, positive_inputs_24_26_port, 
      positive_inputs_24_25_port, positive_inputs_24_24_port, 
      positive_inputs_24_23_port, positive_inputs_24_22_port, 
      positive_inputs_24_21_port, positive_inputs_24_20_port, 
      positive_inputs_24_19_port, positive_inputs_24_18_port, 
      positive_inputs_24_17_port, positive_inputs_24_16_port, 
      positive_inputs_24_15_port, positive_inputs_24_14_port, 
      positive_inputs_24_13_port, positive_inputs_24_12_port, 
      positive_inputs_24_11_port, positive_inputs_24_10_port, 
      positive_inputs_24_9_port, positive_inputs_24_8_port, 
      positive_inputs_24_7_port, positive_inputs_24_6_port, 
      positive_inputs_24_5_port, positive_inputs_24_4_port, 
      positive_inputs_24_3_port, positive_inputs_24_2_port, 
      positive_inputs_24_1_port, positive_inputs_23_63_port, 
      positive_inputs_23_62_port, positive_inputs_23_61_port, 
      positive_inputs_23_60_port, positive_inputs_23_59_port, 
      positive_inputs_23_58_port, positive_inputs_23_57_port, 
      positive_inputs_23_56_port, positive_inputs_23_55_port, 
      positive_inputs_23_54_port, positive_inputs_23_53_port, 
      positive_inputs_23_52_port, positive_inputs_23_51_port, 
      positive_inputs_23_50_port, positive_inputs_23_49_port, 
      positive_inputs_23_48_port, positive_inputs_23_47_port, 
      positive_inputs_23_46_port, positive_inputs_23_45_port, 
      positive_inputs_23_44_port, positive_inputs_23_43_port, 
      positive_inputs_23_42_port, positive_inputs_23_41_port, 
      positive_inputs_23_40_port, positive_inputs_23_39_port, 
      positive_inputs_23_38_port, positive_inputs_23_37_port, 
      positive_inputs_23_36_port, positive_inputs_23_35_port, 
      positive_inputs_23_34_port, positive_inputs_23_33_port, 
      positive_inputs_23_32_port, positive_inputs_23_31_port, 
      positive_inputs_23_30_port, positive_inputs_23_29_port, 
      positive_inputs_23_28_port, positive_inputs_23_27_port, 
      positive_inputs_23_26_port, positive_inputs_23_25_port, 
      positive_inputs_23_24_port, positive_inputs_23_23_port, 
      positive_inputs_23_22_port, positive_inputs_23_21_port, 
      positive_inputs_23_20_port, positive_inputs_23_19_port, 
      positive_inputs_23_18_port, positive_inputs_23_17_port, 
      positive_inputs_23_16_port, positive_inputs_23_15_port, 
      positive_inputs_23_14_port, positive_inputs_23_13_port, 
      positive_inputs_23_12_port, positive_inputs_23_11_port, 
      positive_inputs_23_10_port, positive_inputs_23_9_port, 
      positive_inputs_23_8_port, positive_inputs_23_7_port, 
      positive_inputs_23_6_port, positive_inputs_23_5_port, 
      positive_inputs_23_4_port, positive_inputs_23_3_port, 
      positive_inputs_23_2_port, positive_inputs_23_1_port, 
      positive_inputs_22_63_port, positive_inputs_22_62_port, 
      positive_inputs_22_61_port, positive_inputs_22_60_port, 
      positive_inputs_22_59_port, positive_inputs_22_58_port, 
      positive_inputs_22_57_port, positive_inputs_22_56_port, 
      positive_inputs_22_55_port, positive_inputs_22_54_port, 
      positive_inputs_22_53_port, positive_inputs_22_52_port, 
      positive_inputs_22_51_port, positive_inputs_22_50_port, 
      positive_inputs_22_49_port, positive_inputs_22_48_port, 
      positive_inputs_22_47_port, positive_inputs_22_46_port, 
      positive_inputs_22_45_port, positive_inputs_22_44_port, 
      positive_inputs_22_43_port, positive_inputs_22_42_port, 
      positive_inputs_22_41_port, positive_inputs_22_40_port, 
      positive_inputs_22_39_port, positive_inputs_22_38_port, 
      positive_inputs_22_37_port, positive_inputs_22_36_port, 
      positive_inputs_22_35_port, positive_inputs_22_34_port, 
      positive_inputs_22_33_port, positive_inputs_22_32_port, 
      positive_inputs_22_31_port, positive_inputs_22_30_port, 
      positive_inputs_22_29_port, positive_inputs_22_28_port, 
      positive_inputs_22_27_port, positive_inputs_22_26_port, 
      positive_inputs_22_25_port, positive_inputs_22_24_port, 
      positive_inputs_22_23_port, positive_inputs_22_22_port, 
      positive_inputs_22_21_port, positive_inputs_22_20_port, 
      positive_inputs_22_19_port, positive_inputs_22_18_port, 
      positive_inputs_22_17_port, positive_inputs_22_16_port, 
      positive_inputs_22_15_port, positive_inputs_22_14_port, 
      positive_inputs_22_13_port, positive_inputs_22_12_port, 
      positive_inputs_22_11_port, positive_inputs_22_10_port, 
      positive_inputs_22_9_port, positive_inputs_22_8_port, 
      positive_inputs_22_7_port, positive_inputs_22_6_port, 
      positive_inputs_22_5_port, positive_inputs_22_4_port, 
      positive_inputs_22_3_port, positive_inputs_22_2_port, 
      positive_inputs_22_1_port, positive_inputs_21_63_port, 
      positive_inputs_21_62_port, positive_inputs_21_61_port, 
      positive_inputs_21_60_port, positive_inputs_21_59_port, 
      positive_inputs_21_58_port, positive_inputs_21_57_port, 
      positive_inputs_21_56_port, positive_inputs_21_55_port, 
      positive_inputs_21_54_port, positive_inputs_21_53_port, 
      positive_inputs_21_52_port, positive_inputs_21_51_port, 
      positive_inputs_21_50_port, positive_inputs_21_49_port, 
      positive_inputs_21_48_port, positive_inputs_21_47_port, 
      positive_inputs_21_46_port, positive_inputs_21_45_port, 
      positive_inputs_21_44_port, positive_inputs_21_43_port, 
      positive_inputs_21_42_port, positive_inputs_21_41_port, 
      positive_inputs_21_40_port, positive_inputs_21_39_port, 
      positive_inputs_21_38_port, positive_inputs_21_37_port, 
      positive_inputs_21_36_port, positive_inputs_21_35_port, 
      positive_inputs_21_34_port, positive_inputs_21_33_port, 
      positive_inputs_21_32_port, positive_inputs_21_31_port, 
      positive_inputs_21_30_port, positive_inputs_21_29_port, 
      positive_inputs_21_28_port, positive_inputs_21_27_port, 
      positive_inputs_21_26_port, positive_inputs_21_25_port, 
      positive_inputs_21_24_port, positive_inputs_21_23_port, 
      positive_inputs_21_22_port, positive_inputs_21_21_port, 
      positive_inputs_21_20_port, positive_inputs_21_19_port, 
      positive_inputs_21_18_port, positive_inputs_21_17_port, 
      positive_inputs_21_16_port, positive_inputs_21_15_port, 
      positive_inputs_21_14_port, positive_inputs_21_13_port, 
      positive_inputs_21_12_port, positive_inputs_21_11_port, 
      positive_inputs_21_10_port, positive_inputs_21_9_port, 
      positive_inputs_21_8_port, positive_inputs_21_7_port, 
      positive_inputs_21_6_port, positive_inputs_21_5_port, 
      positive_inputs_21_4_port, positive_inputs_21_3_port, 
      positive_inputs_21_2_port, positive_inputs_21_1_port, 
      positive_inputs_20_63_port, positive_inputs_20_62_port, 
      positive_inputs_20_61_port, positive_inputs_20_60_port, 
      positive_inputs_20_59_port, positive_inputs_20_58_port, 
      positive_inputs_20_57_port, positive_inputs_20_56_port, 
      positive_inputs_20_55_port, positive_inputs_20_54_port, 
      positive_inputs_20_53_port, positive_inputs_20_52_port, 
      positive_inputs_20_51_port, positive_inputs_20_50_port, 
      positive_inputs_20_49_port, positive_inputs_20_48_port, 
      positive_inputs_20_47_port, positive_inputs_20_46_port, 
      positive_inputs_20_45_port, positive_inputs_20_44_port, 
      positive_inputs_20_43_port, positive_inputs_20_42_port, 
      positive_inputs_20_41_port, positive_inputs_20_40_port, 
      positive_inputs_20_39_port, positive_inputs_20_38_port, 
      positive_inputs_20_37_port, positive_inputs_20_36_port, 
      positive_inputs_20_35_port, positive_inputs_20_34_port, 
      positive_inputs_20_33_port, positive_inputs_20_32_port, 
      positive_inputs_20_31_port, positive_inputs_20_30_port, 
      positive_inputs_20_29_port, positive_inputs_20_28_port, 
      positive_inputs_20_27_port, positive_inputs_20_26_port, 
      positive_inputs_20_25_port, positive_inputs_20_24_port, 
      positive_inputs_20_23_port, positive_inputs_20_22_port, 
      positive_inputs_20_21_port, positive_inputs_20_20_port, 
      positive_inputs_20_19_port, positive_inputs_20_18_port, 
      positive_inputs_20_17_port, positive_inputs_20_16_port, 
      positive_inputs_20_15_port, positive_inputs_20_14_port, 
      positive_inputs_20_13_port, positive_inputs_20_12_port, 
      positive_inputs_20_11_port, positive_inputs_20_10_port, 
      positive_inputs_20_9_port, positive_inputs_20_8_port, 
      positive_inputs_20_7_port, positive_inputs_20_6_port, 
      positive_inputs_20_5_port, positive_inputs_20_4_port, 
      positive_inputs_20_3_port, positive_inputs_20_2_port, 
      positive_inputs_20_1_port, positive_inputs_19_63_port, 
      positive_inputs_19_62_port, positive_inputs_19_61_port, 
      positive_inputs_19_60_port, positive_inputs_19_59_port, 
      positive_inputs_19_58_port, positive_inputs_19_57_port, 
      positive_inputs_19_56_port, positive_inputs_19_55_port, 
      positive_inputs_19_54_port, positive_inputs_19_53_port, 
      positive_inputs_19_52_port, positive_inputs_19_51_port, 
      positive_inputs_19_50_port, positive_inputs_19_49_port, 
      positive_inputs_19_48_port, positive_inputs_19_47_port, 
      positive_inputs_19_46_port, positive_inputs_19_45_port, 
      positive_inputs_19_44_port, positive_inputs_19_43_port, 
      positive_inputs_19_42_port, positive_inputs_19_41_port, 
      positive_inputs_19_40_port, positive_inputs_19_39_port, 
      positive_inputs_19_38_port, positive_inputs_19_37_port, 
      positive_inputs_19_36_port, positive_inputs_19_35_port, 
      positive_inputs_19_34_port, positive_inputs_19_33_port, 
      positive_inputs_19_32_port, positive_inputs_19_31_port, 
      positive_inputs_19_30_port, positive_inputs_19_29_port, 
      positive_inputs_19_28_port, positive_inputs_19_27_port, 
      positive_inputs_19_26_port, positive_inputs_19_25_port, 
      positive_inputs_19_24_port, positive_inputs_19_23_port, 
      positive_inputs_19_22_port, positive_inputs_19_21_port, 
      positive_inputs_19_20_port, positive_inputs_19_19_port, 
      positive_inputs_19_18_port, positive_inputs_19_17_port, 
      positive_inputs_19_16_port, positive_inputs_19_15_port, 
      positive_inputs_19_14_port, positive_inputs_19_13_port, 
      positive_inputs_19_12_port, positive_inputs_19_11_port, 
      positive_inputs_19_10_port, positive_inputs_19_9_port, 
      positive_inputs_19_8_port, positive_inputs_19_7_port, 
      positive_inputs_19_6_port, positive_inputs_19_5_port, 
      positive_inputs_19_4_port, positive_inputs_19_3_port, 
      positive_inputs_19_2_port, positive_inputs_19_1_port, 
      positive_inputs_18_63_port, positive_inputs_18_62_port, 
      positive_inputs_18_61_port, positive_inputs_18_60_port, 
      positive_inputs_18_59_port, positive_inputs_18_58_port, 
      positive_inputs_18_57_port, positive_inputs_18_56_port, 
      positive_inputs_18_55_port, positive_inputs_18_54_port, 
      positive_inputs_18_53_port, positive_inputs_18_52_port, 
      positive_inputs_18_51_port, positive_inputs_18_50_port, 
      positive_inputs_18_49_port, positive_inputs_18_48_port, 
      positive_inputs_18_47_port, positive_inputs_18_46_port, 
      positive_inputs_18_45_port, positive_inputs_18_44_port, 
      positive_inputs_18_43_port, positive_inputs_18_42_port, 
      positive_inputs_18_41_port, positive_inputs_18_40_port, 
      positive_inputs_18_39_port, positive_inputs_18_38_port, 
      positive_inputs_18_37_port, positive_inputs_18_36_port, 
      positive_inputs_18_35_port, positive_inputs_18_34_port, 
      positive_inputs_18_33_port, positive_inputs_18_32_port, 
      positive_inputs_18_31_port, positive_inputs_18_30_port, 
      positive_inputs_18_29_port, positive_inputs_18_28_port, 
      positive_inputs_18_27_port, positive_inputs_18_26_port, 
      positive_inputs_18_25_port, positive_inputs_18_24_port, 
      positive_inputs_18_23_port, positive_inputs_18_22_port, 
      positive_inputs_18_21_port, positive_inputs_18_20_port, 
      positive_inputs_18_19_port, positive_inputs_18_18_port, 
      positive_inputs_18_17_port, positive_inputs_18_16_port, 
      positive_inputs_18_15_port, positive_inputs_18_14_port, 
      positive_inputs_18_13_port, positive_inputs_18_12_port, 
      positive_inputs_18_11_port, positive_inputs_18_10_port, 
      positive_inputs_18_9_port, positive_inputs_18_8_port, 
      positive_inputs_18_7_port, positive_inputs_18_6_port, 
      positive_inputs_18_5_port, positive_inputs_18_4_port, 
      positive_inputs_18_3_port, positive_inputs_18_2_port, 
      positive_inputs_18_1_port, positive_inputs_17_63_port, 
      positive_inputs_17_62_port, positive_inputs_17_61_port, 
      positive_inputs_17_60_port, positive_inputs_17_59_port, 
      positive_inputs_17_58_port, positive_inputs_17_57_port, 
      positive_inputs_17_56_port, positive_inputs_17_55_port, 
      positive_inputs_17_54_port, positive_inputs_17_53_port, 
      positive_inputs_17_52_port, positive_inputs_17_51_port, 
      positive_inputs_17_50_port, positive_inputs_17_49_port, 
      positive_inputs_17_48_port, positive_inputs_17_47_port, 
      positive_inputs_17_46_port, positive_inputs_17_45_port, 
      positive_inputs_17_44_port, positive_inputs_17_43_port, 
      positive_inputs_17_42_port, positive_inputs_17_41_port, 
      positive_inputs_17_40_port, positive_inputs_17_39_port, 
      positive_inputs_17_38_port, positive_inputs_17_37_port, 
      positive_inputs_17_36_port, positive_inputs_17_35_port, 
      positive_inputs_17_34_port, positive_inputs_17_33_port, 
      positive_inputs_17_32_port, positive_inputs_17_31_port, 
      positive_inputs_17_30_port, positive_inputs_17_29_port, 
      positive_inputs_17_28_port, positive_inputs_17_27_port, 
      positive_inputs_17_26_port, positive_inputs_17_25_port, 
      positive_inputs_17_24_port, positive_inputs_17_23_port, 
      positive_inputs_17_22_port, positive_inputs_17_21_port, 
      positive_inputs_17_20_port, positive_inputs_17_19_port, 
      positive_inputs_17_18_port, positive_inputs_17_17_port, 
      positive_inputs_17_16_port, positive_inputs_17_15_port, 
      positive_inputs_17_14_port, positive_inputs_17_13_port, 
      positive_inputs_17_12_port, positive_inputs_17_11_port, 
      positive_inputs_17_10_port, positive_inputs_17_9_port, 
      positive_inputs_17_8_port, positive_inputs_17_7_port, 
      positive_inputs_17_6_port, positive_inputs_17_5_port, 
      positive_inputs_17_4_port, positive_inputs_17_3_port, 
      positive_inputs_17_2_port, positive_inputs_17_1_port, 
      positive_inputs_31_63_port, positive_inputs_31_62_port, 
      positive_inputs_31_61_port, positive_inputs_31_60_port, 
      positive_inputs_31_59_port, positive_inputs_31_58_port, 
      positive_inputs_31_57_port, positive_inputs_31_56_port, 
      positive_inputs_31_55_port, positive_inputs_31_54_port, 
      positive_inputs_31_53_port, positive_inputs_31_52_port, 
      positive_inputs_31_51_port, positive_inputs_31_50_port, 
      positive_inputs_31_49_port, positive_inputs_31_48_port, 
      positive_inputs_31_47_port, positive_inputs_31_46_port, 
      positive_inputs_31_45_port, positive_inputs_31_44_port, 
      positive_inputs_31_43_port, positive_inputs_31_42_port, 
      positive_inputs_31_41_port, positive_inputs_31_40_port, 
      positive_inputs_31_39_port, positive_inputs_31_38_port, 
      positive_inputs_31_37_port, positive_inputs_31_36_port, 
      positive_inputs_31_35_port, positive_inputs_31_34_port, 
      positive_inputs_31_33_port, positive_inputs_31_32_port, 
      positive_inputs_31_31_port, positive_inputs_31_30_port, 
      positive_inputs_31_29_port, positive_inputs_31_28_port, 
      positive_inputs_31_27_port, positive_inputs_31_26_port, 
      positive_inputs_31_25_port, positive_inputs_31_24_port, 
      positive_inputs_31_23_port, positive_inputs_31_22_port, 
      positive_inputs_31_21_port, positive_inputs_31_20_port, 
      positive_inputs_31_19_port, positive_inputs_31_18_port, 
      positive_inputs_31_17_port, positive_inputs_31_16_port, 
      positive_inputs_31_15_port, positive_inputs_31_14_port, 
      positive_inputs_31_13_port, positive_inputs_31_12_port, 
      positive_inputs_31_11_port, positive_inputs_31_10_port, 
      positive_inputs_31_9_port, positive_inputs_31_8_port, 
      positive_inputs_31_7_port, positive_inputs_31_6_port, 
      positive_inputs_31_5_port, positive_inputs_31_4_port, 
      positive_inputs_31_3_port, positive_inputs_31_2_port, 
      positive_inputs_31_1_port, positive_inputs_30_63_port, 
      positive_inputs_30_62_port, positive_inputs_30_61_port, 
      positive_inputs_30_60_port, positive_inputs_30_59_port, 
      positive_inputs_30_58_port, positive_inputs_30_57_port, 
      positive_inputs_30_56_port, positive_inputs_30_55_port, 
      positive_inputs_30_54_port, positive_inputs_30_53_port, 
      positive_inputs_30_52_port, positive_inputs_30_51_port, 
      positive_inputs_30_50_port, positive_inputs_30_49_port, 
      positive_inputs_30_48_port, positive_inputs_30_47_port, 
      positive_inputs_30_46_port, positive_inputs_30_45_port, 
      positive_inputs_30_44_port, positive_inputs_30_43_port, 
      positive_inputs_30_42_port, positive_inputs_30_41_port, 
      positive_inputs_30_40_port, positive_inputs_30_39_port, 
      positive_inputs_30_38_port, positive_inputs_30_37_port, 
      positive_inputs_30_36_port, positive_inputs_30_35_port, 
      positive_inputs_30_34_port, positive_inputs_30_33_port, 
      positive_inputs_30_32_port, positive_inputs_30_31_port, 
      positive_inputs_30_30_port, positive_inputs_30_29_port, 
      positive_inputs_30_28_port, positive_inputs_30_27_port, 
      positive_inputs_30_26_port, positive_inputs_30_25_port, 
      positive_inputs_30_24_port, positive_inputs_30_23_port, 
      positive_inputs_30_22_port, positive_inputs_30_21_port, 
      positive_inputs_30_20_port, positive_inputs_30_19_port, 
      positive_inputs_30_18_port, positive_inputs_30_17_port, 
      positive_inputs_30_16_port, positive_inputs_30_15_port, 
      positive_inputs_30_14_port, positive_inputs_30_13_port, 
      positive_inputs_30_12_port, positive_inputs_30_11_port, 
      positive_inputs_30_10_port, positive_inputs_30_9_port, 
      positive_inputs_30_8_port, positive_inputs_30_7_port, 
      positive_inputs_30_6_port, positive_inputs_30_5_port, 
      positive_inputs_30_4_port, positive_inputs_30_3_port, 
      positive_inputs_30_2_port, positive_inputs_30_1_port, 
      positive_inputs_29_63_port, positive_inputs_29_62_port, 
      positive_inputs_29_61_port, positive_inputs_29_60_port, 
      positive_inputs_29_59_port, positive_inputs_29_58_port, 
      positive_inputs_29_57_port, positive_inputs_29_56_port, 
      positive_inputs_29_55_port, positive_inputs_29_54_port, 
      positive_inputs_29_53_port, positive_inputs_29_52_port, 
      positive_inputs_29_51_port, positive_inputs_29_50_port, 
      positive_inputs_29_49_port, positive_inputs_29_48_port, 
      positive_inputs_29_47_port, positive_inputs_29_46_port, 
      positive_inputs_29_45_port, positive_inputs_29_44_port, 
      positive_inputs_29_43_port, positive_inputs_29_42_port, 
      positive_inputs_29_41_port, positive_inputs_29_40_port, 
      positive_inputs_29_39_port, positive_inputs_29_38_port, 
      positive_inputs_29_37_port, positive_inputs_29_36_port, 
      positive_inputs_29_35_port, positive_inputs_29_34_port, 
      positive_inputs_29_33_port, positive_inputs_29_32_port, 
      positive_inputs_29_31_port, positive_inputs_29_30_port, 
      positive_inputs_29_29_port, positive_inputs_29_28_port, 
      positive_inputs_29_27_port, positive_inputs_29_26_port, 
      positive_inputs_29_25_port, positive_inputs_29_24_port, 
      positive_inputs_29_23_port, positive_inputs_29_22_port, 
      positive_inputs_29_21_port, positive_inputs_29_20_port, 
      positive_inputs_29_19_port, positive_inputs_29_18_port, 
      positive_inputs_29_17_port, positive_inputs_29_16_port, 
      positive_inputs_29_15_port, positive_inputs_29_14_port, 
      positive_inputs_29_13_port, positive_inputs_29_12_port, 
      positive_inputs_29_11_port, positive_inputs_29_10_port, 
      positive_inputs_29_9_port, positive_inputs_29_8_port, 
      positive_inputs_29_7_port, positive_inputs_29_6_port, 
      positive_inputs_29_5_port, positive_inputs_29_4_port, 
      positive_inputs_29_3_port, positive_inputs_29_2_port, 
      positive_inputs_29_1_port, positive_inputs_28_63_port, 
      positive_inputs_28_62_port, positive_inputs_28_61_port, 
      positive_inputs_28_60_port, positive_inputs_28_59_port, 
      positive_inputs_28_58_port, positive_inputs_28_57_port, 
      positive_inputs_28_56_port, positive_inputs_28_55_port, 
      positive_inputs_28_54_port, positive_inputs_28_53_port, 
      positive_inputs_28_52_port, positive_inputs_28_51_port, 
      positive_inputs_28_50_port, positive_inputs_28_49_port, 
      positive_inputs_28_48_port, positive_inputs_28_47_port, 
      positive_inputs_28_46_port, positive_inputs_28_45_port, 
      positive_inputs_28_44_port, positive_inputs_28_43_port, 
      positive_inputs_28_42_port, positive_inputs_28_41_port, 
      positive_inputs_28_40_port, positive_inputs_28_39_port, 
      positive_inputs_28_38_port, positive_inputs_28_37_port, 
      positive_inputs_28_36_port, positive_inputs_28_35_port, 
      positive_inputs_28_34_port, positive_inputs_28_33_port, 
      positive_inputs_28_32_port, positive_inputs_28_31_port, 
      positive_inputs_28_30_port, positive_inputs_28_29_port, 
      positive_inputs_28_28_port, positive_inputs_28_27_port, 
      positive_inputs_28_26_port, positive_inputs_28_25_port, 
      positive_inputs_28_24_port, positive_inputs_28_23_port, 
      positive_inputs_28_22_port, positive_inputs_28_21_port, 
      positive_inputs_28_20_port, positive_inputs_28_19_port, 
      positive_inputs_28_18_port, positive_inputs_28_17_port, 
      positive_inputs_28_16_port, positive_inputs_28_15_port, 
      positive_inputs_28_14_port, positive_inputs_28_13_port, 
      positive_inputs_28_12_port, positive_inputs_28_11_port, 
      positive_inputs_28_10_port, positive_inputs_28_9_port, 
      positive_inputs_28_8_port, positive_inputs_28_7_port, 
      positive_inputs_28_6_port, positive_inputs_28_5_port, 
      positive_inputs_28_4_port, positive_inputs_28_3_port, 
      positive_inputs_28_2_port, positive_inputs_28_1_port, 
      positive_inputs_27_63_port, positive_inputs_27_62_port, 
      positive_inputs_27_61_port, positive_inputs_27_60_port, 
      positive_inputs_27_59_port, positive_inputs_27_58_port, 
      positive_inputs_27_57_port, positive_inputs_27_56_port, 
      positive_inputs_27_55_port, positive_inputs_27_54_port, 
      positive_inputs_27_53_port, positive_inputs_27_52_port, 
      positive_inputs_27_51_port, positive_inputs_27_50_port, 
      positive_inputs_27_49_port, positive_inputs_27_48_port, 
      positive_inputs_27_47_port, positive_inputs_27_46_port, 
      positive_inputs_27_45_port, positive_inputs_27_44_port, 
      positive_inputs_27_43_port, positive_inputs_27_42_port, 
      positive_inputs_27_41_port, positive_inputs_27_40_port, 
      positive_inputs_27_39_port, positive_inputs_27_38_port, 
      positive_inputs_27_37_port, positive_inputs_27_36_port, 
      positive_inputs_27_35_port, positive_inputs_27_34_port, 
      positive_inputs_27_33_port, positive_inputs_27_32_port, 
      positive_inputs_27_31_port, positive_inputs_27_30_port, 
      positive_inputs_27_29_port, positive_inputs_27_28_port, 
      positive_inputs_27_27_port, positive_inputs_27_26_port, 
      positive_inputs_27_25_port, positive_inputs_27_24_port, 
      positive_inputs_27_23_port, positive_inputs_27_22_port, 
      positive_inputs_27_21_port, positive_inputs_27_20_port, 
      positive_inputs_27_19_port, positive_inputs_27_18_port, 
      positive_inputs_27_17_port, positive_inputs_27_16_port, 
      positive_inputs_27_15_port, positive_inputs_27_14_port, 
      positive_inputs_27_13_port, positive_inputs_27_12_port, 
      positive_inputs_27_11_port, positive_inputs_27_10_port, 
      positive_inputs_27_9_port, positive_inputs_27_8_port, 
      positive_inputs_27_7_port, positive_inputs_27_6_port, 
      positive_inputs_27_5_port, positive_inputs_27_4_port, 
      positive_inputs_27_3_port, positive_inputs_27_2_port, 
      positive_inputs_27_1_port, positive_inputs_26_63_port, 
      positive_inputs_26_62_port, positive_inputs_26_61_port, 
      positive_inputs_26_60_port, positive_inputs_26_59_port, 
      positive_inputs_26_58_port, positive_inputs_26_57_port, 
      positive_inputs_26_56_port, positive_inputs_26_55_port, 
      positive_inputs_26_54_port, positive_inputs_26_53_port, 
      positive_inputs_26_52_port, positive_inputs_26_51_port, 
      positive_inputs_26_50_port, positive_inputs_26_49_port, 
      positive_inputs_26_48_port, positive_inputs_26_47_port, 
      positive_inputs_26_46_port, positive_inputs_26_45_port, 
      positive_inputs_26_44_port, positive_inputs_26_43_port, 
      positive_inputs_26_42_port, positive_inputs_26_41_port, 
      positive_inputs_26_40_port, positive_inputs_26_39_port, 
      positive_inputs_26_38_port, positive_inputs_26_37_port, 
      positive_inputs_26_36_port, positive_inputs_26_35_port, 
      positive_inputs_26_34_port, positive_inputs_26_33_port, 
      positive_inputs_26_32_port, positive_inputs_26_31_port, 
      positive_inputs_26_30_port, positive_inputs_26_29_port, 
      positive_inputs_26_28_port, positive_inputs_26_27_port, 
      positive_inputs_26_26_port, positive_inputs_26_25_port, 
      positive_inputs_26_24_port, positive_inputs_26_23_port, 
      positive_inputs_26_22_port, positive_inputs_26_21_port, 
      positive_inputs_26_20_port, positive_inputs_26_19_port, 
      positive_inputs_26_18_port, positive_inputs_26_17_port, 
      positive_inputs_26_16_port, positive_inputs_26_15_port, 
      positive_inputs_26_14_port, positive_inputs_26_13_port, 
      positive_inputs_26_12_port, positive_inputs_26_11_port, 
      positive_inputs_26_10_port, positive_inputs_26_9_port, 
      positive_inputs_26_8_port, positive_inputs_26_7_port, 
      positive_inputs_26_6_port, positive_inputs_26_5_port, 
      positive_inputs_26_4_port, positive_inputs_26_3_port, 
      positive_inputs_26_2_port, positive_inputs_26_1_port, 
      positive_inputs_25_63_port, positive_inputs_25_62_port, 
      positive_inputs_25_61_port, positive_inputs_25_60_port, 
      positive_inputs_25_59_port, positive_inputs_25_58_port, 
      positive_inputs_25_57_port, positive_inputs_25_56_port, 
      positive_inputs_25_55_port, positive_inputs_25_54_port, 
      positive_inputs_25_53_port, positive_inputs_25_52_port, 
      positive_inputs_25_51_port, positive_inputs_25_50_port, 
      positive_inputs_25_49_port, positive_inputs_25_48_port, 
      positive_inputs_25_47_port, positive_inputs_25_46_port, 
      positive_inputs_25_45_port, positive_inputs_25_44_port, 
      positive_inputs_25_43_port, positive_inputs_25_42_port, 
      positive_inputs_25_41_port, positive_inputs_25_40_port, 
      positive_inputs_25_39_port, positive_inputs_25_38_port, 
      positive_inputs_25_37_port, positive_inputs_25_36_port, 
      positive_inputs_25_35_port, positive_inputs_25_34_port, 
      positive_inputs_25_33_port, positive_inputs_25_32_port, 
      positive_inputs_25_31_port, positive_inputs_25_30_port, 
      positive_inputs_25_29_port, positive_inputs_25_28_port, 
      positive_inputs_25_27_port, positive_inputs_25_26_port, 
      positive_inputs_25_25_port, positive_inputs_25_24_port, 
      positive_inputs_25_23_port, positive_inputs_25_22_port, 
      positive_inputs_25_21_port, positive_inputs_25_20_port, 
      positive_inputs_25_19_port, positive_inputs_25_18_port, 
      positive_inputs_25_17_port, positive_inputs_25_16_port, 
      positive_inputs_25_15_port, positive_inputs_25_14_port, 
      positive_inputs_25_13_port, positive_inputs_25_12_port, 
      positive_inputs_25_11_port, positive_inputs_25_10_port, 
      positive_inputs_25_9_port, positive_inputs_25_8_port, 
      positive_inputs_25_7_port, positive_inputs_25_6_port, 
      positive_inputs_25_5_port, positive_inputs_25_4_port, 
      positive_inputs_25_3_port, positive_inputs_25_2_port, 
      positive_inputs_25_1_port, negative_inputs_8_63_port, 
      negative_inputs_8_62_port, negative_inputs_8_61_port, 
      negative_inputs_8_60_port, negative_inputs_8_59_port, 
      negative_inputs_8_58_port, negative_inputs_8_57_port, 
      negative_inputs_8_56_port, negative_inputs_8_55_port, 
      negative_inputs_8_54_port, negative_inputs_8_53_port, 
      negative_inputs_8_52_port, negative_inputs_8_51_port, 
      negative_inputs_8_50_port, negative_inputs_8_49_port, 
      negative_inputs_8_48_port, negative_inputs_8_47_port, 
      negative_inputs_8_46_port, negative_inputs_8_45_port, 
      negative_inputs_8_44_port, negative_inputs_8_43_port, 
      negative_inputs_8_42_port, negative_inputs_8_41_port, 
      negative_inputs_8_40_port, negative_inputs_8_39_port, 
      negative_inputs_8_38_port, negative_inputs_8_37_port, 
      negative_inputs_8_36_port, negative_inputs_8_35_port, 
      negative_inputs_8_34_port, negative_inputs_8_33_port, 
      negative_inputs_8_32_port, negative_inputs_8_31_port, 
      negative_inputs_8_30_port, negative_inputs_8_29_port, 
      negative_inputs_8_28_port, negative_inputs_8_27_port, 
      negative_inputs_8_26_port, negative_inputs_8_25_port, 
      negative_inputs_8_24_port, negative_inputs_8_23_port, 
      negative_inputs_8_22_port, negative_inputs_8_21_port, 
      negative_inputs_8_20_port, negative_inputs_8_19_port, 
      negative_inputs_8_18_port, negative_inputs_8_17_port, 
      negative_inputs_8_16_port, negative_inputs_8_15_port, 
      negative_inputs_8_14_port, negative_inputs_8_13_port, 
      negative_inputs_8_12_port, negative_inputs_8_11_port, 
      negative_inputs_8_10_port, negative_inputs_8_9_port, 
      negative_inputs_8_8_port, negative_inputs_8_7_port, 
      negative_inputs_8_6_port, negative_inputs_8_5_port, 
      negative_inputs_8_4_port, negative_inputs_8_3_port, 
      negative_inputs_8_2_port, negative_inputs_8_1_port, 
      negative_inputs_7_63_port, negative_inputs_7_62_port, 
      negative_inputs_7_61_port, negative_inputs_7_60_port, 
      negative_inputs_7_59_port, negative_inputs_7_58_port, 
      negative_inputs_7_57_port, negative_inputs_7_56_port, 
      negative_inputs_7_55_port, negative_inputs_7_54_port, 
      negative_inputs_7_53_port, negative_inputs_7_52_port, 
      negative_inputs_7_51_port, negative_inputs_7_50_port, 
      negative_inputs_7_49_port, negative_inputs_7_48_port, 
      negative_inputs_7_47_port, negative_inputs_7_46_port, 
      negative_inputs_7_45_port, negative_inputs_7_44_port, 
      negative_inputs_7_43_port, negative_inputs_7_42_port, 
      negative_inputs_7_41_port, negative_inputs_7_40_port, 
      negative_inputs_7_39_port, negative_inputs_7_38_port, 
      negative_inputs_7_37_port, negative_inputs_7_36_port, 
      negative_inputs_7_35_port, negative_inputs_7_34_port, 
      negative_inputs_7_33_port, negative_inputs_7_32_port, 
      negative_inputs_7_31_port, negative_inputs_7_30_port, 
      negative_inputs_7_29_port, negative_inputs_7_28_port, 
      negative_inputs_7_27_port, negative_inputs_7_26_port, 
      negative_inputs_7_25_port, negative_inputs_7_24_port, 
      negative_inputs_7_23_port, negative_inputs_7_22_port, 
      negative_inputs_7_21_port, negative_inputs_7_20_port, 
      negative_inputs_7_19_port, negative_inputs_7_18_port, 
      negative_inputs_7_17_port, negative_inputs_7_16_port, 
      negative_inputs_7_15_port, negative_inputs_7_14_port, 
      negative_inputs_7_13_port, negative_inputs_7_12_port, 
      negative_inputs_7_11_port, negative_inputs_7_10_port, 
      negative_inputs_7_9_port, negative_inputs_7_8_port, 
      negative_inputs_7_7_port, negative_inputs_7_6_port, 
      negative_inputs_7_5_port, negative_inputs_7_4_port, 
      negative_inputs_7_3_port, negative_inputs_7_2_port, 
      negative_inputs_7_1_port, negative_inputs_6_63_port, 
      negative_inputs_6_62_port, negative_inputs_6_61_port, 
      negative_inputs_6_60_port, negative_inputs_6_59_port, 
      negative_inputs_6_58_port, negative_inputs_6_57_port, 
      negative_inputs_6_56_port, negative_inputs_6_55_port, 
      negative_inputs_6_54_port, negative_inputs_6_53_port, 
      negative_inputs_6_52_port, negative_inputs_6_51_port, 
      negative_inputs_6_50_port, negative_inputs_6_49_port, 
      negative_inputs_6_48_port, negative_inputs_6_47_port, 
      negative_inputs_6_46_port, negative_inputs_6_45_port, 
      negative_inputs_6_44_port, negative_inputs_6_43_port, 
      negative_inputs_6_42_port, negative_inputs_6_41_port, 
      negative_inputs_6_40_port, negative_inputs_6_39_port, 
      negative_inputs_6_38_port, negative_inputs_6_37_port, 
      negative_inputs_6_36_port, negative_inputs_6_35_port, 
      negative_inputs_6_34_port, negative_inputs_6_33_port, 
      negative_inputs_6_32_port, negative_inputs_6_31_port, 
      negative_inputs_6_30_port, negative_inputs_6_29_port, 
      negative_inputs_6_28_port, negative_inputs_6_27_port, 
      negative_inputs_6_26_port, negative_inputs_6_25_port, 
      negative_inputs_6_24_port, negative_inputs_6_23_port, 
      negative_inputs_6_22_port, negative_inputs_6_21_port, 
      negative_inputs_6_20_port, negative_inputs_6_19_port, 
      negative_inputs_6_18_port, negative_inputs_6_17_port, 
      negative_inputs_6_16_port, negative_inputs_6_15_port, 
      negative_inputs_6_14_port, negative_inputs_6_13_port, 
      negative_inputs_6_12_port, negative_inputs_6_11_port, 
      negative_inputs_6_10_port, negative_inputs_6_9_port, 
      negative_inputs_6_8_port, negative_inputs_6_7_port, 
      negative_inputs_6_6_port, negative_inputs_6_5_port, 
      negative_inputs_6_4_port, negative_inputs_6_3_port, 
      negative_inputs_6_2_port, negative_inputs_6_1_port, 
      negative_inputs_5_63_port, negative_inputs_5_62_port, 
      negative_inputs_5_61_port, negative_inputs_5_60_port, 
      negative_inputs_5_59_port, negative_inputs_5_58_port, 
      negative_inputs_5_57_port, negative_inputs_5_56_port, 
      negative_inputs_5_55_port, negative_inputs_5_54_port, 
      negative_inputs_5_53_port, negative_inputs_5_52_port, 
      negative_inputs_5_51_port, negative_inputs_5_50_port, 
      negative_inputs_5_49_port, negative_inputs_5_48_port, 
      negative_inputs_5_47_port, negative_inputs_5_46_port, 
      negative_inputs_5_45_port, negative_inputs_5_44_port, 
      negative_inputs_5_43_port, negative_inputs_5_42_port, 
      negative_inputs_5_41_port, negative_inputs_5_40_port, 
      negative_inputs_5_39_port, negative_inputs_5_38_port, 
      negative_inputs_5_37_port, negative_inputs_5_36_port, 
      negative_inputs_5_35_port, negative_inputs_5_34_port, 
      negative_inputs_5_33_port, negative_inputs_5_32_port, 
      negative_inputs_5_31_port, negative_inputs_5_30_port, 
      negative_inputs_5_29_port, negative_inputs_5_28_port, 
      negative_inputs_5_27_port, negative_inputs_5_26_port, 
      negative_inputs_5_25_port, negative_inputs_5_24_port, 
      negative_inputs_5_23_port, negative_inputs_5_22_port, 
      negative_inputs_5_21_port, negative_inputs_5_20_port, 
      negative_inputs_5_19_port, negative_inputs_5_18_port, 
      negative_inputs_5_17_port, negative_inputs_5_16_port, 
      negative_inputs_5_15_port, negative_inputs_5_14_port, 
      negative_inputs_5_13_port, negative_inputs_5_12_port, 
      negative_inputs_5_11_port, negative_inputs_5_10_port, 
      negative_inputs_5_9_port, negative_inputs_5_8_port, 
      negative_inputs_5_7_port, negative_inputs_5_6_port, 
      negative_inputs_5_5_port, negative_inputs_5_4_port, 
      negative_inputs_5_3_port, negative_inputs_5_2_port, 
      negative_inputs_5_1_port, negative_inputs_4_63_port, 
      negative_inputs_4_62_port, negative_inputs_4_61_port, 
      negative_inputs_4_60_port, negative_inputs_4_59_port, 
      negative_inputs_4_58_port, negative_inputs_4_57_port, 
      negative_inputs_4_56_port, negative_inputs_4_55_port, 
      negative_inputs_4_54_port, negative_inputs_4_53_port, 
      negative_inputs_4_52_port, negative_inputs_4_51_port, 
      negative_inputs_4_50_port, negative_inputs_4_49_port, 
      negative_inputs_4_48_port, negative_inputs_4_47_port, 
      negative_inputs_4_46_port, negative_inputs_4_45_port, 
      negative_inputs_4_44_port, negative_inputs_4_43_port, 
      negative_inputs_4_42_port, negative_inputs_4_41_port, 
      negative_inputs_4_40_port, negative_inputs_4_39_port, 
      negative_inputs_4_38_port, negative_inputs_4_37_port, 
      negative_inputs_4_36_port, negative_inputs_4_35_port, 
      negative_inputs_4_34_port, negative_inputs_4_33_port, 
      negative_inputs_4_32_port, negative_inputs_4_31_port, 
      negative_inputs_4_30_port, negative_inputs_4_29_port, 
      negative_inputs_4_28_port, negative_inputs_4_27_port, 
      negative_inputs_4_26_port, negative_inputs_4_25_port, 
      negative_inputs_4_24_port, negative_inputs_4_23_port, 
      negative_inputs_4_22_port, negative_inputs_4_21_port, 
      negative_inputs_4_20_port, negative_inputs_4_19_port, 
      negative_inputs_4_18_port, negative_inputs_4_17_port, 
      negative_inputs_4_16_port, negative_inputs_4_15_port, 
      negative_inputs_4_14_port, negative_inputs_4_13_port, 
      negative_inputs_4_12_port, negative_inputs_4_11_port, 
      negative_inputs_4_10_port, negative_inputs_4_9_port, 
      negative_inputs_4_8_port, negative_inputs_4_7_port, 
      negative_inputs_4_6_port, negative_inputs_4_5_port, 
      negative_inputs_4_4_port, negative_inputs_4_3_port, 
      negative_inputs_4_2_port, negative_inputs_4_1_port, 
      negative_inputs_3_63_port, negative_inputs_3_62_port, 
      negative_inputs_3_61_port, negative_inputs_3_60_port, 
      negative_inputs_3_59_port, negative_inputs_3_58_port, 
      negative_inputs_3_57_port, negative_inputs_3_56_port, 
      negative_inputs_3_55_port, negative_inputs_3_54_port, 
      negative_inputs_3_53_port, negative_inputs_3_52_port, 
      negative_inputs_3_51_port, negative_inputs_3_50_port, 
      negative_inputs_3_49_port, negative_inputs_3_48_port, 
      negative_inputs_3_47_port, negative_inputs_3_46_port, 
      negative_inputs_3_45_port, negative_inputs_3_44_port, 
      negative_inputs_3_43_port, negative_inputs_3_42_port, 
      negative_inputs_3_41_port, negative_inputs_3_40_port, 
      negative_inputs_3_39_port, negative_inputs_3_38_port, 
      negative_inputs_3_37_port, negative_inputs_3_36_port, 
      negative_inputs_3_35_port, negative_inputs_3_34_port, 
      negative_inputs_3_33_port, negative_inputs_3_32_port, 
      negative_inputs_3_31_port, negative_inputs_3_30_port, 
      negative_inputs_3_29_port, negative_inputs_3_28_port, 
      negative_inputs_3_27_port, negative_inputs_3_26_port, 
      negative_inputs_3_25_port, negative_inputs_3_24_port, 
      negative_inputs_3_23_port, negative_inputs_3_22_port, 
      negative_inputs_3_21_port, negative_inputs_3_20_port, 
      negative_inputs_3_19_port, negative_inputs_3_18_port, 
      negative_inputs_3_17_port, negative_inputs_3_16_port, 
      negative_inputs_3_15_port, negative_inputs_3_14_port, 
      negative_inputs_3_13_port, negative_inputs_3_12_port, 
      negative_inputs_3_11_port, negative_inputs_3_10_port, 
      negative_inputs_3_9_port, negative_inputs_3_8_port, 
      negative_inputs_3_7_port, negative_inputs_3_6_port, 
      negative_inputs_3_5_port, negative_inputs_3_4_port, 
      negative_inputs_3_3_port, negative_inputs_3_2_port, 
      negative_inputs_3_1_port, negative_inputs_2_63_port, 
      negative_inputs_2_62_port, negative_inputs_2_61_port, 
      negative_inputs_2_60_port, negative_inputs_2_59_port, 
      negative_inputs_2_58_port, negative_inputs_2_57_port, 
      negative_inputs_2_56_port, negative_inputs_2_55_port, 
      negative_inputs_2_54_port, negative_inputs_2_53_port, 
      negative_inputs_2_52_port, negative_inputs_2_51_port, 
      negative_inputs_2_50_port, negative_inputs_2_49_port, 
      negative_inputs_2_48_port, negative_inputs_2_47_port, 
      negative_inputs_2_46_port, negative_inputs_2_45_port, 
      negative_inputs_2_44_port, negative_inputs_2_43_port, 
      negative_inputs_2_42_port, negative_inputs_2_41_port, 
      negative_inputs_2_40_port, negative_inputs_2_39_port, 
      negative_inputs_2_38_port, negative_inputs_2_37_port, 
      negative_inputs_2_36_port, negative_inputs_2_35_port, 
      negative_inputs_2_34_port, negative_inputs_2_33_port, 
      negative_inputs_2_32_port, negative_inputs_2_31_port, 
      negative_inputs_2_30_port, negative_inputs_2_29_port, 
      negative_inputs_2_28_port, negative_inputs_2_27_port, 
      negative_inputs_2_26_port, negative_inputs_2_25_port, 
      negative_inputs_2_24_port, negative_inputs_2_23_port, 
      negative_inputs_2_22_port, negative_inputs_2_21_port, 
      negative_inputs_2_20_port, negative_inputs_2_19_port, 
      negative_inputs_2_18_port, negative_inputs_2_17_port, 
      negative_inputs_2_16_port, negative_inputs_2_15_port, 
      negative_inputs_2_14_port, negative_inputs_2_13_port, 
      negative_inputs_2_12_port, negative_inputs_2_11_port, 
      negative_inputs_2_10_port, negative_inputs_2_9_port, 
      negative_inputs_2_8_port, negative_inputs_2_7_port, 
      negative_inputs_2_6_port, negative_inputs_2_5_port, 
      negative_inputs_2_4_port, negative_inputs_2_3_port, 
      negative_inputs_2_2_port, negative_inputs_2_1_port, 
      negative_inputs_1_63_port, negative_inputs_1_62_port, 
      negative_inputs_1_61_port, negative_inputs_1_60_port, 
      negative_inputs_1_59_port, negative_inputs_1_58_port, 
      negative_inputs_1_57_port, negative_inputs_1_56_port, 
      negative_inputs_1_55_port, negative_inputs_1_54_port, 
      negative_inputs_1_53_port, negative_inputs_1_52_port, 
      negative_inputs_1_51_port, negative_inputs_1_50_port, 
      negative_inputs_1_49_port, negative_inputs_1_48_port, 
      negative_inputs_1_47_port, negative_inputs_1_46_port, 
      negative_inputs_1_45_port, negative_inputs_1_44_port, 
      negative_inputs_1_43_port, negative_inputs_1_42_port, 
      negative_inputs_1_41_port, negative_inputs_1_40_port, 
      negative_inputs_1_39_port, negative_inputs_1_38_port, 
      negative_inputs_1_37_port, negative_inputs_1_36_port, 
      negative_inputs_1_35_port, negative_inputs_1_34_port, 
      negative_inputs_1_33_port, negative_inputs_1_32_port, 
      negative_inputs_1_31_port, negative_inputs_1_30_port, 
      negative_inputs_1_29_port, negative_inputs_1_28_port, 
      negative_inputs_1_27_port, negative_inputs_1_26_port, 
      negative_inputs_1_25_port, negative_inputs_1_24_port, 
      negative_inputs_1_23_port, negative_inputs_1_22_port, 
      negative_inputs_1_21_port, negative_inputs_1_20_port, 
      negative_inputs_1_19_port, negative_inputs_1_18_port, 
      negative_inputs_1_17_port, negative_inputs_1_16_port, 
      negative_inputs_1_15_port, negative_inputs_1_14_port, 
      negative_inputs_1_13_port, negative_inputs_1_12_port, 
      negative_inputs_1_11_port, negative_inputs_1_10_port, 
      negative_inputs_1_9_port, negative_inputs_1_8_port, 
      negative_inputs_1_7_port, negative_inputs_1_6_port, 
      negative_inputs_1_5_port, negative_inputs_1_4_port, 
      negative_inputs_1_3_port, negative_inputs_1_2_port, 
      negative_inputs_1_1_port, negative_inputs_16_63_port, 
      negative_inputs_16_62_port, negative_inputs_16_61_port, 
      negative_inputs_16_60_port, negative_inputs_16_59_port, 
      negative_inputs_16_58_port, negative_inputs_16_57_port, 
      negative_inputs_16_56_port, negative_inputs_16_55_port, 
      negative_inputs_16_54_port, negative_inputs_16_53_port, 
      negative_inputs_16_52_port, negative_inputs_16_51_port, 
      negative_inputs_16_50_port, negative_inputs_16_49_port, 
      negative_inputs_16_48_port, negative_inputs_16_47_port, 
      negative_inputs_16_46_port, negative_inputs_16_45_port, 
      negative_inputs_16_44_port, negative_inputs_16_43_port, 
      negative_inputs_16_42_port, negative_inputs_16_41_port, 
      negative_inputs_16_40_port, negative_inputs_16_39_port, 
      negative_inputs_16_38_port, negative_inputs_16_37_port, 
      negative_inputs_16_36_port, negative_inputs_16_35_port, 
      negative_inputs_16_34_port, negative_inputs_16_33_port, 
      negative_inputs_16_32_port, negative_inputs_16_31_port, 
      negative_inputs_16_30_port, negative_inputs_16_29_port, 
      negative_inputs_16_28_port, negative_inputs_16_27_port, 
      negative_inputs_16_26_port, negative_inputs_16_25_port, 
      negative_inputs_16_24_port, negative_inputs_16_23_port, 
      negative_inputs_16_22_port, negative_inputs_16_21_port, 
      negative_inputs_16_20_port, negative_inputs_16_19_port, 
      negative_inputs_16_18_port, negative_inputs_16_17_port, 
      negative_inputs_16_16_port, negative_inputs_16_15_port, 
      negative_inputs_16_14_port, negative_inputs_16_13_port, 
      negative_inputs_16_12_port, negative_inputs_16_11_port, 
      negative_inputs_16_10_port, negative_inputs_16_9_port, 
      negative_inputs_16_8_port, negative_inputs_16_7_port, 
      negative_inputs_16_6_port, negative_inputs_16_5_port, 
      negative_inputs_16_4_port, negative_inputs_16_3_port, 
      negative_inputs_16_2_port, negative_inputs_16_1_port, 
      negative_inputs_15_63_port, negative_inputs_15_62_port, 
      negative_inputs_15_61_port, negative_inputs_15_60_port, 
      negative_inputs_15_59_port, negative_inputs_15_58_port, 
      negative_inputs_15_57_port, negative_inputs_15_56_port, 
      negative_inputs_15_55_port, negative_inputs_15_54_port, 
      negative_inputs_15_53_port, negative_inputs_15_52_port, 
      negative_inputs_15_51_port, negative_inputs_15_50_port, 
      negative_inputs_15_49_port, negative_inputs_15_48_port, 
      negative_inputs_15_47_port, negative_inputs_15_46_port, 
      negative_inputs_15_45_port, negative_inputs_15_44_port, 
      negative_inputs_15_43_port, negative_inputs_15_42_port, 
      negative_inputs_15_41_port, negative_inputs_15_40_port, 
      negative_inputs_15_39_port, negative_inputs_15_38_port, 
      negative_inputs_15_37_port, negative_inputs_15_36_port, 
      negative_inputs_15_35_port, negative_inputs_15_34_port, 
      negative_inputs_15_33_port, negative_inputs_15_32_port, 
      negative_inputs_15_31_port, negative_inputs_15_30_port, 
      negative_inputs_15_29_port, negative_inputs_15_28_port, 
      negative_inputs_15_27_port, negative_inputs_15_26_port, 
      negative_inputs_15_25_port, negative_inputs_15_24_port, 
      negative_inputs_15_23_port, negative_inputs_15_22_port, 
      negative_inputs_15_21_port, negative_inputs_15_20_port, 
      negative_inputs_15_19_port, negative_inputs_15_18_port, 
      negative_inputs_15_17_port, negative_inputs_15_16_port, 
      negative_inputs_15_15_port, negative_inputs_15_14_port, 
      negative_inputs_15_13_port, negative_inputs_15_12_port, 
      negative_inputs_15_11_port, negative_inputs_15_10_port, 
      negative_inputs_15_9_port, negative_inputs_15_8_port, 
      negative_inputs_15_7_port, negative_inputs_15_6_port, 
      negative_inputs_15_5_port, negative_inputs_15_4_port, 
      negative_inputs_15_3_port, negative_inputs_15_2_port, 
      negative_inputs_15_1_port, negative_inputs_14_63_port, 
      negative_inputs_14_62_port, negative_inputs_14_61_port, 
      negative_inputs_14_60_port, negative_inputs_14_59_port, 
      negative_inputs_14_58_port, negative_inputs_14_57_port, 
      negative_inputs_14_56_port, negative_inputs_14_55_port, 
      negative_inputs_14_54_port, negative_inputs_14_53_port, 
      negative_inputs_14_52_port, negative_inputs_14_51_port, 
      negative_inputs_14_50_port, negative_inputs_14_49_port, 
      negative_inputs_14_48_port, negative_inputs_14_47_port, 
      negative_inputs_14_46_port, negative_inputs_14_45_port, 
      negative_inputs_14_44_port, negative_inputs_14_43_port, 
      negative_inputs_14_42_port, negative_inputs_14_41_port, 
      negative_inputs_14_40_port, negative_inputs_14_39_port, 
      negative_inputs_14_38_port, negative_inputs_14_37_port, 
      negative_inputs_14_36_port, negative_inputs_14_35_port, 
      negative_inputs_14_34_port, negative_inputs_14_33_port, 
      negative_inputs_14_32_port, negative_inputs_14_31_port, 
      negative_inputs_14_30_port, negative_inputs_14_29_port, 
      negative_inputs_14_28_port, negative_inputs_14_27_port, 
      negative_inputs_14_26_port, negative_inputs_14_25_port, 
      negative_inputs_14_24_port, negative_inputs_14_23_port, 
      negative_inputs_14_22_port, negative_inputs_14_21_port, 
      negative_inputs_14_20_port, negative_inputs_14_19_port, 
      negative_inputs_14_18_port, negative_inputs_14_17_port, 
      negative_inputs_14_16_port, negative_inputs_14_15_port, 
      negative_inputs_14_14_port, negative_inputs_14_13_port, 
      negative_inputs_14_12_port, negative_inputs_14_11_port, 
      negative_inputs_14_10_port, negative_inputs_14_9_port, 
      negative_inputs_14_8_port, negative_inputs_14_7_port, 
      negative_inputs_14_6_port, negative_inputs_14_5_port, 
      negative_inputs_14_4_port, negative_inputs_14_3_port, 
      negative_inputs_14_2_port, negative_inputs_14_1_port, 
      negative_inputs_13_63_port, negative_inputs_13_62_port, 
      negative_inputs_13_61_port, negative_inputs_13_60_port, 
      negative_inputs_13_59_port, negative_inputs_13_58_port, 
      negative_inputs_13_57_port, negative_inputs_13_56_port, 
      negative_inputs_13_55_port, negative_inputs_13_54_port, 
      negative_inputs_13_53_port, negative_inputs_13_52_port, 
      negative_inputs_13_51_port, negative_inputs_13_50_port, 
      negative_inputs_13_49_port, negative_inputs_13_48_port, 
      negative_inputs_13_47_port, negative_inputs_13_46_port, 
      negative_inputs_13_45_port, negative_inputs_13_44_port, 
      negative_inputs_13_43_port, negative_inputs_13_42_port, 
      negative_inputs_13_41_port, negative_inputs_13_40_port, 
      negative_inputs_13_39_port, negative_inputs_13_38_port, 
      negative_inputs_13_37_port, negative_inputs_13_36_port, 
      negative_inputs_13_35_port, negative_inputs_13_34_port, 
      negative_inputs_13_33_port, negative_inputs_13_32_port, 
      negative_inputs_13_31_port, negative_inputs_13_30_port, 
      negative_inputs_13_29_port, negative_inputs_13_28_port, 
      negative_inputs_13_27_port, negative_inputs_13_26_port, 
      negative_inputs_13_25_port, negative_inputs_13_24_port, 
      negative_inputs_13_23_port, negative_inputs_13_22_port, 
      negative_inputs_13_21_port, negative_inputs_13_20_port, 
      negative_inputs_13_19_port, negative_inputs_13_18_port, 
      negative_inputs_13_17_port, negative_inputs_13_16_port, 
      negative_inputs_13_15_port, negative_inputs_13_14_port, 
      negative_inputs_13_13_port, negative_inputs_13_12_port, 
      negative_inputs_13_11_port, negative_inputs_13_10_port, 
      negative_inputs_13_9_port, negative_inputs_13_8_port, 
      negative_inputs_13_7_port, negative_inputs_13_6_port, 
      negative_inputs_13_5_port, negative_inputs_13_4_port, 
      negative_inputs_13_3_port, negative_inputs_13_2_port, 
      negative_inputs_13_1_port, negative_inputs_12_63_port, 
      negative_inputs_12_62_port, negative_inputs_12_61_port, 
      negative_inputs_12_60_port, negative_inputs_12_59_port, 
      negative_inputs_12_58_port, negative_inputs_12_57_port, 
      negative_inputs_12_56_port, negative_inputs_12_55_port, 
      negative_inputs_12_54_port, negative_inputs_12_53_port, 
      negative_inputs_12_52_port, negative_inputs_12_51_port, 
      negative_inputs_12_50_port, negative_inputs_12_49_port, 
      negative_inputs_12_48_port, negative_inputs_12_47_port, 
      negative_inputs_12_46_port, negative_inputs_12_45_port, 
      negative_inputs_12_44_port, negative_inputs_12_43_port, 
      negative_inputs_12_42_port, negative_inputs_12_41_port, 
      negative_inputs_12_40_port, negative_inputs_12_39_port, 
      negative_inputs_12_38_port, negative_inputs_12_37_port, 
      negative_inputs_12_36_port, negative_inputs_12_35_port, 
      negative_inputs_12_34_port, negative_inputs_12_33_port, 
      negative_inputs_12_32_port, negative_inputs_12_31_port, 
      negative_inputs_12_30_port, negative_inputs_12_29_port, 
      negative_inputs_12_28_port, negative_inputs_12_27_port, 
      negative_inputs_12_26_port, negative_inputs_12_25_port, 
      negative_inputs_12_24_port, negative_inputs_12_23_port, 
      negative_inputs_12_22_port, negative_inputs_12_21_port, 
      negative_inputs_12_20_port, negative_inputs_12_19_port, 
      negative_inputs_12_18_port, negative_inputs_12_17_port, 
      negative_inputs_12_16_port, negative_inputs_12_15_port, 
      negative_inputs_12_14_port, negative_inputs_12_13_port, 
      negative_inputs_12_12_port, negative_inputs_12_11_port, 
      negative_inputs_12_10_port, negative_inputs_12_9_port, 
      negative_inputs_12_8_port, negative_inputs_12_7_port, 
      negative_inputs_12_6_port, negative_inputs_12_5_port, 
      negative_inputs_12_4_port, negative_inputs_12_3_port, 
      negative_inputs_12_2_port, negative_inputs_12_1_port, 
      negative_inputs_11_63_port, negative_inputs_11_62_port, 
      negative_inputs_11_61_port, negative_inputs_11_60_port, 
      negative_inputs_11_59_port, negative_inputs_11_58_port, 
      negative_inputs_11_57_port, negative_inputs_11_56_port, 
      negative_inputs_11_55_port, negative_inputs_11_54_port, 
      negative_inputs_11_53_port, negative_inputs_11_52_port, 
      negative_inputs_11_51_port, negative_inputs_11_50_port, 
      negative_inputs_11_49_port, negative_inputs_11_48_port, 
      negative_inputs_11_47_port, negative_inputs_11_46_port, 
      negative_inputs_11_45_port, negative_inputs_11_44_port, 
      negative_inputs_11_43_port, negative_inputs_11_42_port, 
      negative_inputs_11_41_port, negative_inputs_11_40_port, 
      negative_inputs_11_39_port, negative_inputs_11_38_port, 
      negative_inputs_11_37_port, negative_inputs_11_36_port, 
      negative_inputs_11_35_port, negative_inputs_11_34_port, 
      negative_inputs_11_33_port, negative_inputs_11_32_port, 
      negative_inputs_11_31_port, negative_inputs_11_30_port, 
      negative_inputs_11_29_port, negative_inputs_11_28_port, 
      negative_inputs_11_27_port, negative_inputs_11_26_port, 
      negative_inputs_11_25_port, negative_inputs_11_24_port, 
      negative_inputs_11_23_port, negative_inputs_11_22_port, 
      negative_inputs_11_21_port, negative_inputs_11_20_port, 
      negative_inputs_11_19_port, negative_inputs_11_18_port, 
      negative_inputs_11_17_port, negative_inputs_11_16_port, 
      negative_inputs_11_15_port, negative_inputs_11_14_port, 
      negative_inputs_11_13_port, negative_inputs_11_12_port, 
      negative_inputs_11_11_port, negative_inputs_11_10_port, 
      negative_inputs_11_9_port, negative_inputs_11_8_port, 
      negative_inputs_11_7_port, negative_inputs_11_6_port, 
      negative_inputs_11_5_port, negative_inputs_11_4_port, 
      negative_inputs_11_3_port, negative_inputs_11_2_port, 
      negative_inputs_11_1_port, negative_inputs_10_63_port, 
      negative_inputs_10_62_port, negative_inputs_10_61_port, 
      negative_inputs_10_60_port, negative_inputs_10_59_port, 
      negative_inputs_10_58_port, negative_inputs_10_57_port, 
      negative_inputs_10_56_port, negative_inputs_10_55_port, 
      negative_inputs_10_54_port, negative_inputs_10_53_port, 
      negative_inputs_10_52_port, negative_inputs_10_51_port, 
      negative_inputs_10_50_port, negative_inputs_10_49_port, 
      negative_inputs_10_48_port, negative_inputs_10_47_port, 
      negative_inputs_10_46_port, negative_inputs_10_45_port, 
      negative_inputs_10_44_port, negative_inputs_10_43_port, 
      negative_inputs_10_42_port, negative_inputs_10_41_port, 
      negative_inputs_10_40_port, negative_inputs_10_39_port, 
      negative_inputs_10_38_port, negative_inputs_10_37_port, 
      negative_inputs_10_36_port, negative_inputs_10_35_port, 
      negative_inputs_10_34_port, negative_inputs_10_33_port, 
      negative_inputs_10_32_port, negative_inputs_10_31_port, 
      negative_inputs_10_30_port, negative_inputs_10_29_port, 
      negative_inputs_10_28_port, negative_inputs_10_27_port, 
      negative_inputs_10_26_port, negative_inputs_10_25_port, 
      negative_inputs_10_24_port, negative_inputs_10_23_port, 
      negative_inputs_10_22_port, negative_inputs_10_21_port, 
      negative_inputs_10_20_port, negative_inputs_10_19_port, 
      negative_inputs_10_18_port, negative_inputs_10_17_port, 
      negative_inputs_10_16_port, negative_inputs_10_15_port, 
      negative_inputs_10_14_port, negative_inputs_10_13_port, 
      negative_inputs_10_12_port, negative_inputs_10_11_port, 
      negative_inputs_10_10_port, negative_inputs_10_9_port, 
      negative_inputs_10_8_port, negative_inputs_10_7_port, 
      negative_inputs_10_6_port, negative_inputs_10_5_port, 
      negative_inputs_10_4_port, negative_inputs_10_3_port, 
      negative_inputs_10_2_port, negative_inputs_10_1_port, 
      negative_inputs_9_63_port, negative_inputs_9_62_port, 
      negative_inputs_9_61_port, negative_inputs_9_60_port, 
      negative_inputs_9_59_port, negative_inputs_9_58_port, 
      negative_inputs_9_57_port, negative_inputs_9_56_port, 
      negative_inputs_9_55_port, negative_inputs_9_54_port, 
      negative_inputs_9_53_port, negative_inputs_9_52_port, 
      negative_inputs_9_51_port, negative_inputs_9_50_port, 
      negative_inputs_9_49_port, negative_inputs_9_48_port, 
      negative_inputs_9_47_port, negative_inputs_9_46_port, 
      negative_inputs_9_45_port, negative_inputs_9_44_port, 
      negative_inputs_9_43_port, negative_inputs_9_42_port, 
      negative_inputs_9_41_port, negative_inputs_9_40_port, 
      negative_inputs_9_39_port, negative_inputs_9_38_port, 
      negative_inputs_9_37_port, negative_inputs_9_36_port, 
      negative_inputs_9_35_port, negative_inputs_9_34_port, 
      negative_inputs_9_33_port, negative_inputs_9_32_port, 
      negative_inputs_9_31_port, negative_inputs_9_30_port, 
      negative_inputs_9_29_port, negative_inputs_9_28_port, 
      negative_inputs_9_27_port, negative_inputs_9_26_port, 
      negative_inputs_9_25_port, negative_inputs_9_24_port, 
      negative_inputs_9_23_port, negative_inputs_9_22_port, 
      negative_inputs_9_21_port, negative_inputs_9_20_port, 
      negative_inputs_9_19_port, negative_inputs_9_18_port, 
      negative_inputs_9_17_port, negative_inputs_9_16_port, 
      negative_inputs_9_15_port, negative_inputs_9_14_port, 
      negative_inputs_9_13_port, negative_inputs_9_12_port, 
      negative_inputs_9_11_port, negative_inputs_9_10_port, 
      negative_inputs_9_9_port, negative_inputs_9_8_port, 
      negative_inputs_9_7_port, negative_inputs_9_6_port, 
      negative_inputs_9_5_port, negative_inputs_9_4_port, 
      negative_inputs_9_3_port, negative_inputs_9_2_port, 
      negative_inputs_9_1_port, negative_inputs_24_63_port, 
      negative_inputs_24_62_port, negative_inputs_24_61_port, 
      negative_inputs_24_60_port, negative_inputs_24_59_port, 
      negative_inputs_24_58_port, negative_inputs_24_57_port, 
      negative_inputs_24_56_port, negative_inputs_24_55_port, 
      negative_inputs_24_54_port, negative_inputs_24_53_port, 
      negative_inputs_24_52_port, negative_inputs_24_51_port, 
      negative_inputs_24_50_port, negative_inputs_24_49_port, 
      negative_inputs_24_48_port, negative_inputs_24_47_port, 
      negative_inputs_24_46_port, negative_inputs_24_45_port, 
      negative_inputs_24_44_port, negative_inputs_24_43_port, 
      negative_inputs_24_42_port, negative_inputs_24_41_port, 
      negative_inputs_24_40_port, negative_inputs_24_39_port, 
      negative_inputs_24_38_port, negative_inputs_24_37_port, 
      negative_inputs_24_36_port, negative_inputs_24_35_port, 
      negative_inputs_24_34_port, negative_inputs_24_33_port, 
      negative_inputs_24_32_port, negative_inputs_24_31_port, 
      negative_inputs_24_30_port, negative_inputs_24_29_port, 
      negative_inputs_24_28_port, negative_inputs_24_27_port, 
      negative_inputs_24_26_port, negative_inputs_24_25_port, 
      negative_inputs_24_24_port, negative_inputs_24_23_port, 
      negative_inputs_24_22_port, negative_inputs_24_21_port, 
      negative_inputs_24_20_port, negative_inputs_24_19_port, 
      negative_inputs_24_18_port, negative_inputs_24_17_port, 
      negative_inputs_24_16_port, negative_inputs_24_15_port, 
      negative_inputs_24_14_port, negative_inputs_24_13_port, 
      negative_inputs_24_12_port, negative_inputs_24_11_port, 
      negative_inputs_24_10_port, negative_inputs_24_9_port, 
      negative_inputs_24_8_port, negative_inputs_24_7_port, 
      negative_inputs_24_6_port, negative_inputs_24_5_port, 
      negative_inputs_24_4_port, negative_inputs_24_3_port, 
      negative_inputs_24_2_port, negative_inputs_24_1_port, 
      negative_inputs_23_63_port, negative_inputs_23_62_port, 
      negative_inputs_23_61_port, negative_inputs_23_60_port, 
      negative_inputs_23_59_port, negative_inputs_23_58_port, 
      negative_inputs_23_57_port, negative_inputs_23_56_port, 
      negative_inputs_23_55_port, negative_inputs_23_54_port, 
      negative_inputs_23_53_port, negative_inputs_23_52_port, 
      negative_inputs_23_51_port, negative_inputs_23_50_port, 
      negative_inputs_23_49_port, negative_inputs_23_48_port, 
      negative_inputs_23_47_port, negative_inputs_23_46_port, 
      negative_inputs_23_45_port, negative_inputs_23_44_port, 
      negative_inputs_23_43_port, negative_inputs_23_42_port, 
      negative_inputs_23_41_port, negative_inputs_23_40_port, 
      negative_inputs_23_39_port, negative_inputs_23_38_port, 
      negative_inputs_23_37_port, negative_inputs_23_36_port, 
      negative_inputs_23_35_port, negative_inputs_23_34_port, 
      negative_inputs_23_33_port, negative_inputs_23_32_port, 
      negative_inputs_23_31_port, negative_inputs_23_30_port, 
      negative_inputs_23_29_port, negative_inputs_23_28_port, 
      negative_inputs_23_27_port, negative_inputs_23_26_port, 
      negative_inputs_23_25_port, negative_inputs_23_24_port, 
      negative_inputs_23_23_port, negative_inputs_23_22_port, 
      negative_inputs_23_21_port, negative_inputs_23_20_port, 
      negative_inputs_23_19_port, negative_inputs_23_18_port, 
      negative_inputs_23_17_port, negative_inputs_23_16_port, 
      negative_inputs_23_15_port, negative_inputs_23_14_port, 
      negative_inputs_23_13_port, negative_inputs_23_12_port, 
      negative_inputs_23_11_port, negative_inputs_23_10_port, 
      negative_inputs_23_9_port, negative_inputs_23_8_port, 
      negative_inputs_23_7_port, negative_inputs_23_6_port, 
      negative_inputs_23_5_port, negative_inputs_23_4_port, 
      negative_inputs_23_3_port, negative_inputs_23_2_port, 
      negative_inputs_23_1_port, negative_inputs_22_63_port, 
      negative_inputs_22_62_port, negative_inputs_22_61_port, 
      negative_inputs_22_60_port, negative_inputs_22_59_port, 
      negative_inputs_22_58_port, negative_inputs_22_57_port, 
      negative_inputs_22_56_port, negative_inputs_22_55_port, 
      negative_inputs_22_54_port, negative_inputs_22_53_port, 
      negative_inputs_22_52_port, negative_inputs_22_51_port, 
      negative_inputs_22_50_port, negative_inputs_22_49_port, 
      negative_inputs_22_48_port, negative_inputs_22_47_port, 
      negative_inputs_22_46_port, negative_inputs_22_45_port, 
      negative_inputs_22_44_port, negative_inputs_22_43_port, 
      negative_inputs_22_42_port, negative_inputs_22_41_port, 
      negative_inputs_22_40_port, negative_inputs_22_39_port, 
      negative_inputs_22_38_port, negative_inputs_22_37_port, 
      negative_inputs_22_36_port, negative_inputs_22_35_port, 
      negative_inputs_22_34_port, negative_inputs_22_33_port, 
      negative_inputs_22_32_port, negative_inputs_22_31_port, 
      negative_inputs_22_30_port, negative_inputs_22_29_port, 
      negative_inputs_22_28_port, negative_inputs_22_27_port, 
      negative_inputs_22_26_port, negative_inputs_22_25_port, 
      negative_inputs_22_24_port, negative_inputs_22_23_port, 
      negative_inputs_22_22_port, negative_inputs_22_21_port, 
      negative_inputs_22_20_port, negative_inputs_22_19_port, 
      negative_inputs_22_18_port, negative_inputs_22_17_port, 
      negative_inputs_22_16_port, negative_inputs_22_15_port, 
      negative_inputs_22_14_port, negative_inputs_22_13_port, 
      negative_inputs_22_12_port, negative_inputs_22_11_port, 
      negative_inputs_22_10_port, negative_inputs_22_9_port, 
      negative_inputs_22_8_port, negative_inputs_22_7_port, 
      negative_inputs_22_6_port, negative_inputs_22_5_port, 
      negative_inputs_22_4_port, negative_inputs_22_3_port, 
      negative_inputs_22_2_port, negative_inputs_22_1_port, 
      negative_inputs_21_63_port, negative_inputs_21_62_port, 
      negative_inputs_21_61_port, negative_inputs_21_60_port, 
      negative_inputs_21_59_port, negative_inputs_21_58_port, 
      negative_inputs_21_57_port, negative_inputs_21_56_port, 
      negative_inputs_21_55_port, negative_inputs_21_54_port, 
      negative_inputs_21_53_port, negative_inputs_21_52_port, 
      negative_inputs_21_51_port, negative_inputs_21_50_port, 
      negative_inputs_21_49_port, negative_inputs_21_48_port, 
      negative_inputs_21_47_port, negative_inputs_21_46_port, 
      negative_inputs_21_45_port, negative_inputs_21_44_port, 
      negative_inputs_21_43_port, negative_inputs_21_42_port, 
      negative_inputs_21_41_port, negative_inputs_21_40_port, 
      negative_inputs_21_39_port, negative_inputs_21_38_port, 
      negative_inputs_21_37_port, negative_inputs_21_36_port, 
      negative_inputs_21_35_port, negative_inputs_21_34_port, 
      negative_inputs_21_33_port, negative_inputs_21_32_port, 
      negative_inputs_21_31_port, negative_inputs_21_30_port, 
      negative_inputs_21_29_port, negative_inputs_21_28_port, 
      negative_inputs_21_27_port, negative_inputs_21_26_port, 
      negative_inputs_21_25_port, negative_inputs_21_24_port, 
      negative_inputs_21_23_port, negative_inputs_21_22_port, 
      negative_inputs_21_21_port, negative_inputs_21_20_port, 
      negative_inputs_21_19_port, negative_inputs_21_18_port, 
      negative_inputs_21_17_port, negative_inputs_21_16_port, 
      negative_inputs_21_15_port, negative_inputs_21_14_port, 
      negative_inputs_21_13_port, negative_inputs_21_12_port, 
      negative_inputs_21_11_port, negative_inputs_21_10_port, 
      negative_inputs_21_9_port, negative_inputs_21_8_port, 
      negative_inputs_21_7_port, negative_inputs_21_6_port, 
      negative_inputs_21_5_port, negative_inputs_21_4_port, 
      negative_inputs_21_3_port, negative_inputs_21_2_port, 
      negative_inputs_21_1_port, negative_inputs_20_63_port, 
      negative_inputs_20_62_port, negative_inputs_20_61_port, 
      negative_inputs_20_60_port, negative_inputs_20_59_port, 
      negative_inputs_20_58_port, negative_inputs_20_57_port, 
      negative_inputs_20_56_port, negative_inputs_20_55_port, 
      negative_inputs_20_54_port, negative_inputs_20_53_port, 
      negative_inputs_20_52_port, negative_inputs_20_51_port, 
      negative_inputs_20_50_port, negative_inputs_20_49_port, 
      negative_inputs_20_48_port, negative_inputs_20_47_port, 
      negative_inputs_20_46_port, negative_inputs_20_45_port, 
      negative_inputs_20_44_port, negative_inputs_20_43_port, 
      negative_inputs_20_42_port, negative_inputs_20_41_port, 
      negative_inputs_20_40_port, negative_inputs_20_39_port, 
      negative_inputs_20_38_port, negative_inputs_20_37_port, 
      negative_inputs_20_36_port, negative_inputs_20_35_port, 
      negative_inputs_20_34_port, negative_inputs_20_33_port, 
      negative_inputs_20_32_port, negative_inputs_20_31_port, 
      negative_inputs_20_30_port, negative_inputs_20_29_port, 
      negative_inputs_20_28_port, negative_inputs_20_27_port, 
      negative_inputs_20_26_port, negative_inputs_20_25_port, 
      negative_inputs_20_24_port, negative_inputs_20_23_port, 
      negative_inputs_20_22_port, negative_inputs_20_21_port, 
      negative_inputs_20_20_port, negative_inputs_20_19_port, 
      negative_inputs_20_18_port, negative_inputs_20_17_port, 
      negative_inputs_20_16_port, negative_inputs_20_15_port, 
      negative_inputs_20_14_port, negative_inputs_20_13_port, 
      negative_inputs_20_12_port, negative_inputs_20_11_port, 
      negative_inputs_20_10_port, negative_inputs_20_9_port, 
      negative_inputs_20_8_port, negative_inputs_20_7_port, 
      negative_inputs_20_6_port, negative_inputs_20_5_port, 
      negative_inputs_20_4_port, negative_inputs_20_3_port, 
      negative_inputs_20_2_port, negative_inputs_20_1_port, 
      negative_inputs_19_63_port, negative_inputs_19_62_port, 
      negative_inputs_19_61_port, negative_inputs_19_60_port, 
      negative_inputs_19_59_port, negative_inputs_19_58_port, 
      negative_inputs_19_57_port, negative_inputs_19_56_port, 
      negative_inputs_19_55_port, negative_inputs_19_54_port, 
      negative_inputs_19_53_port, negative_inputs_19_52_port, 
      negative_inputs_19_51_port, negative_inputs_19_50_port, 
      negative_inputs_19_49_port, negative_inputs_19_48_port, 
      negative_inputs_19_47_port, negative_inputs_19_46_port, 
      negative_inputs_19_45_port, negative_inputs_19_44_port, 
      negative_inputs_19_43_port, negative_inputs_19_42_port, 
      negative_inputs_19_41_port, negative_inputs_19_40_port, 
      negative_inputs_19_39_port, negative_inputs_19_38_port, 
      negative_inputs_19_37_port, negative_inputs_19_36_port, 
      negative_inputs_19_35_port, negative_inputs_19_34_port, 
      negative_inputs_19_33_port, negative_inputs_19_32_port, 
      negative_inputs_19_31_port, negative_inputs_19_30_port, 
      negative_inputs_19_29_port, negative_inputs_19_28_port, 
      negative_inputs_19_27_port, negative_inputs_19_26_port, 
      negative_inputs_19_25_port, negative_inputs_19_24_port, 
      negative_inputs_19_23_port, negative_inputs_19_22_port, 
      negative_inputs_19_21_port, negative_inputs_19_20_port, 
      negative_inputs_19_19_port, negative_inputs_19_18_port, 
      negative_inputs_19_17_port, negative_inputs_19_16_port, 
      negative_inputs_19_15_port, negative_inputs_19_14_port, 
      negative_inputs_19_13_port, negative_inputs_19_12_port, 
      negative_inputs_19_11_port, negative_inputs_19_10_port, 
      negative_inputs_19_9_port, negative_inputs_19_8_port, 
      negative_inputs_19_7_port, negative_inputs_19_6_port, 
      negative_inputs_19_5_port, negative_inputs_19_4_port, 
      negative_inputs_19_3_port, negative_inputs_19_2_port, 
      negative_inputs_19_1_port, negative_inputs_18_63_port, 
      negative_inputs_18_62_port, negative_inputs_18_61_port, 
      negative_inputs_18_60_port, negative_inputs_18_59_port, 
      negative_inputs_18_58_port, negative_inputs_18_57_port, 
      negative_inputs_18_56_port, negative_inputs_18_55_port, 
      negative_inputs_18_54_port, negative_inputs_18_53_port, 
      negative_inputs_18_52_port, negative_inputs_18_51_port, 
      negative_inputs_18_50_port, negative_inputs_18_49_port, 
      negative_inputs_18_48_port, negative_inputs_18_47_port, 
      negative_inputs_18_46_port, negative_inputs_18_45_port, 
      negative_inputs_18_44_port, negative_inputs_18_43_port, 
      negative_inputs_18_42_port, negative_inputs_18_41_port, 
      negative_inputs_18_40_port, negative_inputs_18_39_port, 
      negative_inputs_18_38_port, negative_inputs_18_37_port, 
      negative_inputs_18_36_port, negative_inputs_18_35_port, 
      negative_inputs_18_34_port, negative_inputs_18_33_port, 
      negative_inputs_18_32_port, negative_inputs_18_31_port, 
      negative_inputs_18_30_port, negative_inputs_18_29_port, 
      negative_inputs_18_28_port, negative_inputs_18_27_port, 
      negative_inputs_18_26_port, negative_inputs_18_25_port, 
      negative_inputs_18_24_port, negative_inputs_18_23_port, 
      negative_inputs_18_22_port, negative_inputs_18_21_port, 
      negative_inputs_18_20_port, negative_inputs_18_19_port, 
      negative_inputs_18_18_port, negative_inputs_18_17_port, 
      negative_inputs_18_16_port, negative_inputs_18_15_port, 
      negative_inputs_18_14_port, negative_inputs_18_13_port, 
      negative_inputs_18_12_port, negative_inputs_18_11_port, 
      negative_inputs_18_10_port, negative_inputs_18_9_port, 
      negative_inputs_18_8_port, negative_inputs_18_7_port, 
      negative_inputs_18_6_port, negative_inputs_18_5_port, 
      negative_inputs_18_4_port, negative_inputs_18_3_port, 
      negative_inputs_18_2_port, negative_inputs_18_1_port, 
      negative_inputs_17_63_port, negative_inputs_17_62_port, 
      negative_inputs_17_61_port, negative_inputs_17_60_port, 
      negative_inputs_17_59_port, negative_inputs_17_58_port, 
      negative_inputs_17_57_port, negative_inputs_17_56_port, 
      negative_inputs_17_55_port, negative_inputs_17_54_port, 
      negative_inputs_17_53_port, negative_inputs_17_52_port, 
      negative_inputs_17_51_port, negative_inputs_17_50_port, 
      negative_inputs_17_49_port, negative_inputs_17_48_port, 
      negative_inputs_17_47_port, negative_inputs_17_46_port, 
      negative_inputs_17_45_port, negative_inputs_17_44_port, 
      negative_inputs_17_43_port, negative_inputs_17_42_port, 
      negative_inputs_17_41_port, negative_inputs_17_40_port, 
      negative_inputs_17_39_port, negative_inputs_17_38_port, 
      negative_inputs_17_37_port, negative_inputs_17_36_port, 
      negative_inputs_17_35_port, negative_inputs_17_34_port, 
      negative_inputs_17_33_port, negative_inputs_17_32_port, 
      negative_inputs_17_31_port, negative_inputs_17_30_port, 
      negative_inputs_17_29_port, negative_inputs_17_28_port, 
      negative_inputs_17_27_port, negative_inputs_17_26_port, 
      negative_inputs_17_25_port, negative_inputs_17_24_port, 
      negative_inputs_17_23_port, negative_inputs_17_22_port, 
      negative_inputs_17_21_port, negative_inputs_17_20_port, 
      negative_inputs_17_19_port, negative_inputs_17_18_port, 
      negative_inputs_17_17_port, negative_inputs_17_16_port, 
      negative_inputs_17_15_port, negative_inputs_17_14_port, 
      negative_inputs_17_13_port, negative_inputs_17_12_port, 
      negative_inputs_17_11_port, negative_inputs_17_10_port, 
      negative_inputs_17_9_port, negative_inputs_17_8_port, 
      negative_inputs_17_7_port, negative_inputs_17_6_port, 
      negative_inputs_17_5_port, negative_inputs_17_4_port, 
      negative_inputs_17_3_port, negative_inputs_17_2_port, 
      negative_inputs_17_1_port, negative_inputs_31_63_port, 
      negative_inputs_31_62_port, negative_inputs_31_61_port, 
      negative_inputs_31_60_port, negative_inputs_31_59_port, 
      negative_inputs_31_58_port, negative_inputs_31_57_port, 
      negative_inputs_31_56_port, negative_inputs_31_55_port, 
      negative_inputs_31_54_port, negative_inputs_31_53_port, 
      negative_inputs_31_52_port, negative_inputs_31_51_port, 
      negative_inputs_31_50_port, negative_inputs_31_49_port, 
      negative_inputs_31_48_port, negative_inputs_31_47_port, 
      negative_inputs_31_46_port, negative_inputs_31_45_port, 
      negative_inputs_31_44_port, negative_inputs_31_43_port, 
      negative_inputs_31_42_port, negative_inputs_31_41_port, 
      negative_inputs_31_40_port, negative_inputs_31_39_port, 
      negative_inputs_31_38_port, negative_inputs_31_37_port, 
      negative_inputs_31_36_port, negative_inputs_31_35_port, 
      negative_inputs_31_34_port, negative_inputs_31_33_port, 
      negative_inputs_31_32_port, negative_inputs_31_31_port, 
      negative_inputs_31_30_port, negative_inputs_31_29_port, 
      negative_inputs_31_28_port, negative_inputs_31_27_port, 
      negative_inputs_31_26_port, negative_inputs_31_25_port, 
      negative_inputs_31_24_port, negative_inputs_31_23_port, 
      negative_inputs_31_22_port, negative_inputs_31_21_port, 
      negative_inputs_31_20_port, negative_inputs_31_19_port, 
      negative_inputs_31_18_port, negative_inputs_31_17_port, 
      negative_inputs_31_16_port, negative_inputs_31_15_port, 
      negative_inputs_31_14_port, negative_inputs_31_13_port, 
      negative_inputs_31_12_port, negative_inputs_31_11_port, 
      negative_inputs_31_10_port, negative_inputs_31_9_port, 
      negative_inputs_31_8_port, negative_inputs_31_7_port, 
      negative_inputs_31_6_port, negative_inputs_31_5_port, 
      negative_inputs_31_4_port, negative_inputs_31_3_port, 
      negative_inputs_31_2_port, negative_inputs_31_1_port, 
      negative_inputs_30_63_port, negative_inputs_30_62_port, 
      negative_inputs_30_61_port, negative_inputs_30_60_port, 
      negative_inputs_30_59_port, negative_inputs_30_58_port, 
      negative_inputs_30_57_port, negative_inputs_30_56_port, 
      negative_inputs_30_55_port, negative_inputs_30_54_port, 
      negative_inputs_30_53_port, negative_inputs_30_52_port, 
      negative_inputs_30_51_port, negative_inputs_30_50_port, 
      negative_inputs_30_49_port, negative_inputs_30_48_port, 
      negative_inputs_30_47_port, negative_inputs_30_46_port, 
      negative_inputs_30_45_port, negative_inputs_30_44_port, 
      negative_inputs_30_43_port, negative_inputs_30_42_port, 
      negative_inputs_30_41_port, negative_inputs_30_40_port, 
      negative_inputs_30_39_port, negative_inputs_30_38_port, 
      negative_inputs_30_37_port, negative_inputs_30_36_port, 
      negative_inputs_30_35_port, negative_inputs_30_34_port, 
      negative_inputs_30_33_port, negative_inputs_30_32_port, 
      negative_inputs_30_31_port, negative_inputs_30_30_port, 
      negative_inputs_30_29_port, negative_inputs_30_28_port, 
      negative_inputs_30_27_port, negative_inputs_30_26_port, 
      negative_inputs_30_25_port, negative_inputs_30_24_port, 
      negative_inputs_30_23_port, negative_inputs_30_22_port, 
      negative_inputs_30_21_port, negative_inputs_30_20_port, 
      negative_inputs_30_19_port, negative_inputs_30_18_port, 
      negative_inputs_30_17_port, negative_inputs_30_16_port, 
      negative_inputs_30_15_port, negative_inputs_30_14_port, 
      negative_inputs_30_13_port, negative_inputs_30_12_port, 
      negative_inputs_30_11_port, negative_inputs_30_10_port, 
      negative_inputs_30_9_port, negative_inputs_30_8_port, 
      negative_inputs_30_7_port, negative_inputs_30_6_port, 
      negative_inputs_30_5_port, negative_inputs_30_4_port, 
      negative_inputs_30_3_port, negative_inputs_30_2_port, 
      negative_inputs_30_1_port, negative_inputs_29_63_port, 
      negative_inputs_29_62_port, negative_inputs_29_61_port, 
      negative_inputs_29_60_port, negative_inputs_29_59_port, 
      negative_inputs_29_58_port, negative_inputs_29_57_port, 
      negative_inputs_29_56_port, negative_inputs_29_55_port, 
      negative_inputs_29_54_port, negative_inputs_29_53_port, 
      negative_inputs_29_52_port, negative_inputs_29_51_port, 
      negative_inputs_29_50_port, negative_inputs_29_49_port, 
      negative_inputs_29_48_port, negative_inputs_29_47_port, 
      negative_inputs_29_46_port, negative_inputs_29_45_port, 
      negative_inputs_29_44_port, negative_inputs_29_43_port, 
      negative_inputs_29_42_port, negative_inputs_29_41_port, 
      negative_inputs_29_40_port, negative_inputs_29_39_port, 
      negative_inputs_29_38_port, negative_inputs_29_37_port, 
      negative_inputs_29_36_port, negative_inputs_29_35_port, 
      negative_inputs_29_34_port, negative_inputs_29_33_port, 
      negative_inputs_29_32_port, negative_inputs_29_31_port, 
      negative_inputs_29_30_port, negative_inputs_29_29_port, 
      negative_inputs_29_28_port, negative_inputs_29_27_port, 
      negative_inputs_29_26_port, negative_inputs_29_25_port, 
      negative_inputs_29_24_port, negative_inputs_29_23_port, 
      negative_inputs_29_22_port, negative_inputs_29_21_port, 
      negative_inputs_29_20_port, negative_inputs_29_19_port, 
      negative_inputs_29_18_port, negative_inputs_29_17_port, 
      negative_inputs_29_16_port, negative_inputs_29_15_port, 
      negative_inputs_29_14_port, negative_inputs_29_13_port, 
      negative_inputs_29_12_port, negative_inputs_29_11_port, 
      negative_inputs_29_10_port, negative_inputs_29_9_port, 
      negative_inputs_29_8_port, negative_inputs_29_7_port, 
      negative_inputs_29_6_port, negative_inputs_29_5_port, 
      negative_inputs_29_4_port, negative_inputs_29_3_port, 
      negative_inputs_29_2_port, negative_inputs_29_1_port, 
      negative_inputs_28_63_port, negative_inputs_28_62_port, 
      negative_inputs_28_61_port, negative_inputs_28_60_port, 
      negative_inputs_28_59_port, negative_inputs_28_58_port, 
      negative_inputs_28_57_port, negative_inputs_28_56_port, 
      negative_inputs_28_55_port, negative_inputs_28_54_port, 
      negative_inputs_28_53_port, negative_inputs_28_52_port, 
      negative_inputs_28_51_port, negative_inputs_28_50_port, 
      negative_inputs_28_49_port, negative_inputs_28_48_port, 
      negative_inputs_28_47_port, negative_inputs_28_46_port, 
      negative_inputs_28_45_port, negative_inputs_28_44_port, 
      negative_inputs_28_43_port, negative_inputs_28_42_port, 
      negative_inputs_28_41_port, negative_inputs_28_40_port, 
      negative_inputs_28_39_port, negative_inputs_28_38_port, 
      negative_inputs_28_37_port, negative_inputs_28_36_port, 
      negative_inputs_28_35_port, negative_inputs_28_34_port, 
      negative_inputs_28_33_port, negative_inputs_28_32_port, 
      negative_inputs_28_31_port, negative_inputs_28_30_port, 
      negative_inputs_28_29_port, negative_inputs_28_28_port, 
      negative_inputs_28_27_port, negative_inputs_28_26_port, 
      negative_inputs_28_25_port, negative_inputs_28_24_port, 
      negative_inputs_28_23_port, negative_inputs_28_22_port, 
      negative_inputs_28_21_port, negative_inputs_28_20_port, 
      negative_inputs_28_19_port, negative_inputs_28_18_port, 
      negative_inputs_28_17_port, negative_inputs_28_16_port, 
      negative_inputs_28_15_port, negative_inputs_28_14_port, 
      negative_inputs_28_13_port, negative_inputs_28_12_port, 
      negative_inputs_28_11_port, negative_inputs_28_10_port, 
      negative_inputs_28_9_port, negative_inputs_28_8_port, 
      negative_inputs_28_7_port, negative_inputs_28_6_port, 
      negative_inputs_28_5_port, negative_inputs_28_4_port, 
      negative_inputs_28_3_port, negative_inputs_28_2_port, 
      negative_inputs_28_1_port, negative_inputs_27_63_port, 
      negative_inputs_27_62_port, negative_inputs_27_61_port, 
      negative_inputs_27_60_port, negative_inputs_27_59_port, 
      negative_inputs_27_58_port, negative_inputs_27_57_port, 
      negative_inputs_27_56_port, negative_inputs_27_55_port, 
      negative_inputs_27_54_port, negative_inputs_27_53_port, 
      negative_inputs_27_52_port, negative_inputs_27_51_port, 
      negative_inputs_27_50_port, negative_inputs_27_49_port, 
      negative_inputs_27_48_port, negative_inputs_27_47_port, 
      negative_inputs_27_46_port, negative_inputs_27_45_port, 
      negative_inputs_27_44_port, negative_inputs_27_43_port, 
      negative_inputs_27_42_port, negative_inputs_27_41_port, 
      negative_inputs_27_40_port, negative_inputs_27_39_port, 
      negative_inputs_27_38_port, negative_inputs_27_37_port, 
      negative_inputs_27_36_port, negative_inputs_27_35_port, 
      negative_inputs_27_34_port, negative_inputs_27_33_port, 
      negative_inputs_27_32_port, negative_inputs_27_31_port, 
      negative_inputs_27_30_port, negative_inputs_27_29_port, 
      negative_inputs_27_28_port, negative_inputs_27_27_port, 
      negative_inputs_27_26_port, negative_inputs_27_25_port, 
      negative_inputs_27_24_port, negative_inputs_27_23_port, 
      negative_inputs_27_22_port, negative_inputs_27_21_port, 
      negative_inputs_27_20_port, negative_inputs_27_19_port, 
      negative_inputs_27_18_port, negative_inputs_27_17_port, 
      negative_inputs_27_16_port, negative_inputs_27_15_port, 
      negative_inputs_27_14_port, negative_inputs_27_13_port, 
      negative_inputs_27_12_port, negative_inputs_27_11_port, 
      negative_inputs_27_10_port, negative_inputs_27_9_port, 
      negative_inputs_27_8_port, negative_inputs_27_7_port, 
      negative_inputs_27_6_port, negative_inputs_27_5_port, 
      negative_inputs_27_4_port, negative_inputs_27_3_port, 
      negative_inputs_27_2_port, negative_inputs_27_1_port, 
      negative_inputs_26_63_port, negative_inputs_26_62_port, 
      negative_inputs_26_61_port, negative_inputs_26_60_port, 
      negative_inputs_26_59_port, negative_inputs_26_58_port, 
      negative_inputs_26_57_port, negative_inputs_26_56_port, 
      negative_inputs_26_55_port, negative_inputs_26_54_port, 
      negative_inputs_26_53_port, negative_inputs_26_52_port, 
      negative_inputs_26_51_port, negative_inputs_26_50_port, 
      negative_inputs_26_49_port, negative_inputs_26_48_port, 
      negative_inputs_26_47_port, negative_inputs_26_46_port, 
      negative_inputs_26_45_port, negative_inputs_26_44_port, 
      negative_inputs_26_43_port, negative_inputs_26_42_port, 
      negative_inputs_26_41_port, negative_inputs_26_40_port, 
      negative_inputs_26_39_port, negative_inputs_26_38_port, 
      negative_inputs_26_37_port, negative_inputs_26_36_port, 
      negative_inputs_26_35_port, negative_inputs_26_34_port, 
      negative_inputs_26_33_port, negative_inputs_26_32_port, 
      negative_inputs_26_31_port, negative_inputs_26_30_port, 
      negative_inputs_26_29_port, negative_inputs_26_28_port, 
      negative_inputs_26_27_port, negative_inputs_26_26_port, 
      negative_inputs_26_25_port, negative_inputs_26_24_port, 
      negative_inputs_26_23_port, negative_inputs_26_22_port, 
      negative_inputs_26_21_port, negative_inputs_26_20_port, 
      negative_inputs_26_19_port, negative_inputs_26_18_port, 
      negative_inputs_26_17_port, negative_inputs_26_16_port, 
      negative_inputs_26_15_port, negative_inputs_26_14_port, 
      negative_inputs_26_13_port, negative_inputs_26_12_port, 
      negative_inputs_26_11_port, negative_inputs_26_10_port, 
      negative_inputs_26_9_port, negative_inputs_26_8_port, 
      negative_inputs_26_7_port, negative_inputs_26_6_port, 
      negative_inputs_26_5_port, negative_inputs_26_4_port, 
      negative_inputs_26_3_port, negative_inputs_26_2_port, 
      negative_inputs_26_1_port, negative_inputs_25_63_port, 
      negative_inputs_25_62_port, negative_inputs_25_61_port, 
      negative_inputs_25_60_port, negative_inputs_25_59_port, 
      negative_inputs_25_58_port, negative_inputs_25_57_port, 
      negative_inputs_25_56_port, negative_inputs_25_55_port, 
      negative_inputs_25_54_port, negative_inputs_25_53_port, 
      negative_inputs_25_52_port, negative_inputs_25_51_port, 
      negative_inputs_25_50_port, negative_inputs_25_49_port, 
      negative_inputs_25_48_port, negative_inputs_25_47_port, 
      negative_inputs_25_46_port, negative_inputs_25_45_port, 
      negative_inputs_25_44_port, negative_inputs_25_43_port, 
      negative_inputs_25_42_port, negative_inputs_25_41_port, 
      negative_inputs_25_40_port, negative_inputs_25_39_port, 
      negative_inputs_25_38_port, negative_inputs_25_37_port, 
      negative_inputs_25_36_port, negative_inputs_25_35_port, 
      negative_inputs_25_34_port, negative_inputs_25_33_port, 
      negative_inputs_25_32_port, negative_inputs_25_31_port, 
      negative_inputs_25_30_port, negative_inputs_25_29_port, 
      negative_inputs_25_28_port, negative_inputs_25_27_port, 
      negative_inputs_25_26_port, negative_inputs_25_25_port, 
      negative_inputs_25_24_port, negative_inputs_25_23_port, 
      negative_inputs_25_22_port, negative_inputs_25_21_port, 
      negative_inputs_25_20_port, negative_inputs_25_19_port, 
      negative_inputs_25_18_port, negative_inputs_25_17_port, 
      negative_inputs_25_16_port, negative_inputs_25_15_port, 
      negative_inputs_25_14_port, negative_inputs_25_13_port, 
      negative_inputs_25_12_port, negative_inputs_25_11_port, 
      negative_inputs_25_10_port, negative_inputs_25_9_port, 
      negative_inputs_25_8_port, negative_inputs_25_7_port, 
      negative_inputs_25_6_port, negative_inputs_25_5_port, 
      negative_inputs_25_4_port, negative_inputs_25_3_port, 
      negative_inputs_25_2_port, negative_inputs_25_1_port, sel_15_2_port, 
      sel_15_1_port, sel_15_0_port, sel_14_2_port, sel_14_1_port, sel_14_0_port
      , sel_13_2_port, sel_13_1_port, sel_13_0_port, sel_12_2_port, 
      sel_12_1_port, sel_12_0_port, sel_11_2_port, sel_11_1_port, sel_11_0_port
      , sel_10_2_port, sel_10_1_port, sel_10_0_port, sel_9_2_port, sel_9_1_port
      , sel_9_0_port, sel_8_2_port, sel_8_1_port, sel_8_0_port, sel_7_2_port, 
      sel_7_1_port, sel_7_0_port, sel_6_2_port, sel_6_1_port, sel_6_0_port, 
      sel_5_2_port, sel_5_1_port, sel_5_0_port, sel_4_2_port, sel_4_1_port, 
      sel_4_0_port, sel_3_2_port, sel_3_1_port, sel_3_0_port, sel_2_2_port, 
      sel_2_1_port, sel_2_0_port, sel_1_2_port, sel_1_1_port, sel_1_0_port, 
      sel_0_2_port, sel_0_1_port, sel_0_0_port, MuxOutputs_7_63_port, 
      MuxOutputs_7_62_port, MuxOutputs_7_61_port, MuxOutputs_7_60_port, 
      MuxOutputs_7_59_port, MuxOutputs_7_58_port, MuxOutputs_7_57_port, 
      MuxOutputs_7_56_port, MuxOutputs_7_55_port, MuxOutputs_7_54_port, 
      MuxOutputs_7_53_port, MuxOutputs_7_52_port, MuxOutputs_7_51_port, 
      MuxOutputs_7_50_port, MuxOutputs_7_49_port, MuxOutputs_7_48_port, 
      MuxOutputs_7_47_port, MuxOutputs_7_46_port, MuxOutputs_7_45_port, 
      MuxOutputs_7_44_port, MuxOutputs_7_43_port, MuxOutputs_7_42_port, 
      MuxOutputs_7_41_port, MuxOutputs_7_40_port, MuxOutputs_7_39_port, 
      MuxOutputs_7_38_port, MuxOutputs_7_37_port, MuxOutputs_7_36_port, 
      MuxOutputs_7_35_port, MuxOutputs_7_34_port, MuxOutputs_7_33_port, 
      MuxOutputs_7_32_port, MuxOutputs_7_31_port, MuxOutputs_7_30_port, 
      MuxOutputs_7_29_port, MuxOutputs_7_28_port, MuxOutputs_7_27_port, 
      MuxOutputs_7_26_port, MuxOutputs_7_25_port, MuxOutputs_7_24_port, 
      MuxOutputs_7_23_port, MuxOutputs_7_22_port, MuxOutputs_7_21_port, 
      MuxOutputs_7_20_port, MuxOutputs_7_19_port, MuxOutputs_7_18_port, 
      MuxOutputs_7_17_port, MuxOutputs_7_16_port, MuxOutputs_7_15_port, 
      MuxOutputs_7_14_port, MuxOutputs_7_13_port, MuxOutputs_7_12_port, 
      MuxOutputs_7_11_port, MuxOutputs_7_10_port, MuxOutputs_7_9_port, 
      MuxOutputs_7_8_port, MuxOutputs_7_7_port, MuxOutputs_7_6_port, 
      MuxOutputs_7_5_port, MuxOutputs_7_4_port, MuxOutputs_7_3_port, 
      MuxOutputs_7_2_port, MuxOutputs_7_1_port, MuxOutputs_7_0_port, 
      MuxOutputs_6_63_port, MuxOutputs_6_62_port, MuxOutputs_6_61_port, 
      MuxOutputs_6_60_port, MuxOutputs_6_59_port, MuxOutputs_6_58_port, 
      MuxOutputs_6_57_port, MuxOutputs_6_56_port, MuxOutputs_6_55_port, 
      MuxOutputs_6_54_port, MuxOutputs_6_53_port, MuxOutputs_6_52_port, 
      MuxOutputs_6_51_port, MuxOutputs_6_50_port, MuxOutputs_6_49_port, 
      MuxOutputs_6_48_port, MuxOutputs_6_47_port, MuxOutputs_6_46_port, 
      MuxOutputs_6_45_port, MuxOutputs_6_44_port, MuxOutputs_6_43_port, 
      MuxOutputs_6_42_port, MuxOutputs_6_41_port, MuxOutputs_6_40_port, 
      MuxOutputs_6_39_port, MuxOutputs_6_38_port, MuxOutputs_6_37_port, 
      MuxOutputs_6_36_port, MuxOutputs_6_35_port, MuxOutputs_6_34_port, 
      MuxOutputs_6_33_port, MuxOutputs_6_32_port, MuxOutputs_6_31_port, 
      MuxOutputs_6_30_port, MuxOutputs_6_29_port, MuxOutputs_6_28_port, 
      MuxOutputs_6_27_port, MuxOutputs_6_26_port, MuxOutputs_6_25_port, 
      MuxOutputs_6_24_port, MuxOutputs_6_23_port, MuxOutputs_6_22_port, 
      MuxOutputs_6_21_port, MuxOutputs_6_20_port, MuxOutputs_6_19_port, 
      MuxOutputs_6_18_port, MuxOutputs_6_17_port, MuxOutputs_6_16_port, 
      MuxOutputs_6_15_port, MuxOutputs_6_14_port, MuxOutputs_6_13_port, 
      MuxOutputs_6_12_port, MuxOutputs_6_11_port, MuxOutputs_6_10_port, 
      MuxOutputs_6_9_port, MuxOutputs_6_8_port, MuxOutputs_6_7_port, 
      MuxOutputs_6_6_port, MuxOutputs_6_5_port, MuxOutputs_6_4_port, 
      MuxOutputs_6_3_port, MuxOutputs_6_2_port, MuxOutputs_6_1_port, 
      MuxOutputs_6_0_port, MuxOutputs_5_63_port, MuxOutputs_5_62_port, 
      MuxOutputs_5_61_port, MuxOutputs_5_60_port, MuxOutputs_5_59_port, 
      MuxOutputs_5_58_port, MuxOutputs_5_57_port, MuxOutputs_5_56_port, 
      MuxOutputs_5_55_port, MuxOutputs_5_54_port, MuxOutputs_5_53_port, 
      MuxOutputs_5_52_port, MuxOutputs_5_51_port, MuxOutputs_5_50_port, 
      MuxOutputs_5_49_port, MuxOutputs_5_48_port, MuxOutputs_5_47_port, 
      MuxOutputs_5_46_port, MuxOutputs_5_45_port, MuxOutputs_5_44_port, 
      MuxOutputs_5_43_port, MuxOutputs_5_42_port, MuxOutputs_5_41_port, 
      MuxOutputs_5_40_port, MuxOutputs_5_39_port, MuxOutputs_5_38_port, 
      MuxOutputs_5_37_port, MuxOutputs_5_36_port, MuxOutputs_5_35_port, 
      MuxOutputs_5_34_port, MuxOutputs_5_33_port, MuxOutputs_5_32_port, 
      MuxOutputs_5_31_port, MuxOutputs_5_30_port, MuxOutputs_5_29_port, 
      MuxOutputs_5_28_port, MuxOutputs_5_27_port, MuxOutputs_5_26_port, 
      MuxOutputs_5_25_port, MuxOutputs_5_24_port, MuxOutputs_5_23_port, 
      MuxOutputs_5_22_port, MuxOutputs_5_21_port, MuxOutputs_5_20_port, 
      MuxOutputs_5_19_port, MuxOutputs_5_18_port, MuxOutputs_5_17_port, 
      MuxOutputs_5_16_port, MuxOutputs_5_15_port, MuxOutputs_5_14_port, 
      MuxOutputs_5_13_port, MuxOutputs_5_12_port, MuxOutputs_5_11_port, 
      MuxOutputs_5_10_port, MuxOutputs_5_9_port, MuxOutputs_5_8_port, 
      MuxOutputs_5_7_port, MuxOutputs_5_6_port, MuxOutputs_5_5_port, 
      MuxOutputs_5_4_port, MuxOutputs_5_3_port, MuxOutputs_5_2_port, 
      MuxOutputs_5_1_port, MuxOutputs_5_0_port, MuxOutputs_4_63_port, 
      MuxOutputs_4_62_port, MuxOutputs_4_61_port, MuxOutputs_4_60_port, 
      MuxOutputs_4_59_port, MuxOutputs_4_58_port, MuxOutputs_4_57_port, 
      MuxOutputs_4_56_port, MuxOutputs_4_55_port, MuxOutputs_4_54_port, 
      MuxOutputs_4_53_port, MuxOutputs_4_52_port, MuxOutputs_4_51_port, 
      MuxOutputs_4_50_port, MuxOutputs_4_49_port, MuxOutputs_4_48_port, 
      MuxOutputs_4_47_port, MuxOutputs_4_46_port, MuxOutputs_4_45_port, 
      MuxOutputs_4_44_port, MuxOutputs_4_43_port, MuxOutputs_4_42_port, 
      MuxOutputs_4_41_port, MuxOutputs_4_40_port, MuxOutputs_4_39_port, 
      MuxOutputs_4_38_port, MuxOutputs_4_37_port, MuxOutputs_4_36_port, 
      MuxOutputs_4_35_port, MuxOutputs_4_34_port, MuxOutputs_4_33_port, 
      MuxOutputs_4_32_port, MuxOutputs_4_31_port, MuxOutputs_4_30_port, 
      MuxOutputs_4_29_port, MuxOutputs_4_28_port, MuxOutputs_4_27_port, 
      MuxOutputs_4_26_port, MuxOutputs_4_25_port, MuxOutputs_4_24_port, 
      MuxOutputs_4_23_port, MuxOutputs_4_22_port, MuxOutputs_4_21_port, 
      MuxOutputs_4_20_port, MuxOutputs_4_19_port, MuxOutputs_4_18_port, 
      MuxOutputs_4_17_port, MuxOutputs_4_16_port, MuxOutputs_4_15_port, 
      MuxOutputs_4_14_port, MuxOutputs_4_13_port, MuxOutputs_4_12_port, 
      MuxOutputs_4_11_port, MuxOutputs_4_10_port, MuxOutputs_4_9_port, 
      MuxOutputs_4_8_port, MuxOutputs_4_7_port, MuxOutputs_4_6_port, 
      MuxOutputs_4_5_port, MuxOutputs_4_4_port, MuxOutputs_4_3_port, 
      MuxOutputs_4_2_port, MuxOutputs_4_1_port, MuxOutputs_4_0_port, 
      MuxOutputs_3_63_port, MuxOutputs_3_62_port, MuxOutputs_3_61_port, 
      MuxOutputs_3_60_port, MuxOutputs_3_59_port, MuxOutputs_3_58_port, 
      MuxOutputs_3_57_port, MuxOutputs_3_56_port, MuxOutputs_3_55_port, 
      MuxOutputs_3_54_port, MuxOutputs_3_53_port, MuxOutputs_3_52_port, 
      MuxOutputs_3_51_port, MuxOutputs_3_50_port, MuxOutputs_3_49_port, 
      MuxOutputs_3_48_port, MuxOutputs_3_47_port, MuxOutputs_3_46_port, 
      MuxOutputs_3_45_port, MuxOutputs_3_44_port, MuxOutputs_3_43_port, 
      MuxOutputs_3_42_port, MuxOutputs_3_41_port, MuxOutputs_3_40_port, 
      MuxOutputs_3_39_port, MuxOutputs_3_38_port, MuxOutputs_3_37_port, 
      MuxOutputs_3_36_port, MuxOutputs_3_35_port, MuxOutputs_3_34_port, 
      MuxOutputs_3_33_port, MuxOutputs_3_32_port, MuxOutputs_3_31_port, 
      MuxOutputs_3_30_port, MuxOutputs_3_29_port, MuxOutputs_3_28_port, 
      MuxOutputs_3_27_port, MuxOutputs_3_26_port, MuxOutputs_3_25_port, 
      MuxOutputs_3_24_port, MuxOutputs_3_23_port, MuxOutputs_3_22_port, 
      MuxOutputs_3_21_port, MuxOutputs_3_20_port, MuxOutputs_3_19_port, 
      MuxOutputs_3_18_port, MuxOutputs_3_17_port, MuxOutputs_3_16_port, 
      MuxOutputs_3_15_port, MuxOutputs_3_14_port, MuxOutputs_3_13_port, 
      MuxOutputs_3_12_port, MuxOutputs_3_11_port, MuxOutputs_3_10_port, 
      MuxOutputs_3_9_port, MuxOutputs_3_8_port, MuxOutputs_3_7_port, 
      MuxOutputs_3_6_port, MuxOutputs_3_5_port, MuxOutputs_3_4_port, 
      MuxOutputs_3_3_port, MuxOutputs_3_2_port, MuxOutputs_3_1_port, 
      MuxOutputs_3_0_port, MuxOutputs_2_63_port, MuxOutputs_2_62_port, 
      MuxOutputs_2_61_port, MuxOutputs_2_60_port, MuxOutputs_2_59_port, 
      MuxOutputs_2_58_port, MuxOutputs_2_57_port, MuxOutputs_2_56_port, 
      MuxOutputs_2_55_port, MuxOutputs_2_54_port, MuxOutputs_2_53_port, 
      MuxOutputs_2_52_port, MuxOutputs_2_51_port, MuxOutputs_2_50_port, 
      MuxOutputs_2_49_port, MuxOutputs_2_48_port, MuxOutputs_2_47_port, 
      MuxOutputs_2_46_port, MuxOutputs_2_45_port, MuxOutputs_2_44_port, 
      MuxOutputs_2_43_port, MuxOutputs_2_42_port, MuxOutputs_2_41_port, 
      MuxOutputs_2_40_port, MuxOutputs_2_39_port, MuxOutputs_2_38_port, 
      MuxOutputs_2_37_port, MuxOutputs_2_36_port, MuxOutputs_2_35_port, 
      MuxOutputs_2_34_port, MuxOutputs_2_33_port, MuxOutputs_2_32_port, 
      MuxOutputs_2_31_port, MuxOutputs_2_30_port, MuxOutputs_2_29_port, 
      MuxOutputs_2_28_port, MuxOutputs_2_27_port, MuxOutputs_2_26_port, 
      MuxOutputs_2_25_port, MuxOutputs_2_24_port, MuxOutputs_2_23_port, 
      MuxOutputs_2_22_port, MuxOutputs_2_21_port, MuxOutputs_2_20_port, 
      MuxOutputs_2_19_port, MuxOutputs_2_18_port, MuxOutputs_2_17_port, 
      MuxOutputs_2_16_port, MuxOutputs_2_15_port, MuxOutputs_2_14_port, 
      MuxOutputs_2_13_port, MuxOutputs_2_12_port, MuxOutputs_2_11_port, 
      MuxOutputs_2_10_port, MuxOutputs_2_9_port, MuxOutputs_2_8_port, 
      MuxOutputs_2_7_port, MuxOutputs_2_6_port, MuxOutputs_2_5_port, 
      MuxOutputs_2_4_port, MuxOutputs_2_3_port, MuxOutputs_2_2_port, 
      MuxOutputs_2_1_port, MuxOutputs_2_0_port, MuxOutputs_1_63_port, 
      MuxOutputs_1_62_port, MuxOutputs_1_61_port, MuxOutputs_1_60_port, 
      MuxOutputs_1_59_port, MuxOutputs_1_58_port, MuxOutputs_1_57_port, 
      MuxOutputs_1_56_port, MuxOutputs_1_55_port, MuxOutputs_1_54_port, 
      MuxOutputs_1_53_port, MuxOutputs_1_52_port, MuxOutputs_1_51_port, 
      MuxOutputs_1_50_port, MuxOutputs_1_49_port, MuxOutputs_1_48_port, 
      MuxOutputs_1_47_port, MuxOutputs_1_46_port, MuxOutputs_1_45_port, 
      MuxOutputs_1_44_port, MuxOutputs_1_43_port, MuxOutputs_1_42_port, 
      MuxOutputs_1_41_port, MuxOutputs_1_40_port, MuxOutputs_1_39_port, 
      MuxOutputs_1_38_port, MuxOutputs_1_37_port, MuxOutputs_1_36_port, 
      MuxOutputs_1_35_port, MuxOutputs_1_34_port, MuxOutputs_1_33_port, 
      MuxOutputs_1_32_port, MuxOutputs_1_31_port, MuxOutputs_1_30_port, 
      MuxOutputs_1_29_port, MuxOutputs_1_28_port, MuxOutputs_1_27_port, 
      MuxOutputs_1_26_port, MuxOutputs_1_25_port, MuxOutputs_1_24_port, 
      MuxOutputs_1_23_port, MuxOutputs_1_22_port, MuxOutputs_1_21_port, 
      MuxOutputs_1_20_port, MuxOutputs_1_19_port, MuxOutputs_1_18_port, 
      MuxOutputs_1_17_port, MuxOutputs_1_16_port, MuxOutputs_1_15_port, 
      MuxOutputs_1_14_port, MuxOutputs_1_13_port, MuxOutputs_1_12_port, 
      MuxOutputs_1_11_port, MuxOutputs_1_10_port, MuxOutputs_1_9_port, 
      MuxOutputs_1_8_port, MuxOutputs_1_7_port, MuxOutputs_1_6_port, 
      MuxOutputs_1_5_port, MuxOutputs_1_4_port, MuxOutputs_1_3_port, 
      MuxOutputs_1_2_port, MuxOutputs_1_1_port, MuxOutputs_1_0_port, 
      MuxOutputs_0_63_port, MuxOutputs_0_62_port, MuxOutputs_0_61_port, 
      MuxOutputs_0_60_port, MuxOutputs_0_59_port, MuxOutputs_0_58_port, 
      MuxOutputs_0_57_port, MuxOutputs_0_56_port, MuxOutputs_0_55_port, 
      MuxOutputs_0_54_port, MuxOutputs_0_53_port, MuxOutputs_0_52_port, 
      MuxOutputs_0_51_port, MuxOutputs_0_50_port, MuxOutputs_0_49_port, 
      MuxOutputs_0_48_port, MuxOutputs_0_47_port, MuxOutputs_0_46_port, 
      MuxOutputs_0_45_port, MuxOutputs_0_44_port, MuxOutputs_0_43_port, 
      MuxOutputs_0_42_port, MuxOutputs_0_41_port, MuxOutputs_0_40_port, 
      MuxOutputs_0_39_port, MuxOutputs_0_38_port, MuxOutputs_0_37_port, 
      MuxOutputs_0_36_port, MuxOutputs_0_35_port, MuxOutputs_0_34_port, 
      MuxOutputs_0_33_port, MuxOutputs_0_32_port, MuxOutputs_0_31_port, 
      MuxOutputs_0_30_port, MuxOutputs_0_29_port, MuxOutputs_0_28_port, 
      MuxOutputs_0_27_port, MuxOutputs_0_26_port, MuxOutputs_0_25_port, 
      MuxOutputs_0_24_port, MuxOutputs_0_23_port, MuxOutputs_0_22_port, 
      MuxOutputs_0_21_port, MuxOutputs_0_20_port, MuxOutputs_0_19_port, 
      MuxOutputs_0_18_port, MuxOutputs_0_17_port, MuxOutputs_0_16_port, 
      MuxOutputs_0_15_port, MuxOutputs_0_14_port, MuxOutputs_0_13_port, 
      MuxOutputs_0_12_port, MuxOutputs_0_11_port, MuxOutputs_0_10_port, 
      MuxOutputs_0_9_port, MuxOutputs_0_8_port, MuxOutputs_0_7_port, 
      MuxOutputs_0_6_port, MuxOutputs_0_5_port, MuxOutputs_0_4_port, 
      MuxOutputs_0_3_port, MuxOutputs_0_2_port, MuxOutputs_0_1_port, 
      MuxOutputs_0_0_port, MuxOutputs_15_63_port, MuxOutputs_15_62_port, 
      MuxOutputs_15_61_port, MuxOutputs_15_60_port, MuxOutputs_15_59_port, 
      MuxOutputs_15_58_port, MuxOutputs_15_57_port, MuxOutputs_15_56_port, 
      MuxOutputs_15_55_port, MuxOutputs_15_54_port, MuxOutputs_15_53_port, 
      MuxOutputs_15_52_port, MuxOutputs_15_51_port, MuxOutputs_15_50_port, 
      MuxOutputs_15_49_port, MuxOutputs_15_48_port, MuxOutputs_15_47_port, 
      MuxOutputs_15_46_port, MuxOutputs_15_45_port, MuxOutputs_15_44_port, 
      MuxOutputs_15_43_port, MuxOutputs_15_42_port, MuxOutputs_15_41_port, 
      MuxOutputs_15_40_port, MuxOutputs_15_39_port, MuxOutputs_15_38_port, 
      MuxOutputs_15_37_port, MuxOutputs_15_36_port, MuxOutputs_15_35_port, 
      MuxOutputs_15_34_port, MuxOutputs_15_33_port, MuxOutputs_15_32_port, 
      MuxOutputs_15_31_port, MuxOutputs_15_30_port, MuxOutputs_15_29_port, 
      MuxOutputs_15_28_port, MuxOutputs_15_27_port, MuxOutputs_15_26_port, 
      MuxOutputs_15_25_port, MuxOutputs_15_24_port, MuxOutputs_15_23_port, 
      MuxOutputs_15_22_port, MuxOutputs_15_21_port, MuxOutputs_15_20_port, 
      MuxOutputs_15_19_port, MuxOutputs_15_18_port, MuxOutputs_15_17_port, 
      MuxOutputs_15_16_port, MuxOutputs_15_15_port, MuxOutputs_15_14_port, 
      MuxOutputs_15_13_port, MuxOutputs_15_12_port, MuxOutputs_15_11_port, 
      MuxOutputs_15_10_port, MuxOutputs_15_9_port, MuxOutputs_15_8_port, 
      MuxOutputs_15_7_port, MuxOutputs_15_6_port, MuxOutputs_15_5_port, 
      MuxOutputs_15_4_port, MuxOutputs_15_3_port, MuxOutputs_15_2_port, 
      MuxOutputs_15_1_port, MuxOutputs_15_0_port, MuxOutputs_14_63_port, 
      MuxOutputs_14_62_port, MuxOutputs_14_61_port, MuxOutputs_14_60_port, 
      MuxOutputs_14_59_port, MuxOutputs_14_58_port, MuxOutputs_14_57_port, 
      MuxOutputs_14_56_port, MuxOutputs_14_55_port, MuxOutputs_14_54_port, 
      MuxOutputs_14_53_port, MuxOutputs_14_52_port, MuxOutputs_14_51_port, 
      MuxOutputs_14_50_port, MuxOutputs_14_49_port, MuxOutputs_14_48_port, 
      MuxOutputs_14_47_port, MuxOutputs_14_46_port, MuxOutputs_14_45_port, 
      MuxOutputs_14_44_port, MuxOutputs_14_43_port, MuxOutputs_14_42_port, 
      MuxOutputs_14_41_port, MuxOutputs_14_40_port, MuxOutputs_14_39_port, 
      MuxOutputs_14_38_port, MuxOutputs_14_37_port, MuxOutputs_14_36_port, 
      MuxOutputs_14_35_port, MuxOutputs_14_34_port, MuxOutputs_14_33_port, 
      MuxOutputs_14_32_port, MuxOutputs_14_31_port, MuxOutputs_14_30_port, 
      MuxOutputs_14_29_port, MuxOutputs_14_28_port, MuxOutputs_14_27_port, 
      MuxOutputs_14_26_port, MuxOutputs_14_25_port, MuxOutputs_14_24_port, 
      MuxOutputs_14_23_port, MuxOutputs_14_22_port, MuxOutputs_14_21_port, 
      MuxOutputs_14_20_port, MuxOutputs_14_19_port, MuxOutputs_14_18_port, 
      MuxOutputs_14_17_port, MuxOutputs_14_16_port, MuxOutputs_14_15_port, 
      MuxOutputs_14_14_port, MuxOutputs_14_13_port, MuxOutputs_14_12_port, 
      MuxOutputs_14_11_port, MuxOutputs_14_10_port, MuxOutputs_14_9_port, 
      MuxOutputs_14_8_port, MuxOutputs_14_7_port, MuxOutputs_14_6_port, 
      MuxOutputs_14_5_port, MuxOutputs_14_4_port, MuxOutputs_14_3_port, 
      MuxOutputs_14_2_port, MuxOutputs_14_1_port, MuxOutputs_14_0_port, 
      MuxOutputs_13_63_port, MuxOutputs_13_62_port, MuxOutputs_13_61_port, 
      MuxOutputs_13_60_port, MuxOutputs_13_59_port, MuxOutputs_13_58_port, 
      MuxOutputs_13_57_port, MuxOutputs_13_56_port, MuxOutputs_13_55_port, 
      MuxOutputs_13_54_port, MuxOutputs_13_53_port, MuxOutputs_13_52_port, 
      MuxOutputs_13_51_port, MuxOutputs_13_50_port, MuxOutputs_13_49_port, 
      MuxOutputs_13_48_port, MuxOutputs_13_47_port, MuxOutputs_13_46_port, 
      MuxOutputs_13_45_port, MuxOutputs_13_44_port, MuxOutputs_13_43_port, 
      MuxOutputs_13_42_port, MuxOutputs_13_41_port, MuxOutputs_13_40_port, 
      MuxOutputs_13_39_port, MuxOutputs_13_38_port, MuxOutputs_13_37_port, 
      MuxOutputs_13_36_port, MuxOutputs_13_35_port, MuxOutputs_13_34_port, 
      MuxOutputs_13_33_port, MuxOutputs_13_32_port, MuxOutputs_13_31_port, 
      MuxOutputs_13_30_port, MuxOutputs_13_29_port, MuxOutputs_13_28_port, 
      MuxOutputs_13_27_port, MuxOutputs_13_26_port, MuxOutputs_13_25_port, 
      MuxOutputs_13_24_port, MuxOutputs_13_23_port, MuxOutputs_13_22_port, 
      MuxOutputs_13_21_port, MuxOutputs_13_20_port, MuxOutputs_13_19_port, 
      MuxOutputs_13_18_port, MuxOutputs_13_17_port, MuxOutputs_13_16_port, 
      MuxOutputs_13_15_port, MuxOutputs_13_14_port, MuxOutputs_13_13_port, 
      MuxOutputs_13_12_port, MuxOutputs_13_11_port, MuxOutputs_13_10_port, 
      MuxOutputs_13_9_port, MuxOutputs_13_8_port, MuxOutputs_13_7_port, 
      MuxOutputs_13_6_port, MuxOutputs_13_5_port, MuxOutputs_13_4_port, 
      MuxOutputs_13_3_port, MuxOutputs_13_2_port, MuxOutputs_13_1_port, 
      MuxOutputs_13_0_port, MuxOutputs_12_63_port, MuxOutputs_12_62_port, 
      MuxOutputs_12_61_port, MuxOutputs_12_60_port, MuxOutputs_12_59_port, 
      MuxOutputs_12_58_port, MuxOutputs_12_57_port, MuxOutputs_12_56_port, 
      MuxOutputs_12_55_port, MuxOutputs_12_54_port, MuxOutputs_12_53_port, 
      MuxOutputs_12_52_port, MuxOutputs_12_51_port, MuxOutputs_12_50_port, 
      MuxOutputs_12_49_port, MuxOutputs_12_48_port, MuxOutputs_12_47_port, 
      MuxOutputs_12_46_port, MuxOutputs_12_45_port, MuxOutputs_12_44_port, 
      MuxOutputs_12_43_port, MuxOutputs_12_42_port, MuxOutputs_12_41_port, 
      MuxOutputs_12_40_port, MuxOutputs_12_39_port, MuxOutputs_12_38_port, 
      MuxOutputs_12_37_port, MuxOutputs_12_36_port, MuxOutputs_12_35_port, 
      MuxOutputs_12_34_port, MuxOutputs_12_33_port, MuxOutputs_12_32_port, 
      MuxOutputs_12_31_port, MuxOutputs_12_30_port, MuxOutputs_12_29_port, 
      MuxOutputs_12_28_port, MuxOutputs_12_27_port, MuxOutputs_12_26_port, 
      MuxOutputs_12_25_port, MuxOutputs_12_24_port, MuxOutputs_12_23_port, 
      MuxOutputs_12_22_port, MuxOutputs_12_21_port, MuxOutputs_12_20_port, 
      MuxOutputs_12_19_port, MuxOutputs_12_18_port, MuxOutputs_12_17_port, 
      MuxOutputs_12_16_port, MuxOutputs_12_15_port, MuxOutputs_12_14_port, 
      MuxOutputs_12_13_port, MuxOutputs_12_12_port, MuxOutputs_12_11_port, 
      MuxOutputs_12_10_port, MuxOutputs_12_9_port, MuxOutputs_12_8_port, 
      MuxOutputs_12_7_port, MuxOutputs_12_6_port, MuxOutputs_12_5_port, 
      MuxOutputs_12_4_port, MuxOutputs_12_3_port, MuxOutputs_12_2_port, 
      MuxOutputs_12_1_port, MuxOutputs_12_0_port, MuxOutputs_11_63_port, 
      MuxOutputs_11_62_port, MuxOutputs_11_61_port, MuxOutputs_11_60_port, 
      MuxOutputs_11_59_port, MuxOutputs_11_58_port, MuxOutputs_11_57_port, 
      MuxOutputs_11_56_port, MuxOutputs_11_55_port, MuxOutputs_11_54_port, 
      MuxOutputs_11_53_port, MuxOutputs_11_52_port, MuxOutputs_11_51_port, 
      MuxOutputs_11_50_port, MuxOutputs_11_49_port, MuxOutputs_11_48_port, 
      MuxOutputs_11_47_port, MuxOutputs_11_46_port, MuxOutputs_11_45_port, 
      MuxOutputs_11_44_port, MuxOutputs_11_43_port, MuxOutputs_11_42_port, 
      MuxOutputs_11_41_port, MuxOutputs_11_40_port, MuxOutputs_11_39_port, 
      MuxOutputs_11_38_port, MuxOutputs_11_37_port, MuxOutputs_11_36_port, 
      MuxOutputs_11_35_port, MuxOutputs_11_34_port, MuxOutputs_11_33_port, 
      MuxOutputs_11_32_port, MuxOutputs_11_31_port, MuxOutputs_11_30_port, 
      MuxOutputs_11_29_port, MuxOutputs_11_28_port, MuxOutputs_11_27_port, 
      MuxOutputs_11_26_port, MuxOutputs_11_25_port, MuxOutputs_11_24_port, 
      MuxOutputs_11_23_port, MuxOutputs_11_22_port, MuxOutputs_11_21_port, 
      MuxOutputs_11_20_port, MuxOutputs_11_19_port, MuxOutputs_11_18_port, 
      MuxOutputs_11_17_port, MuxOutputs_11_16_port, MuxOutputs_11_15_port, 
      MuxOutputs_11_14_port, MuxOutputs_11_13_port, MuxOutputs_11_12_port, 
      MuxOutputs_11_11_port, MuxOutputs_11_10_port, MuxOutputs_11_9_port, 
      MuxOutputs_11_8_port, MuxOutputs_11_7_port, MuxOutputs_11_6_port, 
      MuxOutputs_11_5_port, MuxOutputs_11_4_port, MuxOutputs_11_3_port, 
      MuxOutputs_11_2_port, MuxOutputs_11_1_port, MuxOutputs_11_0_port, 
      MuxOutputs_10_63_port, MuxOutputs_10_62_port, MuxOutputs_10_61_port, 
      MuxOutputs_10_60_port, MuxOutputs_10_59_port, MuxOutputs_10_58_port, 
      MuxOutputs_10_57_port, MuxOutputs_10_56_port, MuxOutputs_10_55_port, 
      MuxOutputs_10_54_port, MuxOutputs_10_53_port, MuxOutputs_10_52_port, 
      MuxOutputs_10_51_port, MuxOutputs_10_50_port, MuxOutputs_10_49_port, 
      MuxOutputs_10_48_port, MuxOutputs_10_47_port, MuxOutputs_10_46_port, 
      MuxOutputs_10_45_port, MuxOutputs_10_44_port, MuxOutputs_10_43_port, 
      MuxOutputs_10_42_port, MuxOutputs_10_41_port, MuxOutputs_10_40_port, 
      MuxOutputs_10_39_port, MuxOutputs_10_38_port, MuxOutputs_10_37_port, 
      MuxOutputs_10_36_port, MuxOutputs_10_35_port, MuxOutputs_10_34_port, 
      MuxOutputs_10_33_port, MuxOutputs_10_32_port, MuxOutputs_10_31_port, 
      MuxOutputs_10_30_port, MuxOutputs_10_29_port, MuxOutputs_10_28_port, 
      MuxOutputs_10_27_port, MuxOutputs_10_26_port, MuxOutputs_10_25_port, 
      MuxOutputs_10_24_port, MuxOutputs_10_23_port, MuxOutputs_10_22_port, 
      MuxOutputs_10_21_port, MuxOutputs_10_20_port, MuxOutputs_10_19_port, 
      MuxOutputs_10_18_port, MuxOutputs_10_17_port, MuxOutputs_10_16_port, 
      MuxOutputs_10_15_port, MuxOutputs_10_14_port, MuxOutputs_10_13_port, 
      MuxOutputs_10_12_port, MuxOutputs_10_11_port, MuxOutputs_10_10_port, 
      MuxOutputs_10_9_port, MuxOutputs_10_8_port, MuxOutputs_10_7_port, 
      MuxOutputs_10_6_port, MuxOutputs_10_5_port, MuxOutputs_10_4_port, 
      MuxOutputs_10_3_port, MuxOutputs_10_2_port, MuxOutputs_10_1_port, 
      MuxOutputs_10_0_port, MuxOutputs_9_63_port, MuxOutputs_9_62_port, 
      MuxOutputs_9_61_port, MuxOutputs_9_60_port, MuxOutputs_9_59_port, 
      MuxOutputs_9_58_port, MuxOutputs_9_57_port, MuxOutputs_9_56_port, 
      MuxOutputs_9_55_port, MuxOutputs_9_54_port, MuxOutputs_9_53_port, 
      MuxOutputs_9_52_port, MuxOutputs_9_51_port, MuxOutputs_9_50_port, 
      MuxOutputs_9_49_port, MuxOutputs_9_48_port, MuxOutputs_9_47_port, 
      MuxOutputs_9_46_port, MuxOutputs_9_45_port, MuxOutputs_9_44_port, 
      MuxOutputs_9_43_port, MuxOutputs_9_42_port, MuxOutputs_9_41_port, 
      MuxOutputs_9_40_port, MuxOutputs_9_39_port, MuxOutputs_9_38_port, 
      MuxOutputs_9_37_port, MuxOutputs_9_36_port, MuxOutputs_9_35_port, 
      MuxOutputs_9_34_port, MuxOutputs_9_33_port, MuxOutputs_9_32_port, 
      MuxOutputs_9_31_port, MuxOutputs_9_30_port, MuxOutputs_9_29_port, 
      MuxOutputs_9_28_port, MuxOutputs_9_27_port, MuxOutputs_9_26_port, 
      MuxOutputs_9_25_port, MuxOutputs_9_24_port, MuxOutputs_9_23_port, 
      MuxOutputs_9_22_port, MuxOutputs_9_21_port, MuxOutputs_9_20_port, 
      MuxOutputs_9_19_port, MuxOutputs_9_18_port, MuxOutputs_9_17_port, 
      MuxOutputs_9_16_port, MuxOutputs_9_15_port, MuxOutputs_9_14_port, 
      MuxOutputs_9_13_port, MuxOutputs_9_12_port, MuxOutputs_9_11_port, 
      MuxOutputs_9_10_port, MuxOutputs_9_9_port, MuxOutputs_9_8_port, 
      MuxOutputs_9_7_port, MuxOutputs_9_6_port, MuxOutputs_9_5_port, 
      MuxOutputs_9_4_port, MuxOutputs_9_3_port, MuxOutputs_9_2_port, 
      MuxOutputs_9_1_port, MuxOutputs_9_0_port, MuxOutputs_8_63_port, 
      MuxOutputs_8_62_port, MuxOutputs_8_61_port, MuxOutputs_8_60_port, 
      MuxOutputs_8_59_port, MuxOutputs_8_58_port, MuxOutputs_8_57_port, 
      MuxOutputs_8_56_port, MuxOutputs_8_55_port, MuxOutputs_8_54_port, 
      MuxOutputs_8_53_port, MuxOutputs_8_52_port, MuxOutputs_8_51_port, 
      MuxOutputs_8_50_port, MuxOutputs_8_49_port, MuxOutputs_8_48_port, 
      MuxOutputs_8_47_port, MuxOutputs_8_46_port, MuxOutputs_8_45_port, 
      MuxOutputs_8_44_port, MuxOutputs_8_43_port, MuxOutputs_8_42_port, 
      MuxOutputs_8_41_port, MuxOutputs_8_40_port, MuxOutputs_8_39_port, 
      MuxOutputs_8_38_port, MuxOutputs_8_37_port, MuxOutputs_8_36_port, 
      MuxOutputs_8_35_port, MuxOutputs_8_34_port, MuxOutputs_8_33_port, 
      MuxOutputs_8_32_port, MuxOutputs_8_31_port, MuxOutputs_8_30_port, 
      MuxOutputs_8_29_port, MuxOutputs_8_28_port, MuxOutputs_8_27_port, 
      MuxOutputs_8_26_port, MuxOutputs_8_25_port, MuxOutputs_8_24_port, 
      MuxOutputs_8_23_port, MuxOutputs_8_22_port, MuxOutputs_8_21_port, 
      MuxOutputs_8_20_port, MuxOutputs_8_19_port, MuxOutputs_8_18_port, 
      MuxOutputs_8_17_port, MuxOutputs_8_16_port, MuxOutputs_8_15_port, 
      MuxOutputs_8_14_port, MuxOutputs_8_13_port, MuxOutputs_8_12_port, 
      MuxOutputs_8_11_port, MuxOutputs_8_10_port, MuxOutputs_8_9_port, 
      MuxOutputs_8_8_port, MuxOutputs_8_7_port, MuxOutputs_8_6_port, 
      MuxOutputs_8_5_port, MuxOutputs_8_4_port, MuxOutputs_8_3_port, 
      MuxOutputs_8_2_port, MuxOutputs_8_1_port, MuxOutputs_8_0_port, 
      SumOutputs_7_63_port, SumOutputs_7_62_port, SumOutputs_7_61_port, 
      SumOutputs_7_60_port, SumOutputs_7_59_port, SumOutputs_7_58_port, 
      SumOutputs_7_57_port, SumOutputs_7_56_port, SumOutputs_7_55_port, 
      SumOutputs_7_54_port, SumOutputs_7_53_port, SumOutputs_7_52_port, 
      SumOutputs_7_51_port, SumOutputs_7_50_port, SumOutputs_7_49_port, 
      SumOutputs_7_48_port, SumOutputs_7_47_port, SumOutputs_7_46_port, 
      SumOutputs_7_45_port, SumOutputs_7_44_port, SumOutputs_7_43_port, 
      SumOutputs_7_42_port, SumOutputs_7_41_port, SumOutputs_7_40_port, 
      SumOutputs_7_39_port, SumOutputs_7_38_port, SumOutputs_7_37_port, 
      SumOutputs_7_36_port, SumOutputs_7_35_port, SumOutputs_7_34_port, 
      SumOutputs_7_33_port, SumOutputs_7_32_port, SumOutputs_7_31_port, 
      SumOutputs_7_30_port, SumOutputs_7_29_port, SumOutputs_7_28_port, 
      SumOutputs_7_27_port, SumOutputs_7_26_port, SumOutputs_7_25_port, 
      SumOutputs_7_24_port, SumOutputs_7_23_port, SumOutputs_7_22_port, 
      SumOutputs_7_21_port, SumOutputs_7_20_port, SumOutputs_7_19_port, 
      SumOutputs_7_18_port, SumOutputs_7_17_port, SumOutputs_7_16_port, 
      SumOutputs_7_15_port, SumOutputs_7_14_port, SumOutputs_7_13_port, 
      SumOutputs_7_12_port, SumOutputs_7_11_port, SumOutputs_7_10_port, 
      SumOutputs_7_9_port, SumOutputs_7_8_port, SumOutputs_7_7_port, 
      SumOutputs_7_6_port, SumOutputs_7_5_port, SumOutputs_7_4_port, 
      SumOutputs_7_3_port, SumOutputs_7_2_port, SumOutputs_7_1_port, 
      SumOutputs_7_0_port, SumOutputs_6_63_port, SumOutputs_6_62_port, 
      SumOutputs_6_61_port, SumOutputs_6_60_port, SumOutputs_6_59_port, 
      SumOutputs_6_58_port, SumOutputs_6_57_port, SumOutputs_6_56_port, 
      SumOutputs_6_55_port, SumOutputs_6_54_port, SumOutputs_6_53_port, 
      SumOutputs_6_52_port, SumOutputs_6_51_port, SumOutputs_6_50_port, 
      SumOutputs_6_49_port, SumOutputs_6_48_port, SumOutputs_6_47_port, 
      SumOutputs_6_46_port, SumOutputs_6_45_port, SumOutputs_6_44_port, 
      SumOutputs_6_43_port, SumOutputs_6_42_port, SumOutputs_6_41_port, 
      SumOutputs_6_40_port, SumOutputs_6_39_port, SumOutputs_6_38_port, 
      SumOutputs_6_37_port, SumOutputs_6_36_port, SumOutputs_6_35_port, 
      SumOutputs_6_34_port, SumOutputs_6_33_port, SumOutputs_6_32_port, 
      SumOutputs_6_31_port, SumOutputs_6_30_port, SumOutputs_6_29_port, 
      SumOutputs_6_28_port, SumOutputs_6_27_port, SumOutputs_6_26_port, 
      SumOutputs_6_25_port, SumOutputs_6_24_port, SumOutputs_6_23_port, 
      SumOutputs_6_22_port, SumOutputs_6_21_port, SumOutputs_6_20_port, 
      SumOutputs_6_19_port, SumOutputs_6_18_port, SumOutputs_6_17_port, 
      SumOutputs_6_16_port, SumOutputs_6_15_port, SumOutputs_6_14_port, 
      SumOutputs_6_13_port, SumOutputs_6_12_port, SumOutputs_6_11_port, 
      SumOutputs_6_10_port, SumOutputs_6_9_port, SumOutputs_6_8_port, 
      SumOutputs_6_7_port, SumOutputs_6_6_port, SumOutputs_6_5_port, 
      SumOutputs_6_4_port, SumOutputs_6_3_port, SumOutputs_6_2_port, 
      SumOutputs_6_1_port, SumOutputs_6_0_port, SumOutputs_5_63_port, 
      SumOutputs_5_62_port, SumOutputs_5_61_port, SumOutputs_5_60_port, 
      SumOutputs_5_59_port, SumOutputs_5_58_port, SumOutputs_5_57_port, 
      SumOutputs_5_56_port, SumOutputs_5_55_port, SumOutputs_5_54_port, 
      SumOutputs_5_53_port, SumOutputs_5_52_port, SumOutputs_5_51_port, 
      SumOutputs_5_50_port, SumOutputs_5_49_port, SumOutputs_5_48_port, 
      SumOutputs_5_47_port, SumOutputs_5_46_port, SumOutputs_5_45_port, 
      SumOutputs_5_44_port, SumOutputs_5_43_port, SumOutputs_5_42_port, 
      SumOutputs_5_41_port, SumOutputs_5_40_port, SumOutputs_5_39_port, 
      SumOutputs_5_38_port, SumOutputs_5_37_port, SumOutputs_5_36_port, 
      SumOutputs_5_35_port, SumOutputs_5_34_port, SumOutputs_5_33_port, 
      SumOutputs_5_32_port, SumOutputs_5_31_port, SumOutputs_5_30_port, 
      SumOutputs_5_29_port, SumOutputs_5_28_port, SumOutputs_5_27_port, 
      SumOutputs_5_26_port, SumOutputs_5_25_port, SumOutputs_5_24_port, 
      SumOutputs_5_23_port, SumOutputs_5_22_port, SumOutputs_5_21_port, 
      SumOutputs_5_20_port, SumOutputs_5_19_port, SumOutputs_5_18_port, 
      SumOutputs_5_17_port, SumOutputs_5_16_port, SumOutputs_5_15_port, 
      SumOutputs_5_14_port, SumOutputs_5_13_port, SumOutputs_5_12_port, 
      SumOutputs_5_11_port, SumOutputs_5_10_port, SumOutputs_5_9_port, 
      SumOutputs_5_8_port, SumOutputs_5_7_port, SumOutputs_5_6_port, 
      SumOutputs_5_5_port, SumOutputs_5_4_port, SumOutputs_5_3_port, 
      SumOutputs_5_2_port, SumOutputs_5_1_port, SumOutputs_5_0_port, 
      SumOutputs_4_63_port, SumOutputs_4_62_port, SumOutputs_4_61_port, 
      SumOutputs_4_60_port, SumOutputs_4_59_port, SumOutputs_4_58_port, 
      SumOutputs_4_57_port, SumOutputs_4_56_port, SumOutputs_4_55_port, 
      SumOutputs_4_54_port, SumOutputs_4_53_port, SumOutputs_4_52_port, 
      SumOutputs_4_51_port, SumOutputs_4_50_port, SumOutputs_4_49_port, 
      SumOutputs_4_48_port, SumOutputs_4_47_port, SumOutputs_4_46_port, 
      SumOutputs_4_45_port, SumOutputs_4_44_port, SumOutputs_4_43_port, 
      SumOutputs_4_42_port, SumOutputs_4_41_port, SumOutputs_4_40_port, 
      SumOutputs_4_39_port, SumOutputs_4_38_port, SumOutputs_4_37_port, 
      SumOutputs_4_36_port, SumOutputs_4_35_port, SumOutputs_4_34_port, 
      SumOutputs_4_33_port, SumOutputs_4_32_port, SumOutputs_4_31_port, 
      SumOutputs_4_30_port, SumOutputs_4_29_port, SumOutputs_4_28_port, 
      SumOutputs_4_27_port, SumOutputs_4_26_port, SumOutputs_4_25_port, 
      SumOutputs_4_24_port, SumOutputs_4_23_port, SumOutputs_4_22_port, 
      SumOutputs_4_21_port, SumOutputs_4_20_port, SumOutputs_4_19_port, 
      SumOutputs_4_18_port, SumOutputs_4_17_port, SumOutputs_4_16_port, 
      SumOutputs_4_15_port, SumOutputs_4_14_port, SumOutputs_4_13_port, 
      SumOutputs_4_12_port, SumOutputs_4_11_port, SumOutputs_4_10_port, 
      SumOutputs_4_9_port, SumOutputs_4_8_port, SumOutputs_4_7_port, 
      SumOutputs_4_6_port, SumOutputs_4_5_port, SumOutputs_4_4_port, 
      SumOutputs_4_3_port, SumOutputs_4_2_port, SumOutputs_4_1_port, 
      SumOutputs_4_0_port, SumOutputs_3_63_port, SumOutputs_3_62_port, 
      SumOutputs_3_61_port, SumOutputs_3_60_port, SumOutputs_3_59_port, 
      SumOutputs_3_58_port, SumOutputs_3_57_port, SumOutputs_3_56_port, 
      SumOutputs_3_55_port, SumOutputs_3_54_port, SumOutputs_3_53_port, 
      SumOutputs_3_52_port, SumOutputs_3_51_port, SumOutputs_3_50_port, 
      SumOutputs_3_49_port, SumOutputs_3_48_port, SumOutputs_3_47_port, 
      SumOutputs_3_46_port, SumOutputs_3_45_port, SumOutputs_3_44_port, 
      SumOutputs_3_43_port, SumOutputs_3_42_port, SumOutputs_3_41_port, 
      SumOutputs_3_40_port, SumOutputs_3_39_port, SumOutputs_3_38_port, 
      SumOutputs_3_37_port, SumOutputs_3_36_port, SumOutputs_3_35_port, 
      SumOutputs_3_34_port, SumOutputs_3_33_port, SumOutputs_3_32_port, 
      SumOutputs_3_31_port, SumOutputs_3_30_port, SumOutputs_3_29_port, 
      SumOutputs_3_28_port, SumOutputs_3_27_port, SumOutputs_3_26_port, 
      SumOutputs_3_25_port, SumOutputs_3_24_port, SumOutputs_3_23_port, 
      SumOutputs_3_22_port, SumOutputs_3_21_port, SumOutputs_3_20_port, 
      SumOutputs_3_19_port, SumOutputs_3_18_port, SumOutputs_3_17_port, 
      SumOutputs_3_16_port, SumOutputs_3_15_port, SumOutputs_3_14_port, 
      SumOutputs_3_13_port, SumOutputs_3_12_port, SumOutputs_3_11_port, 
      SumOutputs_3_10_port, SumOutputs_3_9_port, SumOutputs_3_8_port, 
      SumOutputs_3_7_port, SumOutputs_3_6_port, SumOutputs_3_5_port, 
      SumOutputs_3_4_port, SumOutputs_3_3_port, SumOutputs_3_2_port, 
      SumOutputs_3_1_port, SumOutputs_3_0_port, SumOutputs_2_63_port, 
      SumOutputs_2_62_port, SumOutputs_2_61_port, SumOutputs_2_60_port, 
      SumOutputs_2_59_port, SumOutputs_2_58_port, SumOutputs_2_57_port, 
      SumOutputs_2_56_port, SumOutputs_2_55_port, SumOutputs_2_54_port, 
      SumOutputs_2_53_port, SumOutputs_2_52_port, SumOutputs_2_51_port, 
      SumOutputs_2_50_port, SumOutputs_2_49_port, SumOutputs_2_48_port, 
      SumOutputs_2_47_port, SumOutputs_2_46_port, SumOutputs_2_45_port, 
      SumOutputs_2_44_port, SumOutputs_2_43_port, SumOutputs_2_42_port, 
      SumOutputs_2_41_port, SumOutputs_2_40_port, SumOutputs_2_39_port, 
      SumOutputs_2_38_port, SumOutputs_2_37_port, SumOutputs_2_36_port, 
      SumOutputs_2_35_port, SumOutputs_2_34_port, SumOutputs_2_33_port, 
      SumOutputs_2_32_port, SumOutputs_2_31_port, SumOutputs_2_30_port, 
      SumOutputs_2_29_port, SumOutputs_2_28_port, SumOutputs_2_27_port, 
      SumOutputs_2_26_port, SumOutputs_2_25_port, SumOutputs_2_24_port, 
      SumOutputs_2_23_port, SumOutputs_2_22_port, SumOutputs_2_21_port, 
      SumOutputs_2_20_port, SumOutputs_2_19_port, SumOutputs_2_18_port, 
      SumOutputs_2_17_port, SumOutputs_2_16_port, SumOutputs_2_15_port, 
      SumOutputs_2_14_port, SumOutputs_2_13_port, SumOutputs_2_12_port, 
      SumOutputs_2_11_port, SumOutputs_2_10_port, SumOutputs_2_9_port, 
      SumOutputs_2_8_port, SumOutputs_2_7_port, SumOutputs_2_6_port, 
      SumOutputs_2_5_port, SumOutputs_2_4_port, SumOutputs_2_3_port, 
      SumOutputs_2_2_port, SumOutputs_2_1_port, SumOutputs_2_0_port, 
      SumOutputs_1_63_port, SumOutputs_1_62_port, SumOutputs_1_61_port, 
      SumOutputs_1_60_port, SumOutputs_1_59_port, SumOutputs_1_58_port, 
      SumOutputs_1_57_port, SumOutputs_1_56_port, SumOutputs_1_55_port, 
      SumOutputs_1_54_port, SumOutputs_1_53_port, SumOutputs_1_52_port, 
      SumOutputs_1_51_port, SumOutputs_1_50_port, SumOutputs_1_49_port, 
      SumOutputs_1_48_port, SumOutputs_1_47_port, SumOutputs_1_46_port, 
      SumOutputs_1_45_port, SumOutputs_1_44_port, SumOutputs_1_43_port, 
      SumOutputs_1_42_port, SumOutputs_1_41_port, SumOutputs_1_40_port, 
      SumOutputs_1_39_port, SumOutputs_1_38_port, SumOutputs_1_37_port, 
      SumOutputs_1_36_port, SumOutputs_1_35_port, SumOutputs_1_34_port, 
      SumOutputs_1_33_port, SumOutputs_1_32_port, SumOutputs_1_31_port, 
      SumOutputs_1_30_port, SumOutputs_1_29_port, SumOutputs_1_28_port, 
      SumOutputs_1_27_port, SumOutputs_1_26_port, SumOutputs_1_25_port, 
      SumOutputs_1_24_port, SumOutputs_1_23_port, SumOutputs_1_22_port, 
      SumOutputs_1_21_port, SumOutputs_1_20_port, SumOutputs_1_19_port, 
      SumOutputs_1_18_port, SumOutputs_1_17_port, SumOutputs_1_16_port, 
      SumOutputs_1_15_port, SumOutputs_1_14_port, SumOutputs_1_13_port, 
      SumOutputs_1_12_port, SumOutputs_1_11_port, SumOutputs_1_10_port, 
      SumOutputs_1_9_port, SumOutputs_1_8_port, SumOutputs_1_7_port, 
      SumOutputs_1_6_port, SumOutputs_1_5_port, SumOutputs_1_4_port, 
      SumOutputs_1_3_port, SumOutputs_1_2_port, SumOutputs_1_1_port, 
      SumOutputs_1_0_port, SumOutputs_0_63_port, SumOutputs_0_62_port, 
      SumOutputs_0_61_port, SumOutputs_0_60_port, SumOutputs_0_59_port, 
      SumOutputs_0_58_port, SumOutputs_0_57_port, SumOutputs_0_56_port, 
      SumOutputs_0_55_port, SumOutputs_0_54_port, SumOutputs_0_53_port, 
      SumOutputs_0_52_port, SumOutputs_0_51_port, SumOutputs_0_50_port, 
      SumOutputs_0_49_port, SumOutputs_0_48_port, SumOutputs_0_47_port, 
      SumOutputs_0_46_port, SumOutputs_0_45_port, SumOutputs_0_44_port, 
      SumOutputs_0_43_port, SumOutputs_0_42_port, SumOutputs_0_41_port, 
      SumOutputs_0_40_port, SumOutputs_0_39_port, SumOutputs_0_38_port, 
      SumOutputs_0_37_port, SumOutputs_0_36_port, SumOutputs_0_35_port, 
      SumOutputs_0_34_port, SumOutputs_0_33_port, SumOutputs_0_32_port, 
      SumOutputs_0_31_port, SumOutputs_0_30_port, SumOutputs_0_29_port, 
      SumOutputs_0_28_port, SumOutputs_0_27_port, SumOutputs_0_26_port, 
      SumOutputs_0_25_port, SumOutputs_0_24_port, SumOutputs_0_23_port, 
      SumOutputs_0_22_port, SumOutputs_0_21_port, SumOutputs_0_20_port, 
      SumOutputs_0_19_port, SumOutputs_0_18_port, SumOutputs_0_17_port, 
      SumOutputs_0_16_port, SumOutputs_0_15_port, SumOutputs_0_14_port, 
      SumOutputs_0_13_port, SumOutputs_0_12_port, SumOutputs_0_11_port, 
      SumOutputs_0_10_port, SumOutputs_0_9_port, SumOutputs_0_8_port, 
      SumOutputs_0_7_port, SumOutputs_0_6_port, SumOutputs_0_5_port, 
      SumOutputs_0_4_port, SumOutputs_0_3_port, SumOutputs_0_2_port, 
      SumOutputs_0_1_port, SumOutputs_0_0_port, SumOutputs_13_63_port, 
      SumOutputs_13_62_port, SumOutputs_13_61_port, SumOutputs_13_60_port, 
      SumOutputs_13_59_port, SumOutputs_13_58_port, SumOutputs_13_57_port, 
      SumOutputs_13_56_port, SumOutputs_13_55_port, SumOutputs_13_54_port, 
      SumOutputs_13_53_port, SumOutputs_13_52_port, SumOutputs_13_51_port, 
      SumOutputs_13_50_port, SumOutputs_13_49_port, SumOutputs_13_48_port, 
      SumOutputs_13_47_port, SumOutputs_13_46_port, SumOutputs_13_45_port, 
      SumOutputs_13_44_port, SumOutputs_13_43_port, SumOutputs_13_42_port, 
      SumOutputs_13_41_port, SumOutputs_13_40_port, SumOutputs_13_39_port, 
      SumOutputs_13_38_port, SumOutputs_13_37_port, SumOutputs_13_36_port, 
      SumOutputs_13_35_port, SumOutputs_13_34_port, SumOutputs_13_33_port, 
      SumOutputs_13_32_port, SumOutputs_13_31_port, SumOutputs_13_30_port, 
      SumOutputs_13_29_port, SumOutputs_13_28_port, SumOutputs_13_27_port, 
      SumOutputs_13_26_port, SumOutputs_13_25_port, SumOutputs_13_24_port, 
      SumOutputs_13_23_port, SumOutputs_13_22_port, SumOutputs_13_21_port, 
      SumOutputs_13_20_port, SumOutputs_13_19_port, SumOutputs_13_18_port, 
      SumOutputs_13_17_port, SumOutputs_13_16_port, SumOutputs_13_15_port, 
      SumOutputs_13_14_port, SumOutputs_13_13_port, SumOutputs_13_12_port, 
      SumOutputs_13_11_port, SumOutputs_13_10_port, SumOutputs_13_9_port, 
      SumOutputs_13_8_port, SumOutputs_13_7_port, SumOutputs_13_6_port, 
      SumOutputs_13_5_port, SumOutputs_13_4_port, SumOutputs_13_3_port, 
      SumOutputs_13_2_port, SumOutputs_13_1_port, SumOutputs_13_0_port, 
      SumOutputs_12_63_port, SumOutputs_12_62_port, SumOutputs_12_61_port, 
      SumOutputs_12_60_port, SumOutputs_12_59_port, SumOutputs_12_58_port, 
      SumOutputs_12_57_port, SumOutputs_12_56_port, SumOutputs_12_55_port, 
      SumOutputs_12_54_port, SumOutputs_12_53_port, SumOutputs_12_52_port, 
      SumOutputs_12_51_port, SumOutputs_12_50_port, SumOutputs_12_49_port, 
      SumOutputs_12_48_port, SumOutputs_12_47_port, SumOutputs_12_46_port, 
      SumOutputs_12_45_port, SumOutputs_12_44_port, SumOutputs_12_43_port, 
      SumOutputs_12_42_port, SumOutputs_12_41_port, SumOutputs_12_40_port, 
      SumOutputs_12_39_port, SumOutputs_12_38_port, SumOutputs_12_37_port, 
      SumOutputs_12_36_port, SumOutputs_12_35_port, SumOutputs_12_34_port, 
      SumOutputs_12_33_port, SumOutputs_12_32_port, SumOutputs_12_31_port, 
      SumOutputs_12_30_port, SumOutputs_12_29_port, SumOutputs_12_28_port, 
      SumOutputs_12_27_port, SumOutputs_12_26_port, SumOutputs_12_25_port, 
      SumOutputs_12_24_port, SumOutputs_12_23_port, SumOutputs_12_22_port, 
      SumOutputs_12_21_port, SumOutputs_12_20_port, SumOutputs_12_19_port, 
      SumOutputs_12_18_port, SumOutputs_12_17_port, SumOutputs_12_16_port, 
      SumOutputs_12_15_port, SumOutputs_12_14_port, SumOutputs_12_13_port, 
      SumOutputs_12_12_port, SumOutputs_12_11_port, SumOutputs_12_10_port, 
      SumOutputs_12_9_port, SumOutputs_12_8_port, SumOutputs_12_7_port, 
      SumOutputs_12_6_port, SumOutputs_12_5_port, SumOutputs_12_4_port, 
      SumOutputs_12_3_port, SumOutputs_12_2_port, SumOutputs_12_1_port, 
      SumOutputs_12_0_port, SumOutputs_11_63_port, SumOutputs_11_62_port, 
      SumOutputs_11_61_port, SumOutputs_11_60_port, SumOutputs_11_59_port, 
      SumOutputs_11_58_port, SumOutputs_11_57_port, SumOutputs_11_56_port, 
      SumOutputs_11_55_port, SumOutputs_11_54_port, SumOutputs_11_53_port, 
      SumOutputs_11_52_port, SumOutputs_11_51_port, SumOutputs_11_50_port, 
      SumOutputs_11_49_port, SumOutputs_11_48_port, SumOutputs_11_47_port, 
      SumOutputs_11_46_port, SumOutputs_11_45_port, SumOutputs_11_44_port, 
      SumOutputs_11_43_port, SumOutputs_11_42_port, SumOutputs_11_41_port, 
      SumOutputs_11_40_port, SumOutputs_11_39_port, SumOutputs_11_38_port, 
      SumOutputs_11_37_port, SumOutputs_11_36_port, SumOutputs_11_35_port, 
      SumOutputs_11_34_port, SumOutputs_11_33_port, SumOutputs_11_32_port, 
      SumOutputs_11_31_port, SumOutputs_11_30_port, SumOutputs_11_29_port, 
      SumOutputs_11_28_port, SumOutputs_11_27_port, SumOutputs_11_26_port, 
      SumOutputs_11_25_port, SumOutputs_11_24_port, SumOutputs_11_23_port, 
      SumOutputs_11_22_port, SumOutputs_11_21_port, SumOutputs_11_20_port, 
      SumOutputs_11_19_port, SumOutputs_11_18_port, SumOutputs_11_17_port, 
      SumOutputs_11_16_port, SumOutputs_11_15_port, SumOutputs_11_14_port, 
      SumOutputs_11_13_port, SumOutputs_11_12_port, SumOutputs_11_11_port, 
      SumOutputs_11_10_port, SumOutputs_11_9_port, SumOutputs_11_8_port, 
      SumOutputs_11_7_port, SumOutputs_11_6_port, SumOutputs_11_5_port, 
      SumOutputs_11_4_port, SumOutputs_11_3_port, SumOutputs_11_2_port, 
      SumOutputs_11_1_port, SumOutputs_11_0_port, SumOutputs_10_63_port, 
      SumOutputs_10_62_port, SumOutputs_10_61_port, SumOutputs_10_60_port, 
      SumOutputs_10_59_port, SumOutputs_10_58_port, SumOutputs_10_57_port, 
      SumOutputs_10_56_port, SumOutputs_10_55_port, SumOutputs_10_54_port, 
      SumOutputs_10_53_port, SumOutputs_10_52_port, SumOutputs_10_51_port, 
      SumOutputs_10_50_port, SumOutputs_10_49_port, SumOutputs_10_48_port, 
      SumOutputs_10_47_port, SumOutputs_10_46_port, SumOutputs_10_45_port, 
      SumOutputs_10_44_port, SumOutputs_10_43_port, SumOutputs_10_42_port, 
      SumOutputs_10_41_port, SumOutputs_10_40_port, SumOutputs_10_39_port, 
      SumOutputs_10_38_port, SumOutputs_10_37_port, SumOutputs_10_36_port, 
      SumOutputs_10_35_port, SumOutputs_10_34_port, SumOutputs_10_33_port, 
      SumOutputs_10_32_port, SumOutputs_10_31_port, SumOutputs_10_30_port, 
      SumOutputs_10_29_port, SumOutputs_10_28_port, SumOutputs_10_27_port, 
      SumOutputs_10_26_port, SumOutputs_10_25_port, SumOutputs_10_24_port, 
      SumOutputs_10_23_port, SumOutputs_10_22_port, SumOutputs_10_21_port, 
      SumOutputs_10_20_port, SumOutputs_10_19_port, SumOutputs_10_18_port, 
      SumOutputs_10_17_port, SumOutputs_10_16_port, SumOutputs_10_15_port, 
      SumOutputs_10_14_port, SumOutputs_10_13_port, SumOutputs_10_12_port, 
      SumOutputs_10_11_port, SumOutputs_10_10_port, SumOutputs_10_9_port, 
      SumOutputs_10_8_port, SumOutputs_10_7_port, SumOutputs_10_6_port, 
      SumOutputs_10_5_port, SumOutputs_10_4_port, SumOutputs_10_3_port, 
      SumOutputs_10_2_port, SumOutputs_10_1_port, SumOutputs_10_0_port, 
      SumOutputs_9_63_port, SumOutputs_9_62_port, SumOutputs_9_61_port, 
      SumOutputs_9_60_port, SumOutputs_9_59_port, SumOutputs_9_58_port, 
      SumOutputs_9_57_port, SumOutputs_9_56_port, SumOutputs_9_55_port, 
      SumOutputs_9_54_port, SumOutputs_9_53_port, SumOutputs_9_52_port, 
      SumOutputs_9_51_port, SumOutputs_9_50_port, SumOutputs_9_49_port, 
      SumOutputs_9_48_port, SumOutputs_9_47_port, SumOutputs_9_46_port, 
      SumOutputs_9_45_port, SumOutputs_9_44_port, SumOutputs_9_43_port, 
      SumOutputs_9_42_port, SumOutputs_9_41_port, SumOutputs_9_40_port, 
      SumOutputs_9_39_port, SumOutputs_9_38_port, SumOutputs_9_37_port, 
      SumOutputs_9_36_port, SumOutputs_9_35_port, SumOutputs_9_34_port, 
      SumOutputs_9_33_port, SumOutputs_9_32_port, SumOutputs_9_31_port, 
      SumOutputs_9_30_port, SumOutputs_9_29_port, SumOutputs_9_28_port, 
      SumOutputs_9_27_port, SumOutputs_9_26_port, SumOutputs_9_25_port, 
      SumOutputs_9_24_port, SumOutputs_9_23_port, SumOutputs_9_22_port, 
      SumOutputs_9_21_port, SumOutputs_9_20_port, SumOutputs_9_19_port, 
      SumOutputs_9_18_port, SumOutputs_9_17_port, SumOutputs_9_16_port, 
      SumOutputs_9_15_port, SumOutputs_9_14_port, SumOutputs_9_13_port, 
      SumOutputs_9_12_port, SumOutputs_9_11_port, SumOutputs_9_10_port, 
      SumOutputs_9_9_port, SumOutputs_9_8_port, SumOutputs_9_7_port, 
      SumOutputs_9_6_port, SumOutputs_9_5_port, SumOutputs_9_4_port, 
      SumOutputs_9_3_port, SumOutputs_9_2_port, SumOutputs_9_1_port, 
      SumOutputs_9_0_port, SumOutputs_8_63_port, SumOutputs_8_62_port, 
      SumOutputs_8_61_port, SumOutputs_8_60_port, SumOutputs_8_59_port, 
      SumOutputs_8_58_port, SumOutputs_8_57_port, SumOutputs_8_56_port, 
      SumOutputs_8_55_port, SumOutputs_8_54_port, SumOutputs_8_53_port, 
      SumOutputs_8_52_port, SumOutputs_8_51_port, SumOutputs_8_50_port, 
      SumOutputs_8_49_port, SumOutputs_8_48_port, SumOutputs_8_47_port, 
      SumOutputs_8_46_port, SumOutputs_8_45_port, SumOutputs_8_44_port, 
      SumOutputs_8_43_port, SumOutputs_8_42_port, SumOutputs_8_41_port, 
      SumOutputs_8_40_port, SumOutputs_8_39_port, SumOutputs_8_38_port, 
      SumOutputs_8_37_port, SumOutputs_8_36_port, SumOutputs_8_35_port, 
      SumOutputs_8_34_port, SumOutputs_8_33_port, SumOutputs_8_32_port, 
      SumOutputs_8_31_port, SumOutputs_8_30_port, SumOutputs_8_29_port, 
      SumOutputs_8_28_port, SumOutputs_8_27_port, SumOutputs_8_26_port, 
      SumOutputs_8_25_port, SumOutputs_8_24_port, SumOutputs_8_23_port, 
      SumOutputs_8_22_port, SumOutputs_8_21_port, SumOutputs_8_20_port, 
      SumOutputs_8_19_port, SumOutputs_8_18_port, SumOutputs_8_17_port, 
      SumOutputs_8_16_port, SumOutputs_8_15_port, SumOutputs_8_14_port, 
      SumOutputs_8_13_port, SumOutputs_8_12_port, SumOutputs_8_11_port, 
      SumOutputs_8_10_port, SumOutputs_8_9_port, SumOutputs_8_8_port, 
      SumOutputs_8_7_port, SumOutputs_8_6_port, SumOutputs_8_5_port, 
      SumOutputs_8_4_port, SumOutputs_8_3_port, SumOutputs_8_2_port, 
      SumOutputs_8_1_port, SumOutputs_8_0_port, n9, n10, n11, n12, n13, n14, 
      n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29
      , n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, 
      n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58
      , n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, 
      n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87
      , n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
      n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, 
      n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, 
      n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, 
      n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, 
      n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, 
      n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, 
      n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, 
      n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, 
      n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, 
      n210, n211, n212, n213, n214, n215, n_1000, n_1001, n_1002, n_1003, 
      n_1004, n_1005, n_1006, n_1007, n_1008, n_1009, n_1010, n_1011, n_1012, 
      n_1013, n_1014, n_1015, n_1016, n_1017, n_1018, n_1019, n_1020, n_1021, 
      n_1022, n_1023, n_1024, n_1025, n_1026, n_1027, n_1028, n_1029, n_1030, 
      n_1031, n_1032, n_1033, n_1034, n_1035, n_1036, n_1037, n_1038, n_1039, 
      n_1040, n_1041, n_1042, n_1043, n_1044, n_1045, n_1046, n_1047, n_1048, 
      n_1049, n_1050, n_1051, n_1052, n_1053, n_1054, n_1055, n_1056, n_1057, 
      n_1058, n_1059, n_1060, n_1061, n_1062, n_1063, n_1064, n_1065, n_1066, 
      n_1067, n_1068, n_1069, n_1070, n_1071, n_1072, n_1073, n_1074, n_1075, 
      n_1076, n_1077, n_1078, n_1079, n_1080, n_1081, n_1082, n_1083, n_1084, 
      n_1085, n_1086, n_1087, n_1088, n_1089, n_1090, n_1091, n_1092, n_1093, 
      n_1094, n_1095, n_1096, n_1097, n_1098, n_1099, n_1100, n_1101, n_1102, 
      n_1103, n_1104, n_1105, n_1106, n_1107, n_1108, n_1109, n_1110, n_1111, 
      n_1112, n_1113, n_1114, n_1115, n_1116, n_1117, n_1118, n_1119, n_1120, 
      n_1121, n_1122, n_1123, n_1124, n_1125, n_1126, n_1127, n_1128, n_1129, 
      n_1130, n_1131, n_1132, n_1133, n_1134, n_1135, n_1136, n_1137, n_1138, 
      n_1139, n_1140, n_1141 : std_logic;

begin
   
   inverterI_0 : IV_0 port map( A => A(0), Y => A_complement_0_port);
   inverterI_1 : IV_63 port map( A => A(1), Y => A_complement_1_port);
   inverterI_2 : IV_62 port map( A => A(2), Y => A_complement_2_port);
   inverterI_3 : IV_61 port map( A => A(3), Y => A_complement_3_port);
   inverterI_4 : IV_60 port map( A => A(4), Y => A_complement_4_port);
   inverterI_5 : IV_59 port map( A => A(5), Y => A_complement_5_port);
   inverterI_6 : IV_58 port map( A => A(6), Y => A_complement_6_port);
   inverterI_7 : IV_57 port map( A => A(7), Y => A_complement_7_port);
   inverterI_8 : IV_56 port map( A => A(8), Y => A_complement_8_port);
   inverterI_9 : IV_55 port map( A => A(9), Y => A_complement_9_port);
   inverterI_10 : IV_54 port map( A => A(10), Y => A_complement_10_port);
   inverterI_11 : IV_53 port map( A => A(11), Y => A_complement_11_port);
   inverterI_12 : IV_52 port map( A => A(12), Y => A_complement_12_port);
   inverterI_13 : IV_51 port map( A => A(13), Y => A_complement_13_port);
   inverterI_14 : IV_50 port map( A => A(14), Y => A_complement_14_port);
   inverterI_15 : IV_49 port map( A => A(15), Y => A_complement_15_port);
   inverterI_16 : IV_48 port map( A => A(16), Y => A_complement_16_port);
   inverterI_17 : IV_47 port map( A => A(17), Y => A_complement_17_port);
   inverterI_18 : IV_46 port map( A => A(18), Y => A_complement_18_port);
   inverterI_19 : IV_45 port map( A => A(19), Y => A_complement_19_port);
   inverterI_20 : IV_44 port map( A => A(20), Y => A_complement_20_port);
   inverterI_21 : IV_43 port map( A => A(21), Y => A_complement_21_port);
   inverterI_22 : IV_42 port map( A => A(22), Y => A_complement_22_port);
   inverterI_23 : IV_41 port map( A => A(23), Y => A_complement_23_port);
   inverterI_24 : IV_40 port map( A => A(24), Y => A_complement_24_port);
   inverterI_25 : IV_39 port map( A => A(25), Y => A_complement_25_port);
   inverterI_26 : IV_38 port map( A => A(26), Y => A_complement_26_port);
   inverterI_27 : IV_37 port map( A => A(27), Y => A_complement_27_port);
   inverterI_28 : IV_36 port map( A => A(28), Y => A_complement_28_port);
   inverterI_29 : IV_35 port map( A => A(29), Y => A_complement_29_port);
   inverterI_30 : IV_34 port map( A => A(30), Y => A_complement_30_port);
   inverterI_31 : IV_33 port map( A => A(31), Y => A_complement_31_port);
   inverterI_32 : IV_32 port map( A => A(31), Y => A_complement_32_port);
   inverterI_33 : IV_31 port map( A => A(31), Y => A_complement_33_port);
   inverterI_34 : IV_30 port map( A => A(31), Y => A_complement_34_port);
   inverterI_35 : IV_29 port map( A => A(31), Y => A_complement_35_port);
   inverterI_36 : IV_28 port map( A => A(31), Y => A_complement_36_port);
   inverterI_37 : IV_27 port map( A => A(31), Y => A_complement_37_port);
   inverterI_38 : IV_26 port map( A => A(31), Y => A_complement_38_port);
   inverterI_39 : IV_25 port map( A => A(31), Y => A_complement_39_port);
   inverterI_40 : IV_24 port map( A => A(31), Y => A_complement_40_port);
   inverterI_41 : IV_23 port map( A => A(31), Y => A_complement_41_port);
   inverterI_42 : IV_22 port map( A => A(31), Y => A_complement_42_port);
   inverterI_43 : IV_21 port map( A => A(31), Y => A_complement_43_port);
   inverterI_44 : IV_20 port map( A => A(31), Y => A_complement_44_port);
   inverterI_45 : IV_19 port map( A => A(31), Y => A_complement_45_port);
   inverterI_46 : IV_18 port map( A => A(31), Y => A_complement_46_port);
   inverterI_47 : IV_17 port map( A => A(31), Y => A_complement_47_port);
   inverterI_48 : IV_16 port map( A => A(31), Y => A_complement_48_port);
   inverterI_49 : IV_15 port map( A => A(31), Y => A_complement_49_port);
   inverterI_50 : IV_14 port map( A => A(31), Y => A_complement_50_port);
   inverterI_51 : IV_13 port map( A => A(31), Y => A_complement_51_port);
   inverterI_52 : IV_12 port map( A => A(31), Y => A_complement_52_port);
   inverterI_53 : IV_11 port map( A => A(31), Y => A_complement_53_port);
   inverterI_54 : IV_10 port map( A => A(31), Y => A_complement_54_port);
   inverterI_55 : IV_9 port map( A => A(31), Y => A_complement_55_port);
   inverterI_56 : IV_8 port map( A => A(31), Y => A_complement_56_port);
   inverterI_57 : IV_7 port map( A => A(31), Y => A_complement_57_port);
   inverterI_58 : IV_6 port map( A => A(31), Y => A_complement_58_port);
   inverterI_59 : IV_5 port map( A => A(31), Y => A_complement_59_port);
   inverterI_60 : IV_4 port map( A => A(31), Y => A_complement_60_port);
   inverterI_61 : IV_3 port map( A => A(31), Y => A_complement_61_port);
   inverterI_62 : IV_2 port map( A => A(31), Y => A_complement_62_port);
   inverterI_63 : IV_1 port map( A => A(31), Y => A_complement_63_port);
   FinilizingNegativeSignal : RCA_NbitRca64_0 port map( A(63) => 
                           A_complement_63_port, A(62) => A_complement_62_port,
                           A(61) => A_complement_61_port, A(60) => 
                           A_complement_60_port, A(59) => A_complement_59_port,
                           A(58) => A_complement_58_port, A(57) => 
                           A_complement_57_port, A(56) => A_complement_56_port,
                           A(55) => A_complement_55_port, A(54) => 
                           A_complement_54_port, A(53) => A_complement_53_port,
                           A(52) => A_complement_52_port, A(51) => 
                           A_complement_51_port, A(50) => A_complement_50_port,
                           A(49) => A_complement_49_port, A(48) => 
                           A_complement_48_port, A(47) => A_complement_47_port,
                           A(46) => A_complement_46_port, A(45) => 
                           A_complement_45_port, A(44) => A_complement_44_port,
                           A(43) => A_complement_43_port, A(42) => 
                           A_complement_42_port, A(41) => A_complement_41_port,
                           A(40) => A_complement_40_port, A(39) => 
                           A_complement_39_port, A(38) => A_complement_38_port,
                           A(37) => A_complement_37_port, A(36) => 
                           A_complement_36_port, A(35) => A_complement_35_port,
                           A(34) => A_complement_34_port, A(33) => 
                           A_complement_33_port, A(32) => A_complement_32_port,
                           A(31) => A_complement_31_port, A(30) => 
                           A_complement_30_port, A(29) => A_complement_29_port,
                           A(28) => A_complement_28_port, A(27) => 
                           A_complement_27_port, A(26) => A_complement_26_port,
                           A(25) => A_complement_25_port, A(24) => 
                           A_complement_24_port, A(23) => A_complement_23_port,
                           A(22) => A_complement_22_port, A(21) => 
                           A_complement_21_port, A(20) => A_complement_20_port,
                           A(19) => A_complement_19_port, A(18) => 
                           A_complement_18_port, A(17) => A_complement_17_port,
                           A(16) => A_complement_16_port, A(15) => 
                           A_complement_15_port, A(14) => A_complement_14_port,
                           A(13) => A_complement_13_port, A(12) => 
                           A_complement_12_port, A(11) => A_complement_11_port,
                           A(10) => A_complement_10_port, A(9) => 
                           A_complement_9_port, A(8) => A_complement_8_port, 
                           A(7) => A_complement_7_port, A(6) => 
                           A_complement_6_port, A(5) => A_complement_5_port, 
                           A(4) => A_complement_4_port, A(3) => 
                           A_complement_3_port, A(2) => A_complement_2_port, 
                           A(1) => A_complement_1_port, A(0) => 
                           A_complement_0_port, B(63) => X_Logic0_port, B(62) 
                           => X_Logic0_port, B(61) => X_Logic0_port, B(60) => 
                           X_Logic0_port, B(59) => X_Logic0_port, B(58) => 
                           X_Logic0_port, B(57) => X_Logic0_port, B(56) => 
                           X_Logic0_port, B(55) => X_Logic0_port, B(54) => 
                           X_Logic0_port, B(53) => X_Logic0_port, B(52) => 
                           X_Logic0_port, B(51) => X_Logic0_port, B(50) => 
                           X_Logic0_port, B(49) => X_Logic0_port, B(48) => 
                           X_Logic0_port, B(47) => X_Logic0_port, B(46) => 
                           X_Logic0_port, B(45) => X_Logic0_port, B(44) => 
                           X_Logic0_port, B(43) => X_Logic0_port, B(42) => 
                           X_Logic0_port, B(41) => X_Logic0_port, B(40) => 
                           X_Logic0_port, B(39) => X_Logic0_port, B(38) => 
                           X_Logic0_port, B(37) => X_Logic0_port, B(36) => 
                           X_Logic0_port, B(35) => X_Logic0_port, B(34) => 
                           X_Logic0_port, B(33) => X_Logic0_port, B(32) => 
                           X_Logic0_port, B(31) => X_Logic0_port, B(30) => 
                           X_Logic0_port, B(29) => X_Logic0_port, B(28) => 
                           X_Logic0_port, B(27) => X_Logic0_port, B(26) => 
                           X_Logic0_port, B(25) => X_Logic0_port, B(24) => 
                           X_Logic0_port, B(23) => X_Logic0_port, B(22) => 
                           X_Logic0_port, B(21) => X_Logic0_port, B(20) => 
                           X_Logic0_port, B(19) => X_Logic0_port, B(18) => 
                           X_Logic0_port, B(17) => X_Logic0_port, B(16) => 
                           X_Logic0_port, B(15) => X_Logic0_port, B(14) => 
                           X_Logic0_port, B(13) => X_Logic0_port, B(12) => 
                           X_Logic0_port, B(11) => X_Logic0_port, B(10) => 
                           X_Logic0_port, B(9) => X_Logic0_port, B(8) => 
                           X_Logic0_port, B(7) => X_Logic0_port, B(6) => 
                           X_Logic0_port, B(5) => X_Logic0_port, B(4) => 
                           X_Logic0_port, B(3) => X_Logic0_port, B(2) => 
                           X_Logic0_port, B(1) => X_Logic0_port, B(0) => 
                           X_Logic0_port, Ci => X_Logic1_port, S(63) => 
                           negative_inputs_0_63_port, S(62) => 
                           negative_inputs_0_62_port, S(61) => 
                           negative_inputs_0_61_port, S(60) => 
                           negative_inputs_0_60_port, S(59) => 
                           negative_inputs_0_59_port, S(58) => 
                           negative_inputs_0_58_port, S(57) => 
                           negative_inputs_0_57_port, S(56) => 
                           negative_inputs_0_56_port, S(55) => 
                           negative_inputs_0_55_port, S(54) => 
                           negative_inputs_0_54_port, S(53) => 
                           negative_inputs_0_53_port, S(52) => 
                           negative_inputs_0_52_port, S(51) => 
                           negative_inputs_0_51_port, S(50) => 
                           negative_inputs_0_50_port, S(49) => 
                           negative_inputs_0_49_port, S(48) => 
                           negative_inputs_0_48_port, S(47) => 
                           negative_inputs_0_47_port, S(46) => 
                           negative_inputs_0_46_port, S(45) => 
                           negative_inputs_0_45_port, S(44) => 
                           negative_inputs_0_44_port, S(43) => 
                           negative_inputs_0_43_port, S(42) => 
                           negative_inputs_0_42_port, S(41) => 
                           negative_inputs_0_41_port, S(40) => 
                           negative_inputs_0_40_port, S(39) => 
                           negative_inputs_0_39_port, S(38) => 
                           negative_inputs_0_38_port, S(37) => 
                           negative_inputs_0_37_port, S(36) => 
                           negative_inputs_0_36_port, S(35) => 
                           negative_inputs_0_35_port, S(34) => 
                           negative_inputs_0_34_port, S(33) => 
                           negative_inputs_0_33_port, S(32) => 
                           negative_inputs_0_32_port, S(31) => 
                           negative_inputs_0_31_port, S(30) => 
                           negative_inputs_0_30_port, S(29) => 
                           negative_inputs_0_29_port, S(28) => 
                           negative_inputs_0_28_port, S(27) => 
                           negative_inputs_0_27_port, S(26) => 
                           negative_inputs_0_26_port, S(25) => 
                           negative_inputs_0_25_port, S(24) => 
                           negative_inputs_0_24_port, S(23) => 
                           negative_inputs_0_23_port, S(22) => 
                           negative_inputs_0_22_port, S(21) => 
                           negative_inputs_0_21_port, S(20) => 
                           negative_inputs_0_20_port, S(19) => 
                           negative_inputs_0_19_port, S(18) => 
                           negative_inputs_0_18_port, S(17) => 
                           negative_inputs_0_17_port, S(16) => 
                           negative_inputs_0_16_port, S(15) => 
                           negative_inputs_0_15_port, S(14) => 
                           negative_inputs_0_14_port, S(13) => 
                           negative_inputs_0_13_port, S(12) => 
                           negative_inputs_0_12_port, S(11) => 
                           negative_inputs_0_11_port, S(10) => 
                           negative_inputs_0_10_port, S(9) => 
                           negative_inputs_0_9_port, S(8) => 
                           negative_inputs_0_8_port, S(7) => 
                           negative_inputs_0_7_port, S(6) => 
                           negative_inputs_0_6_port, S(5) => 
                           negative_inputs_0_5_port, S(4) => 
                           negative_inputs_0_4_port, S(3) => 
                           negative_inputs_0_3_port, S(2) => 
                           negative_inputs_0_2_port, S(1) => 
                           negative_inputs_0_1_port, S(0) => 
                           negative_inputs_0_0_port, Co => n_1000);
   shifted_pos_1 : leftshifter_NbitShifter64_0 port map( shift_in(63) => A(31),
                           shift_in(62) => A(31), shift_in(61) => A(31), 
                           shift_in(60) => A(31), shift_in(59) => A(31), 
                           shift_in(58) => A(31), shift_in(57) => A(31), 
                           shift_in(56) => A(31), shift_in(55) => A(31), 
                           shift_in(54) => A(31), shift_in(53) => A(31), 
                           shift_in(52) => A(31), shift_in(51) => A(31), 
                           shift_in(50) => A(31), shift_in(49) => A(31), 
                           shift_in(48) => A(31), shift_in(47) => A(31), 
                           shift_in(46) => A(31), shift_in(45) => A(31), 
                           shift_in(44) => A(31), shift_in(43) => A(31), 
                           shift_in(42) => A(31), shift_in(41) => A(31), 
                           shift_in(40) => A(31), shift_in(39) => A(31), 
                           shift_in(38) => A(31), shift_in(37) => A(31), 
                           shift_in(36) => A(31), shift_in(35) => A(31), 
                           shift_in(34) => A(31), shift_in(33) => A(31), 
                           shift_in(32) => A(31), shift_in(31) => A(31), 
                           shift_in(30) => A(30), shift_in(29) => A(29), 
                           shift_in(28) => A(28), shift_in(27) => A(27), 
                           shift_in(26) => A(26), shift_in(25) => A(25), 
                           shift_in(24) => A(24), shift_in(23) => A(23), 
                           shift_in(22) => A(22), shift_in(21) => A(21), 
                           shift_in(20) => A(20), shift_in(19) => A(19), 
                           shift_in(18) => A(18), shift_in(17) => A(17), 
                           shift_in(16) => A(16), shift_in(15) => A(15), 
                           shift_in(14) => A(14), shift_in(13) => A(13), 
                           shift_in(12) => A(12), shift_in(11) => A(11), 
                           shift_in(10) => A(10), shift_in(9) => A(9), 
                           shift_in(8) => A(8), shift_in(7) => A(7), 
                           shift_in(6) => A(6), shift_in(5) => A(5), 
                           shift_in(4) => A(4), shift_in(3) => A(3), 
                           shift_in(2) => A(2), shift_in(1) => n11, shift_in(0)
                           => n72, shift_out(63) => positive_inputs_1_63_port, 
                           shift_out(62) => positive_inputs_1_62_port, 
                           shift_out(61) => positive_inputs_1_61_port, 
                           shift_out(60) => positive_inputs_1_60_port, 
                           shift_out(59) => positive_inputs_1_59_port, 
                           shift_out(58) => positive_inputs_1_58_port, 
                           shift_out(57) => positive_inputs_1_57_port, 
                           shift_out(56) => positive_inputs_1_56_port, 
                           shift_out(55) => positive_inputs_1_55_port, 
                           shift_out(54) => positive_inputs_1_54_port, 
                           shift_out(53) => positive_inputs_1_53_port, 
                           shift_out(52) => positive_inputs_1_52_port, 
                           shift_out(51) => positive_inputs_1_51_port, 
                           shift_out(50) => positive_inputs_1_50_port, 
                           shift_out(49) => positive_inputs_1_49_port, 
                           shift_out(48) => positive_inputs_1_48_port, 
                           shift_out(47) => positive_inputs_1_47_port, 
                           shift_out(46) => positive_inputs_1_46_port, 
                           shift_out(45) => positive_inputs_1_45_port, 
                           shift_out(44) => positive_inputs_1_44_port, 
                           shift_out(43) => positive_inputs_1_43_port, 
                           shift_out(42) => positive_inputs_1_42_port, 
                           shift_out(41) => positive_inputs_1_41_port, 
                           shift_out(40) => positive_inputs_1_40_port, 
                           shift_out(39) => positive_inputs_1_39_port, 
                           shift_out(38) => positive_inputs_1_38_port, 
                           shift_out(37) => positive_inputs_1_37_port, 
                           shift_out(36) => positive_inputs_1_36_port, 
                           shift_out(35) => positive_inputs_1_35_port, 
                           shift_out(34) => positive_inputs_1_34_port, 
                           shift_out(33) => positive_inputs_1_33_port, 
                           shift_out(32) => positive_inputs_1_32_port, 
                           shift_out(31) => positive_inputs_1_31_port, 
                           shift_out(30) => positive_inputs_1_30_port, 
                           shift_out(29) => positive_inputs_1_29_port, 
                           shift_out(28) => positive_inputs_1_28_port, 
                           shift_out(27) => positive_inputs_1_27_port, 
                           shift_out(26) => positive_inputs_1_26_port, 
                           shift_out(25) => positive_inputs_1_25_port, 
                           shift_out(24) => positive_inputs_1_24_port, 
                           shift_out(23) => positive_inputs_1_23_port, 
                           shift_out(22) => positive_inputs_1_22_port, 
                           shift_out(21) => positive_inputs_1_21_port, 
                           shift_out(20) => positive_inputs_1_20_port, 
                           shift_out(19) => positive_inputs_1_19_port, 
                           shift_out(18) => positive_inputs_1_18_port, 
                           shift_out(17) => positive_inputs_1_17_port, 
                           shift_out(16) => positive_inputs_1_16_port, 
                           shift_out(15) => positive_inputs_1_15_port, 
                           shift_out(14) => positive_inputs_1_14_port, 
                           shift_out(13) => positive_inputs_1_13_port, 
                           shift_out(12) => positive_inputs_1_12_port, 
                           shift_out(11) => positive_inputs_1_11_port, 
                           shift_out(10) => positive_inputs_1_10_port, 
                           shift_out(9) => positive_inputs_1_9_port, 
                           shift_out(8) => positive_inputs_1_8_port, 
                           shift_out(7) => positive_inputs_1_7_port, 
                           shift_out(6) => positive_inputs_1_6_port, 
                           shift_out(5) => positive_inputs_1_5_port, 
                           shift_out(4) => positive_inputs_1_4_port, 
                           shift_out(3) => positive_inputs_1_3_port, 
                           shift_out(2) => positive_inputs_1_2_port, 
                           shift_out(1) => positive_inputs_1_1_port, 
                           shift_out(0) => n_1001);
   shifted_pos_2 : leftshifter_NbitShifter64_62 port map( shift_in(63) => 
                           positive_inputs_1_63_port, shift_in(62) => 
                           positive_inputs_1_62_port, shift_in(61) => 
                           positive_inputs_1_61_port, shift_in(60) => 
                           positive_inputs_1_60_port, shift_in(59) => 
                           positive_inputs_1_59_port, shift_in(58) => 
                           positive_inputs_1_58_port, shift_in(57) => 
                           positive_inputs_1_57_port, shift_in(56) => 
                           positive_inputs_1_56_port, shift_in(55) => 
                           positive_inputs_1_55_port, shift_in(54) => 
                           positive_inputs_1_54_port, shift_in(53) => 
                           positive_inputs_1_53_port, shift_in(52) => 
                           positive_inputs_1_52_port, shift_in(51) => 
                           positive_inputs_1_51_port, shift_in(50) => 
                           positive_inputs_1_50_port, shift_in(49) => 
                           positive_inputs_1_49_port, shift_in(48) => n70, 
                           shift_in(47) => positive_inputs_1_47_port, 
                           shift_in(46) => positive_inputs_1_46_port, 
                           shift_in(45) => positive_inputs_1_45_port, 
                           shift_in(44) => positive_inputs_1_44_port, 
                           shift_in(43) => positive_inputs_1_43_port, 
                           shift_in(42) => positive_inputs_1_42_port, 
                           shift_in(41) => positive_inputs_1_41_port, 
                           shift_in(40) => positive_inputs_1_40_port, 
                           shift_in(39) => positive_inputs_1_39_port, 
                           shift_in(38) => n50, shift_in(37) => 
                           positive_inputs_1_37_port, shift_in(36) => 
                           positive_inputs_1_36_port, shift_in(35) => 
                           positive_inputs_1_35_port, shift_in(34) => 
                           positive_inputs_1_34_port, shift_in(33) => 
                           positive_inputs_1_33_port, shift_in(32) => 
                           positive_inputs_1_32_port, shift_in(31) => 
                           positive_inputs_1_31_port, shift_in(30) => 
                           positive_inputs_1_30_port, shift_in(29) => 
                           positive_inputs_1_29_port, shift_in(28) => 
                           positive_inputs_1_28_port, shift_in(27) => 
                           positive_inputs_1_27_port, shift_in(26) => 
                           positive_inputs_1_26_port, shift_in(25) => 
                           positive_inputs_1_25_port, shift_in(24) => 
                           positive_inputs_1_24_port, shift_in(23) => 
                           positive_inputs_1_23_port, shift_in(22) => 
                           positive_inputs_1_22_port, shift_in(21) => 
                           positive_inputs_1_21_port, shift_in(20) => 
                           positive_inputs_1_20_port, shift_in(19) => 
                           positive_inputs_1_19_port, shift_in(18) => 
                           positive_inputs_1_18_port, shift_in(17) => 
                           positive_inputs_1_17_port, shift_in(16) => 
                           positive_inputs_1_16_port, shift_in(15) => 
                           positive_inputs_1_15_port, shift_in(14) => 
                           positive_inputs_1_14_port, shift_in(13) => 
                           positive_inputs_1_13_port, shift_in(12) => 
                           positive_inputs_1_12_port, shift_in(11) => 
                           positive_inputs_1_11_port, shift_in(10) => 
                           positive_inputs_1_10_port, shift_in(9) => 
                           positive_inputs_1_9_port, shift_in(8) => 
                           positive_inputs_1_8_port, shift_in(7) => 
                           positive_inputs_1_7_port, shift_in(6) => 
                           positive_inputs_1_6_port, shift_in(5) => 
                           positive_inputs_1_5_port, shift_in(4) => 
                           positive_inputs_1_4_port, shift_in(3) => 
                           positive_inputs_1_3_port, shift_in(2) => 
                           positive_inputs_1_2_port, shift_in(1) => 
                           positive_inputs_1_1_port, shift_in(0) => n9, 
                           shift_out(63) => positive_inputs_2_63_port, 
                           shift_out(62) => positive_inputs_2_62_port, 
                           shift_out(61) => positive_inputs_2_61_port, 
                           shift_out(60) => positive_inputs_2_60_port, 
                           shift_out(59) => positive_inputs_2_59_port, 
                           shift_out(58) => positive_inputs_2_58_port, 
                           shift_out(57) => positive_inputs_2_57_port, 
                           shift_out(56) => positive_inputs_2_56_port, 
                           shift_out(55) => positive_inputs_2_55_port, 
                           shift_out(54) => positive_inputs_2_54_port, 
                           shift_out(53) => positive_inputs_2_53_port, 
                           shift_out(52) => positive_inputs_2_52_port, 
                           shift_out(51) => positive_inputs_2_51_port, 
                           shift_out(50) => positive_inputs_2_50_port, 
                           shift_out(49) => positive_inputs_2_49_port, 
                           shift_out(48) => positive_inputs_2_48_port, 
                           shift_out(47) => positive_inputs_2_47_port, 
                           shift_out(46) => positive_inputs_2_46_port, 
                           shift_out(45) => positive_inputs_2_45_port, 
                           shift_out(44) => positive_inputs_2_44_port, 
                           shift_out(43) => positive_inputs_2_43_port, 
                           shift_out(42) => positive_inputs_2_42_port, 
                           shift_out(41) => positive_inputs_2_41_port, 
                           shift_out(40) => positive_inputs_2_40_port, 
                           shift_out(39) => positive_inputs_2_39_port, 
                           shift_out(38) => positive_inputs_2_38_port, 
                           shift_out(37) => positive_inputs_2_37_port, 
                           shift_out(36) => positive_inputs_2_36_port, 
                           shift_out(35) => positive_inputs_2_35_port, 
                           shift_out(34) => positive_inputs_2_34_port, 
                           shift_out(33) => positive_inputs_2_33_port, 
                           shift_out(32) => positive_inputs_2_32_port, 
                           shift_out(31) => positive_inputs_2_31_port, 
                           shift_out(30) => positive_inputs_2_30_port, 
                           shift_out(29) => positive_inputs_2_29_port, 
                           shift_out(28) => positive_inputs_2_28_port, 
                           shift_out(27) => positive_inputs_2_27_port, 
                           shift_out(26) => positive_inputs_2_26_port, 
                           shift_out(25) => positive_inputs_2_25_port, 
                           shift_out(24) => positive_inputs_2_24_port, 
                           shift_out(23) => positive_inputs_2_23_port, 
                           shift_out(22) => positive_inputs_2_22_port, 
                           shift_out(21) => positive_inputs_2_21_port, 
                           shift_out(20) => positive_inputs_2_20_port, 
                           shift_out(19) => positive_inputs_2_19_port, 
                           shift_out(18) => positive_inputs_2_18_port, 
                           shift_out(17) => positive_inputs_2_17_port, 
                           shift_out(16) => positive_inputs_2_16_port, 
                           shift_out(15) => positive_inputs_2_15_port, 
                           shift_out(14) => positive_inputs_2_14_port, 
                           shift_out(13) => positive_inputs_2_13_port, 
                           shift_out(12) => positive_inputs_2_12_port, 
                           shift_out(11) => positive_inputs_2_11_port, 
                           shift_out(10) => positive_inputs_2_10_port, 
                           shift_out(9) => positive_inputs_2_9_port, 
                           shift_out(8) => positive_inputs_2_8_port, 
                           shift_out(7) => positive_inputs_2_7_port, 
                           shift_out(6) => positive_inputs_2_6_port, 
                           shift_out(5) => positive_inputs_2_5_port, 
                           shift_out(4) => positive_inputs_2_4_port, 
                           shift_out(3) => positive_inputs_2_3_port, 
                           shift_out(2) => positive_inputs_2_2_port, 
                           shift_out(1) => positive_inputs_2_1_port, 
                           shift_out(0) => n_1002);
   shifted_pos_3 : leftshifter_NbitShifter64_61 port map( shift_in(63) => 
                           positive_inputs_2_63_port, shift_in(62) => 
                           positive_inputs_2_62_port, shift_in(61) => 
                           positive_inputs_2_61_port, shift_in(60) => 
                           positive_inputs_2_60_port, shift_in(59) => 
                           positive_inputs_2_59_port, shift_in(58) => 
                           positive_inputs_2_58_port, shift_in(57) => 
                           positive_inputs_2_57_port, shift_in(56) => 
                           positive_inputs_2_56_port, shift_in(55) => 
                           positive_inputs_2_55_port, shift_in(54) => 
                           positive_inputs_2_54_port, shift_in(53) => 
                           positive_inputs_2_53_port, shift_in(52) => 
                           positive_inputs_2_52_port, shift_in(51) => 
                           positive_inputs_2_51_port, shift_in(50) => 
                           positive_inputs_2_50_port, shift_in(49) => 
                           positive_inputs_2_49_port, shift_in(48) => n69, 
                           shift_in(47) => positive_inputs_2_47_port, 
                           shift_in(46) => positive_inputs_2_46_port, 
                           shift_in(45) => positive_inputs_2_45_port, 
                           shift_in(44) => positive_inputs_2_44_port, 
                           shift_in(43) => positive_inputs_2_43_port, 
                           shift_in(42) => positive_inputs_2_42_port, 
                           shift_in(41) => positive_inputs_2_41_port, 
                           shift_in(40) => positive_inputs_2_40_port, 
                           shift_in(39) => positive_inputs_2_39_port, 
                           shift_in(38) => n49, shift_in(37) => 
                           positive_inputs_2_37_port, shift_in(36) => 
                           positive_inputs_2_36_port, shift_in(35) => 
                           positive_inputs_2_35_port, shift_in(34) => 
                           positive_inputs_2_34_port, shift_in(33) => 
                           positive_inputs_2_33_port, shift_in(32) => 
                           positive_inputs_2_32_port, shift_in(31) => 
                           positive_inputs_2_31_port, shift_in(30) => 
                           positive_inputs_2_30_port, shift_in(29) => 
                           positive_inputs_2_29_port, shift_in(28) => 
                           positive_inputs_2_28_port, shift_in(27) => 
                           positive_inputs_2_27_port, shift_in(26) => 
                           positive_inputs_2_26_port, shift_in(25) => 
                           positive_inputs_2_25_port, shift_in(24) => 
                           positive_inputs_2_24_port, shift_in(23) => 
                           positive_inputs_2_23_port, shift_in(22) => 
                           positive_inputs_2_22_port, shift_in(21) => 
                           positive_inputs_2_21_port, shift_in(20) => 
                           positive_inputs_2_20_port, shift_in(19) => 
                           positive_inputs_2_19_port, shift_in(18) => 
                           positive_inputs_2_18_port, shift_in(17) => 
                           positive_inputs_2_17_port, shift_in(16) => 
                           positive_inputs_2_16_port, shift_in(15) => 
                           positive_inputs_2_15_port, shift_in(14) => 
                           positive_inputs_2_14_port, shift_in(13) => 
                           positive_inputs_2_13_port, shift_in(12) => 
                           positive_inputs_2_12_port, shift_in(11) => 
                           positive_inputs_2_11_port, shift_in(10) => 
                           positive_inputs_2_10_port, shift_in(9) => 
                           positive_inputs_2_9_port, shift_in(8) => 
                           positive_inputs_2_8_port, shift_in(7) => 
                           positive_inputs_2_7_port, shift_in(6) => 
                           positive_inputs_2_6_port, shift_in(5) => 
                           positive_inputs_2_5_port, shift_in(4) => 
                           positive_inputs_2_4_port, shift_in(3) => 
                           positive_inputs_2_3_port, shift_in(2) => 
                           positive_inputs_2_2_port, shift_in(1) => 
                           positive_inputs_2_1_port, shift_in(0) => n9, 
                           shift_out(63) => positive_inputs_3_63_port, 
                           shift_out(62) => positive_inputs_3_62_port, 
                           shift_out(61) => positive_inputs_3_61_port, 
                           shift_out(60) => positive_inputs_3_60_port, 
                           shift_out(59) => positive_inputs_3_59_port, 
                           shift_out(58) => positive_inputs_3_58_port, 
                           shift_out(57) => positive_inputs_3_57_port, 
                           shift_out(56) => positive_inputs_3_56_port, 
                           shift_out(55) => positive_inputs_3_55_port, 
                           shift_out(54) => positive_inputs_3_54_port, 
                           shift_out(53) => positive_inputs_3_53_port, 
                           shift_out(52) => positive_inputs_3_52_port, 
                           shift_out(51) => positive_inputs_3_51_port, 
                           shift_out(50) => positive_inputs_3_50_port, 
                           shift_out(49) => positive_inputs_3_49_port, 
                           shift_out(48) => positive_inputs_3_48_port, 
                           shift_out(47) => positive_inputs_3_47_port, 
                           shift_out(46) => positive_inputs_3_46_port, 
                           shift_out(45) => positive_inputs_3_45_port, 
                           shift_out(44) => positive_inputs_3_44_port, 
                           shift_out(43) => positive_inputs_3_43_port, 
                           shift_out(42) => positive_inputs_3_42_port, 
                           shift_out(41) => positive_inputs_3_41_port, 
                           shift_out(40) => positive_inputs_3_40_port, 
                           shift_out(39) => positive_inputs_3_39_port, 
                           shift_out(38) => positive_inputs_3_38_port, 
                           shift_out(37) => positive_inputs_3_37_port, 
                           shift_out(36) => positive_inputs_3_36_port, 
                           shift_out(35) => positive_inputs_3_35_port, 
                           shift_out(34) => positive_inputs_3_34_port, 
                           shift_out(33) => positive_inputs_3_33_port, 
                           shift_out(32) => positive_inputs_3_32_port, 
                           shift_out(31) => positive_inputs_3_31_port, 
                           shift_out(30) => positive_inputs_3_30_port, 
                           shift_out(29) => positive_inputs_3_29_port, 
                           shift_out(28) => positive_inputs_3_28_port, 
                           shift_out(27) => positive_inputs_3_27_port, 
                           shift_out(26) => positive_inputs_3_26_port, 
                           shift_out(25) => positive_inputs_3_25_port, 
                           shift_out(24) => positive_inputs_3_24_port, 
                           shift_out(23) => positive_inputs_3_23_port, 
                           shift_out(22) => positive_inputs_3_22_port, 
                           shift_out(21) => positive_inputs_3_21_port, 
                           shift_out(20) => positive_inputs_3_20_port, 
                           shift_out(19) => positive_inputs_3_19_port, 
                           shift_out(18) => positive_inputs_3_18_port, 
                           shift_out(17) => positive_inputs_3_17_port, 
                           shift_out(16) => positive_inputs_3_16_port, 
                           shift_out(15) => positive_inputs_3_15_port, 
                           shift_out(14) => positive_inputs_3_14_port, 
                           shift_out(13) => positive_inputs_3_13_port, 
                           shift_out(12) => positive_inputs_3_12_port, 
                           shift_out(11) => positive_inputs_3_11_port, 
                           shift_out(10) => positive_inputs_3_10_port, 
                           shift_out(9) => positive_inputs_3_9_port, 
                           shift_out(8) => positive_inputs_3_8_port, 
                           shift_out(7) => positive_inputs_3_7_port, 
                           shift_out(6) => positive_inputs_3_6_port, 
                           shift_out(5) => positive_inputs_3_5_port, 
                           shift_out(4) => positive_inputs_3_4_port, 
                           shift_out(3) => positive_inputs_3_3_port, 
                           shift_out(2) => positive_inputs_3_2_port, 
                           shift_out(1) => positive_inputs_3_1_port, 
                           shift_out(0) => n_1003);
   shifted_pos_4 : leftshifter_NbitShifter64_60 port map( shift_in(63) => 
                           positive_inputs_3_63_port, shift_in(62) => 
                           positive_inputs_3_62_port, shift_in(61) => 
                           positive_inputs_3_61_port, shift_in(60) => 
                           positive_inputs_3_60_port, shift_in(59) => 
                           positive_inputs_3_59_port, shift_in(58) => 
                           positive_inputs_3_58_port, shift_in(57) => 
                           positive_inputs_3_57_port, shift_in(56) => 
                           positive_inputs_3_56_port, shift_in(55) => 
                           positive_inputs_3_55_port, shift_in(54) => 
                           positive_inputs_3_54_port, shift_in(53) => 
                           positive_inputs_3_53_port, shift_in(52) => 
                           positive_inputs_3_52_port, shift_in(51) => 
                           positive_inputs_3_51_port, shift_in(50) => 
                           positive_inputs_3_50_port, shift_in(49) => 
                           positive_inputs_3_49_port, shift_in(48) => 
                           positive_inputs_3_48_port, shift_in(47) => 
                           positive_inputs_3_47_port, shift_in(46) => 
                           positive_inputs_3_46_port, shift_in(45) => 
                           positive_inputs_3_45_port, shift_in(44) => 
                           positive_inputs_3_44_port, shift_in(43) => 
                           positive_inputs_3_43_port, shift_in(42) => 
                           positive_inputs_3_42_port, shift_in(41) => 
                           positive_inputs_3_41_port, shift_in(40) => 
                           positive_inputs_3_40_port, shift_in(39) => 
                           positive_inputs_3_39_port, shift_in(38) => 
                           positive_inputs_3_38_port, shift_in(37) => 
                           positive_inputs_3_37_port, shift_in(36) => 
                           positive_inputs_3_36_port, shift_in(35) => 
                           positive_inputs_3_35_port, shift_in(34) => 
                           positive_inputs_3_34_port, shift_in(33) => 
                           positive_inputs_3_33_port, shift_in(32) => 
                           positive_inputs_3_32_port, shift_in(31) => 
                           positive_inputs_3_31_port, shift_in(30) => 
                           positive_inputs_3_30_port, shift_in(29) => 
                           positive_inputs_3_29_port, shift_in(28) => 
                           positive_inputs_3_28_port, shift_in(27) => 
                           positive_inputs_3_27_port, shift_in(26) => 
                           positive_inputs_3_26_port, shift_in(25) => 
                           positive_inputs_3_25_port, shift_in(24) => 
                           positive_inputs_3_24_port, shift_in(23) => 
                           positive_inputs_3_23_port, shift_in(22) => 
                           positive_inputs_3_22_port, shift_in(21) => 
                           positive_inputs_3_21_port, shift_in(20) => 
                           positive_inputs_3_20_port, shift_in(19) => 
                           positive_inputs_3_19_port, shift_in(18) => 
                           positive_inputs_3_18_port, shift_in(17) => 
                           positive_inputs_3_17_port, shift_in(16) => 
                           positive_inputs_3_16_port, shift_in(15) => 
                           positive_inputs_3_15_port, shift_in(14) => 
                           positive_inputs_3_14_port, shift_in(13) => 
                           positive_inputs_3_13_port, shift_in(12) => 
                           positive_inputs_3_12_port, shift_in(11) => 
                           positive_inputs_3_11_port, shift_in(10) => 
                           positive_inputs_3_10_port, shift_in(9) => 
                           positive_inputs_3_9_port, shift_in(8) => 
                           positive_inputs_3_8_port, shift_in(7) => 
                           positive_inputs_3_7_port, shift_in(6) => 
                           positive_inputs_3_6_port, shift_in(5) => 
                           positive_inputs_3_5_port, shift_in(4) => 
                           positive_inputs_3_4_port, shift_in(3) => 
                           positive_inputs_3_3_port, shift_in(2) => 
                           positive_inputs_3_2_port, shift_in(1) => 
                           positive_inputs_3_1_port, shift_in(0) => n9, 
                           shift_out(63) => positive_inputs_4_63_port, 
                           shift_out(62) => positive_inputs_4_62_port, 
                           shift_out(61) => positive_inputs_4_61_port, 
                           shift_out(60) => positive_inputs_4_60_port, 
                           shift_out(59) => positive_inputs_4_59_port, 
                           shift_out(58) => positive_inputs_4_58_port, 
                           shift_out(57) => positive_inputs_4_57_port, 
                           shift_out(56) => positive_inputs_4_56_port, 
                           shift_out(55) => positive_inputs_4_55_port, 
                           shift_out(54) => positive_inputs_4_54_port, 
                           shift_out(53) => positive_inputs_4_53_port, 
                           shift_out(52) => positive_inputs_4_52_port, 
                           shift_out(51) => positive_inputs_4_51_port, 
                           shift_out(50) => positive_inputs_4_50_port, 
                           shift_out(49) => positive_inputs_4_49_port, 
                           shift_out(48) => positive_inputs_4_48_port, 
                           shift_out(47) => positive_inputs_4_47_port, 
                           shift_out(46) => positive_inputs_4_46_port, 
                           shift_out(45) => positive_inputs_4_45_port, 
                           shift_out(44) => positive_inputs_4_44_port, 
                           shift_out(43) => positive_inputs_4_43_port, 
                           shift_out(42) => positive_inputs_4_42_port, 
                           shift_out(41) => positive_inputs_4_41_port, 
                           shift_out(40) => positive_inputs_4_40_port, 
                           shift_out(39) => positive_inputs_4_39_port, 
                           shift_out(38) => positive_inputs_4_38_port, 
                           shift_out(37) => positive_inputs_4_37_port, 
                           shift_out(36) => positive_inputs_4_36_port, 
                           shift_out(35) => positive_inputs_4_35_port, 
                           shift_out(34) => positive_inputs_4_34_port, 
                           shift_out(33) => positive_inputs_4_33_port, 
                           shift_out(32) => positive_inputs_4_32_port, 
                           shift_out(31) => positive_inputs_4_31_port, 
                           shift_out(30) => positive_inputs_4_30_port, 
                           shift_out(29) => positive_inputs_4_29_port, 
                           shift_out(28) => positive_inputs_4_28_port, 
                           shift_out(27) => positive_inputs_4_27_port, 
                           shift_out(26) => positive_inputs_4_26_port, 
                           shift_out(25) => positive_inputs_4_25_port, 
                           shift_out(24) => positive_inputs_4_24_port, 
                           shift_out(23) => positive_inputs_4_23_port, 
                           shift_out(22) => positive_inputs_4_22_port, 
                           shift_out(21) => positive_inputs_4_21_port, 
                           shift_out(20) => positive_inputs_4_20_port, 
                           shift_out(19) => positive_inputs_4_19_port, 
                           shift_out(18) => positive_inputs_4_18_port, 
                           shift_out(17) => positive_inputs_4_17_port, 
                           shift_out(16) => positive_inputs_4_16_port, 
                           shift_out(15) => positive_inputs_4_15_port, 
                           shift_out(14) => positive_inputs_4_14_port, 
                           shift_out(13) => positive_inputs_4_13_port, 
                           shift_out(12) => positive_inputs_4_12_port, 
                           shift_out(11) => positive_inputs_4_11_port, 
                           shift_out(10) => positive_inputs_4_10_port, 
                           shift_out(9) => positive_inputs_4_9_port, 
                           shift_out(8) => positive_inputs_4_8_port, 
                           shift_out(7) => positive_inputs_4_7_port, 
                           shift_out(6) => positive_inputs_4_6_port, 
                           shift_out(5) => positive_inputs_4_5_port, 
                           shift_out(4) => positive_inputs_4_4_port, 
                           shift_out(3) => positive_inputs_4_3_port, 
                           shift_out(2) => positive_inputs_4_2_port, 
                           shift_out(1) => positive_inputs_4_1_port, 
                           shift_out(0) => n_1004);
   shifted_pos_5 : leftshifter_NbitShifter64_59 port map( shift_in(63) => 
                           positive_inputs_4_63_port, shift_in(62) => 
                           positive_inputs_4_62_port, shift_in(61) => 
                           positive_inputs_4_61_port, shift_in(60) => 
                           positive_inputs_4_60_port, shift_in(59) => 
                           positive_inputs_4_59_port, shift_in(58) => 
                           positive_inputs_4_58_port, shift_in(57) => 
                           positive_inputs_4_57_port, shift_in(56) => 
                           positive_inputs_4_56_port, shift_in(55) => 
                           positive_inputs_4_55_port, shift_in(54) => 
                           positive_inputs_4_54_port, shift_in(53) => 
                           positive_inputs_4_53_port, shift_in(52) => 
                           positive_inputs_4_52_port, shift_in(51) => 
                           positive_inputs_4_51_port, shift_in(50) => 
                           positive_inputs_4_50_port, shift_in(49) => 
                           positive_inputs_4_49_port, shift_in(48) => n68, 
                           shift_in(47) => positive_inputs_4_47_port, 
                           shift_in(46) => positive_inputs_4_46_port, 
                           shift_in(45) => positive_inputs_4_45_port, 
                           shift_in(44) => positive_inputs_4_44_port, 
                           shift_in(43) => positive_inputs_4_43_port, 
                           shift_in(42) => positive_inputs_4_42_port, 
                           shift_in(41) => positive_inputs_4_41_port, 
                           shift_in(40) => positive_inputs_4_40_port, 
                           shift_in(39) => n55, shift_in(38) => 
                           positive_inputs_4_38_port, shift_in(37) => 
                           positive_inputs_4_37_port, shift_in(36) => 
                           positive_inputs_4_36_port, shift_in(35) => 
                           positive_inputs_4_35_port, shift_in(34) => 
                           positive_inputs_4_34_port, shift_in(33) => 
                           positive_inputs_4_33_port, shift_in(32) => 
                           positive_inputs_4_32_port, shift_in(31) => 
                           positive_inputs_4_31_port, shift_in(30) => 
                           positive_inputs_4_30_port, shift_in(29) => 
                           positive_inputs_4_29_port, shift_in(28) => 
                           positive_inputs_4_28_port, shift_in(27) => 
                           positive_inputs_4_27_port, shift_in(26) => 
                           positive_inputs_4_26_port, shift_in(25) => 
                           positive_inputs_4_25_port, shift_in(24) => 
                           positive_inputs_4_24_port, shift_in(23) => 
                           positive_inputs_4_23_port, shift_in(22) => 
                           positive_inputs_4_22_port, shift_in(21) => 
                           positive_inputs_4_21_port, shift_in(20) => 
                           positive_inputs_4_20_port, shift_in(19) => 
                           positive_inputs_4_19_port, shift_in(18) => 
                           positive_inputs_4_18_port, shift_in(17) => 
                           positive_inputs_4_17_port, shift_in(16) => 
                           positive_inputs_4_16_port, shift_in(15) => 
                           positive_inputs_4_15_port, shift_in(14) => 
                           positive_inputs_4_14_port, shift_in(13) => 
                           positive_inputs_4_13_port, shift_in(12) => 
                           positive_inputs_4_12_port, shift_in(11) => 
                           positive_inputs_4_11_port, shift_in(10) => 
                           positive_inputs_4_10_port, shift_in(9) => 
                           positive_inputs_4_9_port, shift_in(8) => 
                           positive_inputs_4_8_port, shift_in(7) => 
                           positive_inputs_4_7_port, shift_in(6) => 
                           positive_inputs_4_6_port, shift_in(5) => 
                           positive_inputs_4_5_port, shift_in(4) => 
                           positive_inputs_4_4_port, shift_in(3) => 
                           positive_inputs_4_3_port, shift_in(2) => 
                           positive_inputs_4_2_port, shift_in(1) => 
                           positive_inputs_4_1_port, shift_in(0) => n9, 
                           shift_out(63) => positive_inputs_5_63_port, 
                           shift_out(62) => positive_inputs_5_62_port, 
                           shift_out(61) => positive_inputs_5_61_port, 
                           shift_out(60) => positive_inputs_5_60_port, 
                           shift_out(59) => positive_inputs_5_59_port, 
                           shift_out(58) => positive_inputs_5_58_port, 
                           shift_out(57) => positive_inputs_5_57_port, 
                           shift_out(56) => positive_inputs_5_56_port, 
                           shift_out(55) => positive_inputs_5_55_port, 
                           shift_out(54) => positive_inputs_5_54_port, 
                           shift_out(53) => positive_inputs_5_53_port, 
                           shift_out(52) => positive_inputs_5_52_port, 
                           shift_out(51) => positive_inputs_5_51_port, 
                           shift_out(50) => positive_inputs_5_50_port, 
                           shift_out(49) => positive_inputs_5_49_port, 
                           shift_out(48) => positive_inputs_5_48_port, 
                           shift_out(47) => positive_inputs_5_47_port, 
                           shift_out(46) => positive_inputs_5_46_port, 
                           shift_out(45) => positive_inputs_5_45_port, 
                           shift_out(44) => positive_inputs_5_44_port, 
                           shift_out(43) => positive_inputs_5_43_port, 
                           shift_out(42) => positive_inputs_5_42_port, 
                           shift_out(41) => positive_inputs_5_41_port, 
                           shift_out(40) => positive_inputs_5_40_port, 
                           shift_out(39) => positive_inputs_5_39_port, 
                           shift_out(38) => positive_inputs_5_38_port, 
                           shift_out(37) => positive_inputs_5_37_port, 
                           shift_out(36) => positive_inputs_5_36_port, 
                           shift_out(35) => positive_inputs_5_35_port, 
                           shift_out(34) => positive_inputs_5_34_port, 
                           shift_out(33) => positive_inputs_5_33_port, 
                           shift_out(32) => positive_inputs_5_32_port, 
                           shift_out(31) => positive_inputs_5_31_port, 
                           shift_out(30) => positive_inputs_5_30_port, 
                           shift_out(29) => positive_inputs_5_29_port, 
                           shift_out(28) => positive_inputs_5_28_port, 
                           shift_out(27) => positive_inputs_5_27_port, 
                           shift_out(26) => positive_inputs_5_26_port, 
                           shift_out(25) => positive_inputs_5_25_port, 
                           shift_out(24) => positive_inputs_5_24_port, 
                           shift_out(23) => positive_inputs_5_23_port, 
                           shift_out(22) => positive_inputs_5_22_port, 
                           shift_out(21) => positive_inputs_5_21_port, 
                           shift_out(20) => positive_inputs_5_20_port, 
                           shift_out(19) => positive_inputs_5_19_port, 
                           shift_out(18) => positive_inputs_5_18_port, 
                           shift_out(17) => positive_inputs_5_17_port, 
                           shift_out(16) => positive_inputs_5_16_port, 
                           shift_out(15) => positive_inputs_5_15_port, 
                           shift_out(14) => positive_inputs_5_14_port, 
                           shift_out(13) => positive_inputs_5_13_port, 
                           shift_out(12) => positive_inputs_5_12_port, 
                           shift_out(11) => positive_inputs_5_11_port, 
                           shift_out(10) => positive_inputs_5_10_port, 
                           shift_out(9) => positive_inputs_5_9_port, 
                           shift_out(8) => positive_inputs_5_8_port, 
                           shift_out(7) => positive_inputs_5_7_port, 
                           shift_out(6) => positive_inputs_5_6_port, 
                           shift_out(5) => positive_inputs_5_5_port, 
                           shift_out(4) => positive_inputs_5_4_port, 
                           shift_out(3) => positive_inputs_5_3_port, 
                           shift_out(2) => positive_inputs_5_2_port, 
                           shift_out(1) => positive_inputs_5_1_port, 
                           shift_out(0) => n_1005);
   shifted_pos_6 : leftshifter_NbitShifter64_58 port map( shift_in(63) => 
                           positive_inputs_5_63_port, shift_in(62) => 
                           positive_inputs_5_62_port, shift_in(61) => 
                           positive_inputs_5_61_port, shift_in(60) => 
                           positive_inputs_5_60_port, shift_in(59) => 
                           positive_inputs_5_59_port, shift_in(58) => 
                           positive_inputs_5_58_port, shift_in(57) => 
                           positive_inputs_5_57_port, shift_in(56) => 
                           positive_inputs_5_56_port, shift_in(55) => 
                           positive_inputs_5_55_port, shift_in(54) => 
                           positive_inputs_5_54_port, shift_in(53) => 
                           positive_inputs_5_53_port, shift_in(52) => 
                           positive_inputs_5_52_port, shift_in(51) => 
                           positive_inputs_5_51_port, shift_in(50) => 
                           positive_inputs_5_50_port, shift_in(49) => 
                           positive_inputs_5_49_port, shift_in(48) => n67, 
                           shift_in(47) => positive_inputs_5_47_port, 
                           shift_in(46) => positive_inputs_5_46_port, 
                           shift_in(45) => positive_inputs_5_45_port, 
                           shift_in(44) => positive_inputs_5_44_port, 
                           shift_in(43) => positive_inputs_5_43_port, 
                           shift_in(42) => positive_inputs_5_42_port, 
                           shift_in(41) => positive_inputs_5_41_port, 
                           shift_in(40) => positive_inputs_5_40_port, 
                           shift_in(39) => n54, shift_in(38) => 
                           positive_inputs_5_38_port, shift_in(37) => 
                           positive_inputs_5_37_port, shift_in(36) => 
                           positive_inputs_5_36_port, shift_in(35) => 
                           positive_inputs_5_35_port, shift_in(34) => 
                           positive_inputs_5_34_port, shift_in(33) => 
                           positive_inputs_5_33_port, shift_in(32) => 
                           positive_inputs_5_32_port, shift_in(31) => 
                           positive_inputs_5_31_port, shift_in(30) => 
                           positive_inputs_5_30_port, shift_in(29) => 
                           positive_inputs_5_29_port, shift_in(28) => 
                           positive_inputs_5_28_port, shift_in(27) => 
                           positive_inputs_5_27_port, shift_in(26) => 
                           positive_inputs_5_26_port, shift_in(25) => 
                           positive_inputs_5_25_port, shift_in(24) => 
                           positive_inputs_5_24_port, shift_in(23) => 
                           positive_inputs_5_23_port, shift_in(22) => 
                           positive_inputs_5_22_port, shift_in(21) => 
                           positive_inputs_5_21_port, shift_in(20) => 
                           positive_inputs_5_20_port, shift_in(19) => 
                           positive_inputs_5_19_port, shift_in(18) => 
                           positive_inputs_5_18_port, shift_in(17) => 
                           positive_inputs_5_17_port, shift_in(16) => 
                           positive_inputs_5_16_port, shift_in(15) => 
                           positive_inputs_5_15_port, shift_in(14) => 
                           positive_inputs_5_14_port, shift_in(13) => 
                           positive_inputs_5_13_port, shift_in(12) => 
                           positive_inputs_5_12_port, shift_in(11) => 
                           positive_inputs_5_11_port, shift_in(10) => 
                           positive_inputs_5_10_port, shift_in(9) => 
                           positive_inputs_5_9_port, shift_in(8) => 
                           positive_inputs_5_8_port, shift_in(7) => 
                           positive_inputs_5_7_port, shift_in(6) => 
                           positive_inputs_5_6_port, shift_in(5) => 
                           positive_inputs_5_5_port, shift_in(4) => 
                           positive_inputs_5_4_port, shift_in(3) => 
                           positive_inputs_5_3_port, shift_in(2) => 
                           positive_inputs_5_2_port, shift_in(1) => 
                           positive_inputs_5_1_port, shift_in(0) => n9, 
                           shift_out(63) => positive_inputs_6_63_port, 
                           shift_out(62) => positive_inputs_6_62_port, 
                           shift_out(61) => positive_inputs_6_61_port, 
                           shift_out(60) => positive_inputs_6_60_port, 
                           shift_out(59) => positive_inputs_6_59_port, 
                           shift_out(58) => positive_inputs_6_58_port, 
                           shift_out(57) => positive_inputs_6_57_port, 
                           shift_out(56) => positive_inputs_6_56_port, 
                           shift_out(55) => positive_inputs_6_55_port, 
                           shift_out(54) => positive_inputs_6_54_port, 
                           shift_out(53) => positive_inputs_6_53_port, 
                           shift_out(52) => positive_inputs_6_52_port, 
                           shift_out(51) => positive_inputs_6_51_port, 
                           shift_out(50) => positive_inputs_6_50_port, 
                           shift_out(49) => positive_inputs_6_49_port, 
                           shift_out(48) => positive_inputs_6_48_port, 
                           shift_out(47) => positive_inputs_6_47_port, 
                           shift_out(46) => positive_inputs_6_46_port, 
                           shift_out(45) => positive_inputs_6_45_port, 
                           shift_out(44) => positive_inputs_6_44_port, 
                           shift_out(43) => positive_inputs_6_43_port, 
                           shift_out(42) => positive_inputs_6_42_port, 
                           shift_out(41) => positive_inputs_6_41_port, 
                           shift_out(40) => positive_inputs_6_40_port, 
                           shift_out(39) => positive_inputs_6_39_port, 
                           shift_out(38) => positive_inputs_6_38_port, 
                           shift_out(37) => positive_inputs_6_37_port, 
                           shift_out(36) => positive_inputs_6_36_port, 
                           shift_out(35) => positive_inputs_6_35_port, 
                           shift_out(34) => positive_inputs_6_34_port, 
                           shift_out(33) => positive_inputs_6_33_port, 
                           shift_out(32) => positive_inputs_6_32_port, 
                           shift_out(31) => positive_inputs_6_31_port, 
                           shift_out(30) => positive_inputs_6_30_port, 
                           shift_out(29) => positive_inputs_6_29_port, 
                           shift_out(28) => positive_inputs_6_28_port, 
                           shift_out(27) => positive_inputs_6_27_port, 
                           shift_out(26) => positive_inputs_6_26_port, 
                           shift_out(25) => positive_inputs_6_25_port, 
                           shift_out(24) => positive_inputs_6_24_port, 
                           shift_out(23) => positive_inputs_6_23_port, 
                           shift_out(22) => positive_inputs_6_22_port, 
                           shift_out(21) => positive_inputs_6_21_port, 
                           shift_out(20) => positive_inputs_6_20_port, 
                           shift_out(19) => positive_inputs_6_19_port, 
                           shift_out(18) => positive_inputs_6_18_port, 
                           shift_out(17) => positive_inputs_6_17_port, 
                           shift_out(16) => positive_inputs_6_16_port, 
                           shift_out(15) => positive_inputs_6_15_port, 
                           shift_out(14) => positive_inputs_6_14_port, 
                           shift_out(13) => positive_inputs_6_13_port, 
                           shift_out(12) => positive_inputs_6_12_port, 
                           shift_out(11) => positive_inputs_6_11_port, 
                           shift_out(10) => positive_inputs_6_10_port, 
                           shift_out(9) => positive_inputs_6_9_port, 
                           shift_out(8) => positive_inputs_6_8_port, 
                           shift_out(7) => positive_inputs_6_7_port, 
                           shift_out(6) => positive_inputs_6_6_port, 
                           shift_out(5) => positive_inputs_6_5_port, 
                           shift_out(4) => positive_inputs_6_4_port, 
                           shift_out(3) => positive_inputs_6_3_port, 
                           shift_out(2) => positive_inputs_6_2_port, 
                           shift_out(1) => positive_inputs_6_1_port, 
                           shift_out(0) => n_1006);
   shifted_pos_7 : leftshifter_NbitShifter64_57 port map( shift_in(63) => 
                           positive_inputs_6_63_port, shift_in(62) => 
                           positive_inputs_6_62_port, shift_in(61) => 
                           positive_inputs_6_61_port, shift_in(60) => 
                           positive_inputs_6_60_port, shift_in(59) => 
                           positive_inputs_6_59_port, shift_in(58) => 
                           positive_inputs_6_58_port, shift_in(57) => 
                           positive_inputs_6_57_port, shift_in(56) => 
                           positive_inputs_6_56_port, shift_in(55) => 
                           positive_inputs_6_55_port, shift_in(54) => 
                           positive_inputs_6_54_port, shift_in(53) => 
                           positive_inputs_6_53_port, shift_in(52) => 
                           positive_inputs_6_52_port, shift_in(51) => 
                           positive_inputs_6_51_port, shift_in(50) => 
                           positive_inputs_6_50_port, shift_in(49) => 
                           positive_inputs_6_49_port, shift_in(48) => 
                           positive_inputs_6_48_port, shift_in(47) => 
                           positive_inputs_6_47_port, shift_in(46) => 
                           positive_inputs_6_46_port, shift_in(45) => 
                           positive_inputs_6_45_port, shift_in(44) => 
                           positive_inputs_6_44_port, shift_in(43) => 
                           positive_inputs_6_43_port, shift_in(42) => 
                           positive_inputs_6_42_port, shift_in(41) => 
                           positive_inputs_6_41_port, shift_in(40) => 
                           positive_inputs_6_40_port, shift_in(39) => n53, 
                           shift_in(38) => positive_inputs_6_38_port, 
                           shift_in(37) => positive_inputs_6_37_port, 
                           shift_in(36) => positive_inputs_6_36_port, 
                           shift_in(35) => positive_inputs_6_35_port, 
                           shift_in(34) => positive_inputs_6_34_port, 
                           shift_in(33) => positive_inputs_6_33_port, 
                           shift_in(32) => positive_inputs_6_32_port, 
                           shift_in(31) => positive_inputs_6_31_port, 
                           shift_in(30) => positive_inputs_6_30_port, 
                           shift_in(29) => positive_inputs_6_29_port, 
                           shift_in(28) => positive_inputs_6_28_port, 
                           shift_in(27) => positive_inputs_6_27_port, 
                           shift_in(26) => positive_inputs_6_26_port, 
                           shift_in(25) => positive_inputs_6_25_port, 
                           shift_in(24) => positive_inputs_6_24_port, 
                           shift_in(23) => positive_inputs_6_23_port, 
                           shift_in(22) => positive_inputs_6_22_port, 
                           shift_in(21) => positive_inputs_6_21_port, 
                           shift_in(20) => positive_inputs_6_20_port, 
                           shift_in(19) => positive_inputs_6_19_port, 
                           shift_in(18) => positive_inputs_6_18_port, 
                           shift_in(17) => positive_inputs_6_17_port, 
                           shift_in(16) => positive_inputs_6_16_port, 
                           shift_in(15) => positive_inputs_6_15_port, 
                           shift_in(14) => positive_inputs_6_14_port, 
                           shift_in(13) => positive_inputs_6_13_port, 
                           shift_in(12) => positive_inputs_6_12_port, 
                           shift_in(11) => positive_inputs_6_11_port, 
                           shift_in(10) => positive_inputs_6_10_port, 
                           shift_in(9) => positive_inputs_6_9_port, shift_in(8)
                           => positive_inputs_6_8_port, shift_in(7) => 
                           positive_inputs_6_7_port, shift_in(6) => 
                           positive_inputs_6_6_port, shift_in(5) => 
                           positive_inputs_6_5_port, shift_in(4) => 
                           positive_inputs_6_4_port, shift_in(3) => 
                           positive_inputs_6_3_port, shift_in(2) => 
                           positive_inputs_6_2_port, shift_in(1) => 
                           positive_inputs_6_1_port, shift_in(0) => n9, 
                           shift_out(63) => positive_inputs_7_63_port, 
                           shift_out(62) => positive_inputs_7_62_port, 
                           shift_out(61) => positive_inputs_7_61_port, 
                           shift_out(60) => positive_inputs_7_60_port, 
                           shift_out(59) => positive_inputs_7_59_port, 
                           shift_out(58) => positive_inputs_7_58_port, 
                           shift_out(57) => positive_inputs_7_57_port, 
                           shift_out(56) => positive_inputs_7_56_port, 
                           shift_out(55) => positive_inputs_7_55_port, 
                           shift_out(54) => positive_inputs_7_54_port, 
                           shift_out(53) => positive_inputs_7_53_port, 
                           shift_out(52) => positive_inputs_7_52_port, 
                           shift_out(51) => positive_inputs_7_51_port, 
                           shift_out(50) => positive_inputs_7_50_port, 
                           shift_out(49) => positive_inputs_7_49_port, 
                           shift_out(48) => positive_inputs_7_48_port, 
                           shift_out(47) => positive_inputs_7_47_port, 
                           shift_out(46) => positive_inputs_7_46_port, 
                           shift_out(45) => positive_inputs_7_45_port, 
                           shift_out(44) => positive_inputs_7_44_port, 
                           shift_out(43) => positive_inputs_7_43_port, 
                           shift_out(42) => positive_inputs_7_42_port, 
                           shift_out(41) => positive_inputs_7_41_port, 
                           shift_out(40) => positive_inputs_7_40_port, 
                           shift_out(39) => positive_inputs_7_39_port, 
                           shift_out(38) => positive_inputs_7_38_port, 
                           shift_out(37) => positive_inputs_7_37_port, 
                           shift_out(36) => positive_inputs_7_36_port, 
                           shift_out(35) => positive_inputs_7_35_port, 
                           shift_out(34) => positive_inputs_7_34_port, 
                           shift_out(33) => positive_inputs_7_33_port, 
                           shift_out(32) => positive_inputs_7_32_port, 
                           shift_out(31) => positive_inputs_7_31_port, 
                           shift_out(30) => positive_inputs_7_30_port, 
                           shift_out(29) => positive_inputs_7_29_port, 
                           shift_out(28) => positive_inputs_7_28_port, 
                           shift_out(27) => positive_inputs_7_27_port, 
                           shift_out(26) => positive_inputs_7_26_port, 
                           shift_out(25) => positive_inputs_7_25_port, 
                           shift_out(24) => positive_inputs_7_24_port, 
                           shift_out(23) => positive_inputs_7_23_port, 
                           shift_out(22) => positive_inputs_7_22_port, 
                           shift_out(21) => positive_inputs_7_21_port, 
                           shift_out(20) => positive_inputs_7_20_port, 
                           shift_out(19) => positive_inputs_7_19_port, 
                           shift_out(18) => positive_inputs_7_18_port, 
                           shift_out(17) => positive_inputs_7_17_port, 
                           shift_out(16) => positive_inputs_7_16_port, 
                           shift_out(15) => positive_inputs_7_15_port, 
                           shift_out(14) => positive_inputs_7_14_port, 
                           shift_out(13) => positive_inputs_7_13_port, 
                           shift_out(12) => positive_inputs_7_12_port, 
                           shift_out(11) => positive_inputs_7_11_port, 
                           shift_out(10) => positive_inputs_7_10_port, 
                           shift_out(9) => positive_inputs_7_9_port, 
                           shift_out(8) => positive_inputs_7_8_port, 
                           shift_out(7) => positive_inputs_7_7_port, 
                           shift_out(6) => positive_inputs_7_6_port, 
                           shift_out(5) => positive_inputs_7_5_port, 
                           shift_out(4) => positive_inputs_7_4_port, 
                           shift_out(3) => positive_inputs_7_3_port, 
                           shift_out(2) => positive_inputs_7_2_port, 
                           shift_out(1) => positive_inputs_7_1_port, 
                           shift_out(0) => n_1007);
   shifted_pos_8 : leftshifter_NbitShifter64_56 port map( shift_in(63) => 
                           positive_inputs_7_63_port, shift_in(62) => 
                           positive_inputs_7_62_port, shift_in(61) => 
                           positive_inputs_7_61_port, shift_in(60) => 
                           positive_inputs_7_60_port, shift_in(59) => 
                           positive_inputs_7_59_port, shift_in(58) => 
                           positive_inputs_7_58_port, shift_in(57) => 
                           positive_inputs_7_57_port, shift_in(56) => 
                           positive_inputs_7_56_port, shift_in(55) => 
                           positive_inputs_7_55_port, shift_in(54) => 
                           positive_inputs_7_54_port, shift_in(53) => 
                           positive_inputs_7_53_port, shift_in(52) => 
                           positive_inputs_7_52_port, shift_in(51) => 
                           positive_inputs_7_51_port, shift_in(50) => 
                           positive_inputs_7_50_port, shift_in(49) => 
                           positive_inputs_7_49_port, shift_in(48) => n66, 
                           shift_in(47) => positive_inputs_7_47_port, 
                           shift_in(46) => positive_inputs_7_46_port, 
                           shift_in(45) => positive_inputs_7_45_port, 
                           shift_in(44) => positive_inputs_7_44_port, 
                           shift_in(43) => positive_inputs_7_43_port, 
                           shift_in(42) => positive_inputs_7_42_port, 
                           shift_in(41) => positive_inputs_7_41_port, 
                           shift_in(40) => positive_inputs_7_40_port, 
                           shift_in(39) => n52, shift_in(38) => n51, 
                           shift_in(37) => n214, shift_in(36) => n212, 
                           shift_in(35) => n210, shift_in(34) => n208, 
                           shift_in(33) => n206, shift_in(32) => n204, 
                           shift_in(31) => n202, shift_in(30) => n200, 
                           shift_in(29) => n198, shift_in(28) => n196, 
                           shift_in(27) => n194, shift_in(26) => n192, 
                           shift_in(25) => n190, shift_in(24) => n188, 
                           shift_in(23) => n186, shift_in(22) => n184, 
                           shift_in(21) => n182, shift_in(20) => n180, 
                           shift_in(19) => n178, shift_in(18) => n176, 
                           shift_in(17) => n174, shift_in(16) => n172, 
                           shift_in(15) => n170, shift_in(14) => n168, 
                           shift_in(13) => n166, shift_in(12) => n164, 
                           shift_in(11) => n162, shift_in(10) => n160, 
                           shift_in(9) => n158, shift_in(8) => n156, 
                           shift_in(7) => n154, shift_in(6) => 
                           positive_inputs_7_6_port, shift_in(5) => 
                           positive_inputs_7_5_port, shift_in(4) => 
                           positive_inputs_7_4_port, shift_in(3) => 
                           positive_inputs_7_3_port, shift_in(2) => 
                           positive_inputs_7_2_port, shift_in(1) => 
                           positive_inputs_7_1_port, shift_in(0) => n9, 
                           shift_out(63) => positive_inputs_8_63_port, 
                           shift_out(62) => positive_inputs_8_62_port, 
                           shift_out(61) => positive_inputs_8_61_port, 
                           shift_out(60) => positive_inputs_8_60_port, 
                           shift_out(59) => positive_inputs_8_59_port, 
                           shift_out(58) => positive_inputs_8_58_port, 
                           shift_out(57) => positive_inputs_8_57_port, 
                           shift_out(56) => positive_inputs_8_56_port, 
                           shift_out(55) => positive_inputs_8_55_port, 
                           shift_out(54) => positive_inputs_8_54_port, 
                           shift_out(53) => positive_inputs_8_53_port, 
                           shift_out(52) => positive_inputs_8_52_port, 
                           shift_out(51) => positive_inputs_8_51_port, 
                           shift_out(50) => positive_inputs_8_50_port, 
                           shift_out(49) => positive_inputs_8_49_port, 
                           shift_out(48) => positive_inputs_8_48_port, 
                           shift_out(47) => positive_inputs_8_47_port, 
                           shift_out(46) => positive_inputs_8_46_port, 
                           shift_out(45) => positive_inputs_8_45_port, 
                           shift_out(44) => positive_inputs_8_44_port, 
                           shift_out(43) => positive_inputs_8_43_port, 
                           shift_out(42) => positive_inputs_8_42_port, 
                           shift_out(41) => positive_inputs_8_41_port, 
                           shift_out(40) => positive_inputs_8_40_port, 
                           shift_out(39) => positive_inputs_8_39_port, 
                           shift_out(38) => positive_inputs_8_38_port, 
                           shift_out(37) => positive_inputs_8_37_port, 
                           shift_out(36) => positive_inputs_8_36_port, 
                           shift_out(35) => positive_inputs_8_35_port, 
                           shift_out(34) => positive_inputs_8_34_port, 
                           shift_out(33) => positive_inputs_8_33_port, 
                           shift_out(32) => positive_inputs_8_32_port, 
                           shift_out(31) => positive_inputs_8_31_port, 
                           shift_out(30) => positive_inputs_8_30_port, 
                           shift_out(29) => positive_inputs_8_29_port, 
                           shift_out(28) => positive_inputs_8_28_port, 
                           shift_out(27) => positive_inputs_8_27_port, 
                           shift_out(26) => positive_inputs_8_26_port, 
                           shift_out(25) => positive_inputs_8_25_port, 
                           shift_out(24) => positive_inputs_8_24_port, 
                           shift_out(23) => positive_inputs_8_23_port, 
                           shift_out(22) => positive_inputs_8_22_port, 
                           shift_out(21) => positive_inputs_8_21_port, 
                           shift_out(20) => positive_inputs_8_20_port, 
                           shift_out(19) => positive_inputs_8_19_port, 
                           shift_out(18) => positive_inputs_8_18_port, 
                           shift_out(17) => positive_inputs_8_17_port, 
                           shift_out(16) => positive_inputs_8_16_port, 
                           shift_out(15) => positive_inputs_8_15_port, 
                           shift_out(14) => positive_inputs_8_14_port, 
                           shift_out(13) => positive_inputs_8_13_port, 
                           shift_out(12) => positive_inputs_8_12_port, 
                           shift_out(11) => positive_inputs_8_11_port, 
                           shift_out(10) => positive_inputs_8_10_port, 
                           shift_out(9) => positive_inputs_8_9_port, 
                           shift_out(8) => positive_inputs_8_8_port, 
                           shift_out(7) => positive_inputs_8_7_port, 
                           shift_out(6) => positive_inputs_8_6_port, 
                           shift_out(5) => positive_inputs_8_5_port, 
                           shift_out(4) => positive_inputs_8_4_port, 
                           shift_out(3) => positive_inputs_8_3_port, 
                           shift_out(2) => positive_inputs_8_2_port, 
                           shift_out(1) => positive_inputs_8_1_port, 
                           shift_out(0) => n_1008);
   shifted_pos_9 : leftshifter_NbitShifter64_55 port map( shift_in(63) => 
                           positive_inputs_8_63_port, shift_in(62) => 
                           positive_inputs_8_62_port, shift_in(61) => 
                           positive_inputs_8_61_port, shift_in(60) => 
                           positive_inputs_8_60_port, shift_in(59) => 
                           positive_inputs_8_59_port, shift_in(58) => 
                           positive_inputs_8_58_port, shift_in(57) => 
                           positive_inputs_8_57_port, shift_in(56) => 
                           positive_inputs_8_56_port, shift_in(55) => 
                           positive_inputs_8_55_port, shift_in(54) => 
                           positive_inputs_8_54_port, shift_in(53) => 
                           positive_inputs_8_53_port, shift_in(52) => 
                           positive_inputs_8_52_port, shift_in(51) => 
                           positive_inputs_8_51_port, shift_in(50) => 
                           positive_inputs_8_50_port, shift_in(49) => 
                           positive_inputs_8_49_port, shift_in(48) => n65, 
                           shift_in(47) => positive_inputs_8_47_port, 
                           shift_in(46) => positive_inputs_8_46_port, 
                           shift_in(45) => positive_inputs_8_45_port, 
                           shift_in(44) => positive_inputs_8_44_port, 
                           shift_in(43) => positive_inputs_8_43_port, 
                           shift_in(42) => positive_inputs_8_42_port, 
                           shift_in(41) => positive_inputs_8_41_port, 
                           shift_in(40) => positive_inputs_8_40_port, 
                           shift_in(39) => positive_inputs_8_39_port, 
                           shift_in(38) => positive_inputs_8_38_port, 
                           shift_in(37) => positive_inputs_8_37_port, 
                           shift_in(36) => positive_inputs_8_36_port, 
                           shift_in(35) => positive_inputs_8_35_port, 
                           shift_in(34) => positive_inputs_8_34_port, 
                           shift_in(33) => positive_inputs_8_33_port, 
                           shift_in(32) => positive_inputs_8_32_port, 
                           shift_in(31) => positive_inputs_8_31_port, 
                           shift_in(30) => positive_inputs_8_30_port, 
                           shift_in(29) => positive_inputs_8_29_port, 
                           shift_in(28) => positive_inputs_8_28_port, 
                           shift_in(27) => positive_inputs_8_27_port, 
                           shift_in(26) => positive_inputs_8_26_port, 
                           shift_in(25) => positive_inputs_8_25_port, 
                           shift_in(24) => positive_inputs_8_24_port, 
                           shift_in(23) => positive_inputs_8_23_port, 
                           shift_in(22) => positive_inputs_8_22_port, 
                           shift_in(21) => positive_inputs_8_21_port, 
                           shift_in(20) => positive_inputs_8_20_port, 
                           shift_in(19) => positive_inputs_8_19_port, 
                           shift_in(18) => positive_inputs_8_18_port, 
                           shift_in(17) => positive_inputs_8_17_port, 
                           shift_in(16) => positive_inputs_8_16_port, 
                           shift_in(15) => positive_inputs_8_15_port, 
                           shift_in(14) => positive_inputs_8_14_port, 
                           shift_in(13) => positive_inputs_8_13_port, 
                           shift_in(12) => positive_inputs_8_12_port, 
                           shift_in(11) => positive_inputs_8_11_port, 
                           shift_in(10) => positive_inputs_8_10_port, 
                           shift_in(9) => positive_inputs_8_9_port, shift_in(8)
                           => positive_inputs_8_8_port, shift_in(7) => 
                           positive_inputs_8_7_port, shift_in(6) => 
                           positive_inputs_8_6_port, shift_in(5) => 
                           positive_inputs_8_5_port, shift_in(4) => 
                           positive_inputs_8_4_port, shift_in(3) => 
                           positive_inputs_8_3_port, shift_in(2) => 
                           positive_inputs_8_2_port, shift_in(1) => 
                           positive_inputs_8_1_port, shift_in(0) => n9, 
                           shift_out(63) => positive_inputs_9_63_port, 
                           shift_out(62) => positive_inputs_9_62_port, 
                           shift_out(61) => positive_inputs_9_61_port, 
                           shift_out(60) => positive_inputs_9_60_port, 
                           shift_out(59) => positive_inputs_9_59_port, 
                           shift_out(58) => positive_inputs_9_58_port, 
                           shift_out(57) => positive_inputs_9_57_port, 
                           shift_out(56) => positive_inputs_9_56_port, 
                           shift_out(55) => positive_inputs_9_55_port, 
                           shift_out(54) => positive_inputs_9_54_port, 
                           shift_out(53) => positive_inputs_9_53_port, 
                           shift_out(52) => positive_inputs_9_52_port, 
                           shift_out(51) => positive_inputs_9_51_port, 
                           shift_out(50) => positive_inputs_9_50_port, 
                           shift_out(49) => positive_inputs_9_49_port, 
                           shift_out(48) => positive_inputs_9_48_port, 
                           shift_out(47) => positive_inputs_9_47_port, 
                           shift_out(46) => positive_inputs_9_46_port, 
                           shift_out(45) => positive_inputs_9_45_port, 
                           shift_out(44) => positive_inputs_9_44_port, 
                           shift_out(43) => positive_inputs_9_43_port, 
                           shift_out(42) => positive_inputs_9_42_port, 
                           shift_out(41) => positive_inputs_9_41_port, 
                           shift_out(40) => positive_inputs_9_40_port, 
                           shift_out(39) => positive_inputs_9_39_port, 
                           shift_out(38) => positive_inputs_9_38_port, 
                           shift_out(37) => positive_inputs_9_37_port, 
                           shift_out(36) => positive_inputs_9_36_port, 
                           shift_out(35) => positive_inputs_9_35_port, 
                           shift_out(34) => positive_inputs_9_34_port, 
                           shift_out(33) => positive_inputs_9_33_port, 
                           shift_out(32) => positive_inputs_9_32_port, 
                           shift_out(31) => positive_inputs_9_31_port, 
                           shift_out(30) => positive_inputs_9_30_port, 
                           shift_out(29) => positive_inputs_9_29_port, 
                           shift_out(28) => positive_inputs_9_28_port, 
                           shift_out(27) => positive_inputs_9_27_port, 
                           shift_out(26) => positive_inputs_9_26_port, 
                           shift_out(25) => positive_inputs_9_25_port, 
                           shift_out(24) => positive_inputs_9_24_port, 
                           shift_out(23) => positive_inputs_9_23_port, 
                           shift_out(22) => positive_inputs_9_22_port, 
                           shift_out(21) => positive_inputs_9_21_port, 
                           shift_out(20) => positive_inputs_9_20_port, 
                           shift_out(19) => positive_inputs_9_19_port, 
                           shift_out(18) => positive_inputs_9_18_port, 
                           shift_out(17) => positive_inputs_9_17_port, 
                           shift_out(16) => positive_inputs_9_16_port, 
                           shift_out(15) => positive_inputs_9_15_port, 
                           shift_out(14) => positive_inputs_9_14_port, 
                           shift_out(13) => positive_inputs_9_13_port, 
                           shift_out(12) => positive_inputs_9_12_port, 
                           shift_out(11) => positive_inputs_9_11_port, 
                           shift_out(10) => positive_inputs_9_10_port, 
                           shift_out(9) => positive_inputs_9_9_port, 
                           shift_out(8) => positive_inputs_9_8_port, 
                           shift_out(7) => positive_inputs_9_7_port, 
                           shift_out(6) => positive_inputs_9_6_port, 
                           shift_out(5) => positive_inputs_9_5_port, 
                           shift_out(4) => positive_inputs_9_4_port, 
                           shift_out(3) => positive_inputs_9_3_port, 
                           shift_out(2) => positive_inputs_9_2_port, 
                           shift_out(1) => positive_inputs_9_1_port, 
                           shift_out(0) => n_1009);
   shifted_pos_10 : leftshifter_NbitShifter64_54 port map( shift_in(63) => 
                           positive_inputs_9_63_port, shift_in(62) => 
                           positive_inputs_9_62_port, shift_in(61) => 
                           positive_inputs_9_61_port, shift_in(60) => 
                           positive_inputs_9_60_port, shift_in(59) => 
                           positive_inputs_9_59_port, shift_in(58) => 
                           positive_inputs_9_58_port, shift_in(57) => 
                           positive_inputs_9_57_port, shift_in(56) => 
                           positive_inputs_9_56_port, shift_in(55) => 
                           positive_inputs_9_55_port, shift_in(54) => 
                           positive_inputs_9_54_port, shift_in(53) => 
                           positive_inputs_9_53_port, shift_in(52) => 
                           positive_inputs_9_52_port, shift_in(51) => 
                           positive_inputs_9_51_port, shift_in(50) => 
                           positive_inputs_9_50_port, shift_in(49) => 
                           positive_inputs_9_49_port, shift_in(48) => n64, 
                           shift_in(47) => positive_inputs_9_47_port, 
                           shift_in(46) => positive_inputs_9_46_port, 
                           shift_in(45) => positive_inputs_9_45_port, 
                           shift_in(44) => positive_inputs_9_44_port, 
                           shift_in(43) => positive_inputs_9_43_port, 
                           shift_in(42) => positive_inputs_9_42_port, 
                           shift_in(41) => positive_inputs_9_41_port, 
                           shift_in(40) => positive_inputs_9_40_port, 
                           shift_in(39) => positive_inputs_9_39_port, 
                           shift_in(38) => positive_inputs_9_38_port, 
                           shift_in(37) => positive_inputs_9_37_port, 
                           shift_in(36) => positive_inputs_9_36_port, 
                           shift_in(35) => positive_inputs_9_35_port, 
                           shift_in(34) => positive_inputs_9_34_port, 
                           shift_in(33) => positive_inputs_9_33_port, 
                           shift_in(32) => positive_inputs_9_32_port, 
                           shift_in(31) => positive_inputs_9_31_port, 
                           shift_in(30) => positive_inputs_9_30_port, 
                           shift_in(29) => positive_inputs_9_29_port, 
                           shift_in(28) => positive_inputs_9_28_port, 
                           shift_in(27) => positive_inputs_9_27_port, 
                           shift_in(26) => positive_inputs_9_26_port, 
                           shift_in(25) => positive_inputs_9_25_port, 
                           shift_in(24) => positive_inputs_9_24_port, 
                           shift_in(23) => positive_inputs_9_23_port, 
                           shift_in(22) => positive_inputs_9_22_port, 
                           shift_in(21) => positive_inputs_9_21_port, 
                           shift_in(20) => positive_inputs_9_20_port, 
                           shift_in(19) => positive_inputs_9_19_port, 
                           shift_in(18) => positive_inputs_9_18_port, 
                           shift_in(17) => positive_inputs_9_17_port, 
                           shift_in(16) => positive_inputs_9_16_port, 
                           shift_in(15) => positive_inputs_9_15_port, 
                           shift_in(14) => positive_inputs_9_14_port, 
                           shift_in(13) => positive_inputs_9_13_port, 
                           shift_in(12) => positive_inputs_9_12_port, 
                           shift_in(11) => positive_inputs_9_11_port, 
                           shift_in(10) => positive_inputs_9_10_port, 
                           shift_in(9) => positive_inputs_9_9_port, shift_in(8)
                           => positive_inputs_9_8_port, shift_in(7) => 
                           positive_inputs_9_7_port, shift_in(6) => 
                           positive_inputs_9_6_port, shift_in(5) => 
                           positive_inputs_9_5_port, shift_in(4) => 
                           positive_inputs_9_4_port, shift_in(3) => 
                           positive_inputs_9_3_port, shift_in(2) => 
                           positive_inputs_9_2_port, shift_in(1) => 
                           positive_inputs_9_1_port, shift_in(0) => n9, 
                           shift_out(63) => positive_inputs_10_63_port, 
                           shift_out(62) => positive_inputs_10_62_port, 
                           shift_out(61) => positive_inputs_10_61_port, 
                           shift_out(60) => positive_inputs_10_60_port, 
                           shift_out(59) => positive_inputs_10_59_port, 
                           shift_out(58) => positive_inputs_10_58_port, 
                           shift_out(57) => positive_inputs_10_57_port, 
                           shift_out(56) => positive_inputs_10_56_port, 
                           shift_out(55) => positive_inputs_10_55_port, 
                           shift_out(54) => positive_inputs_10_54_port, 
                           shift_out(53) => positive_inputs_10_53_port, 
                           shift_out(52) => positive_inputs_10_52_port, 
                           shift_out(51) => positive_inputs_10_51_port, 
                           shift_out(50) => positive_inputs_10_50_port, 
                           shift_out(49) => positive_inputs_10_49_port, 
                           shift_out(48) => positive_inputs_10_48_port, 
                           shift_out(47) => positive_inputs_10_47_port, 
                           shift_out(46) => positive_inputs_10_46_port, 
                           shift_out(45) => positive_inputs_10_45_port, 
                           shift_out(44) => positive_inputs_10_44_port, 
                           shift_out(43) => positive_inputs_10_43_port, 
                           shift_out(42) => positive_inputs_10_42_port, 
                           shift_out(41) => positive_inputs_10_41_port, 
                           shift_out(40) => positive_inputs_10_40_port, 
                           shift_out(39) => positive_inputs_10_39_port, 
                           shift_out(38) => positive_inputs_10_38_port, 
                           shift_out(37) => positive_inputs_10_37_port, 
                           shift_out(36) => positive_inputs_10_36_port, 
                           shift_out(35) => positive_inputs_10_35_port, 
                           shift_out(34) => positive_inputs_10_34_port, 
                           shift_out(33) => positive_inputs_10_33_port, 
                           shift_out(32) => positive_inputs_10_32_port, 
                           shift_out(31) => positive_inputs_10_31_port, 
                           shift_out(30) => positive_inputs_10_30_port, 
                           shift_out(29) => positive_inputs_10_29_port, 
                           shift_out(28) => positive_inputs_10_28_port, 
                           shift_out(27) => positive_inputs_10_27_port, 
                           shift_out(26) => positive_inputs_10_26_port, 
                           shift_out(25) => positive_inputs_10_25_port, 
                           shift_out(24) => positive_inputs_10_24_port, 
                           shift_out(23) => positive_inputs_10_23_port, 
                           shift_out(22) => positive_inputs_10_22_port, 
                           shift_out(21) => positive_inputs_10_21_port, 
                           shift_out(20) => positive_inputs_10_20_port, 
                           shift_out(19) => positive_inputs_10_19_port, 
                           shift_out(18) => positive_inputs_10_18_port, 
                           shift_out(17) => positive_inputs_10_17_port, 
                           shift_out(16) => positive_inputs_10_16_port, 
                           shift_out(15) => positive_inputs_10_15_port, 
                           shift_out(14) => positive_inputs_10_14_port, 
                           shift_out(13) => positive_inputs_10_13_port, 
                           shift_out(12) => positive_inputs_10_12_port, 
                           shift_out(11) => positive_inputs_10_11_port, 
                           shift_out(10) => positive_inputs_10_10_port, 
                           shift_out(9) => positive_inputs_10_9_port, 
                           shift_out(8) => positive_inputs_10_8_port, 
                           shift_out(7) => positive_inputs_10_7_port, 
                           shift_out(6) => positive_inputs_10_6_port, 
                           shift_out(5) => positive_inputs_10_5_port, 
                           shift_out(4) => positive_inputs_10_4_port, 
                           shift_out(3) => positive_inputs_10_3_port, 
                           shift_out(2) => positive_inputs_10_2_port, 
                           shift_out(1) => positive_inputs_10_1_port, 
                           shift_out(0) => n_1010);
   shifted_pos_11 : leftshifter_NbitShifter64_53 port map( shift_in(63) => 
                           positive_inputs_10_63_port, shift_in(62) => 
                           positive_inputs_10_62_port, shift_in(61) => 
                           positive_inputs_10_61_port, shift_in(60) => 
                           positive_inputs_10_60_port, shift_in(59) => 
                           positive_inputs_10_59_port, shift_in(58) => 
                           positive_inputs_10_58_port, shift_in(57) => 
                           positive_inputs_10_57_port, shift_in(56) => 
                           positive_inputs_10_56_port, shift_in(55) => 
                           positive_inputs_10_55_port, shift_in(54) => 
                           positive_inputs_10_54_port, shift_in(53) => 
                           positive_inputs_10_53_port, shift_in(52) => 
                           positive_inputs_10_52_port, shift_in(51) => 
                           positive_inputs_10_51_port, shift_in(50) => 
                           positive_inputs_10_50_port, shift_in(49) => 
                           positive_inputs_10_49_port, shift_in(48) => n63, 
                           shift_in(47) => positive_inputs_10_47_port, 
                           shift_in(46) => positive_inputs_10_46_port, 
                           shift_in(45) => positive_inputs_10_45_port, 
                           shift_in(44) => positive_inputs_10_44_port, 
                           shift_in(43) => positive_inputs_10_43_port, 
                           shift_in(42) => positive_inputs_10_42_port, 
                           shift_in(41) => positive_inputs_10_41_port, 
                           shift_in(40) => positive_inputs_10_40_port, 
                           shift_in(39) => positive_inputs_10_39_port, 
                           shift_in(38) => positive_inputs_10_38_port, 
                           shift_in(37) => positive_inputs_10_37_port, 
                           shift_in(36) => positive_inputs_10_36_port, 
                           shift_in(35) => positive_inputs_10_35_port, 
                           shift_in(34) => positive_inputs_10_34_port, 
                           shift_in(33) => positive_inputs_10_33_port, 
                           shift_in(32) => positive_inputs_10_32_port, 
                           shift_in(31) => positive_inputs_10_31_port, 
                           shift_in(30) => positive_inputs_10_30_port, 
                           shift_in(29) => positive_inputs_10_29_port, 
                           shift_in(28) => positive_inputs_10_28_port, 
                           shift_in(27) => positive_inputs_10_27_port, 
                           shift_in(26) => positive_inputs_10_26_port, 
                           shift_in(25) => positive_inputs_10_25_port, 
                           shift_in(24) => positive_inputs_10_24_port, 
                           shift_in(23) => positive_inputs_10_23_port, 
                           shift_in(22) => positive_inputs_10_22_port, 
                           shift_in(21) => positive_inputs_10_21_port, 
                           shift_in(20) => positive_inputs_10_20_port, 
                           shift_in(19) => positive_inputs_10_19_port, 
                           shift_in(18) => positive_inputs_10_18_port, 
                           shift_in(17) => positive_inputs_10_17_port, 
                           shift_in(16) => positive_inputs_10_16_port, 
                           shift_in(15) => positive_inputs_10_15_port, 
                           shift_in(14) => positive_inputs_10_14_port, 
                           shift_in(13) => positive_inputs_10_13_port, 
                           shift_in(12) => positive_inputs_10_12_port, 
                           shift_in(11) => positive_inputs_10_11_port, 
                           shift_in(10) => positive_inputs_10_10_port, 
                           shift_in(9) => positive_inputs_10_9_port, 
                           shift_in(8) => positive_inputs_10_8_port, 
                           shift_in(7) => positive_inputs_10_7_port, 
                           shift_in(6) => positive_inputs_10_6_port, 
                           shift_in(5) => positive_inputs_10_5_port, 
                           shift_in(4) => positive_inputs_10_4_port, 
                           shift_in(3) => positive_inputs_10_3_port, 
                           shift_in(2) => positive_inputs_10_2_port, 
                           shift_in(1) => positive_inputs_10_1_port, 
                           shift_in(0) => n9, shift_out(63) => 
                           positive_inputs_11_63_port, shift_out(62) => 
                           positive_inputs_11_62_port, shift_out(61) => 
                           positive_inputs_11_61_port, shift_out(60) => 
                           positive_inputs_11_60_port, shift_out(59) => 
                           positive_inputs_11_59_port, shift_out(58) => 
                           positive_inputs_11_58_port, shift_out(57) => 
                           positive_inputs_11_57_port, shift_out(56) => 
                           positive_inputs_11_56_port, shift_out(55) => 
                           positive_inputs_11_55_port, shift_out(54) => 
                           positive_inputs_11_54_port, shift_out(53) => 
                           positive_inputs_11_53_port, shift_out(52) => 
                           positive_inputs_11_52_port, shift_out(51) => 
                           positive_inputs_11_51_port, shift_out(50) => 
                           positive_inputs_11_50_port, shift_out(49) => 
                           positive_inputs_11_49_port, shift_out(48) => 
                           positive_inputs_11_48_port, shift_out(47) => 
                           positive_inputs_11_47_port, shift_out(46) => 
                           positive_inputs_11_46_port, shift_out(45) => 
                           positive_inputs_11_45_port, shift_out(44) => 
                           positive_inputs_11_44_port, shift_out(43) => 
                           positive_inputs_11_43_port, shift_out(42) => 
                           positive_inputs_11_42_port, shift_out(41) => 
                           positive_inputs_11_41_port, shift_out(40) => 
                           positive_inputs_11_40_port, shift_out(39) => 
                           positive_inputs_11_39_port, shift_out(38) => 
                           positive_inputs_11_38_port, shift_out(37) => 
                           positive_inputs_11_37_port, shift_out(36) => 
                           positive_inputs_11_36_port, shift_out(35) => 
                           positive_inputs_11_35_port, shift_out(34) => 
                           positive_inputs_11_34_port, shift_out(33) => 
                           positive_inputs_11_33_port, shift_out(32) => 
                           positive_inputs_11_32_port, shift_out(31) => 
                           positive_inputs_11_31_port, shift_out(30) => 
                           positive_inputs_11_30_port, shift_out(29) => 
                           positive_inputs_11_29_port, shift_out(28) => 
                           positive_inputs_11_28_port, shift_out(27) => 
                           positive_inputs_11_27_port, shift_out(26) => 
                           positive_inputs_11_26_port, shift_out(25) => 
                           positive_inputs_11_25_port, shift_out(24) => 
                           positive_inputs_11_24_port, shift_out(23) => 
                           positive_inputs_11_23_port, shift_out(22) => 
                           positive_inputs_11_22_port, shift_out(21) => 
                           positive_inputs_11_21_port, shift_out(20) => 
                           positive_inputs_11_20_port, shift_out(19) => 
                           positive_inputs_11_19_port, shift_out(18) => 
                           positive_inputs_11_18_port, shift_out(17) => 
                           positive_inputs_11_17_port, shift_out(16) => 
                           positive_inputs_11_16_port, shift_out(15) => 
                           positive_inputs_11_15_port, shift_out(14) => 
                           positive_inputs_11_14_port, shift_out(13) => 
                           positive_inputs_11_13_port, shift_out(12) => 
                           positive_inputs_11_12_port, shift_out(11) => 
                           positive_inputs_11_11_port, shift_out(10) => 
                           positive_inputs_11_10_port, shift_out(9) => 
                           positive_inputs_11_9_port, shift_out(8) => 
                           positive_inputs_11_8_port, shift_out(7) => 
                           positive_inputs_11_7_port, shift_out(6) => 
                           positive_inputs_11_6_port, shift_out(5) => 
                           positive_inputs_11_5_port, shift_out(4) => 
                           positive_inputs_11_4_port, shift_out(3) => 
                           positive_inputs_11_3_port, shift_out(2) => 
                           positive_inputs_11_2_port, shift_out(1) => 
                           positive_inputs_11_1_port, shift_out(0) => n_1011);
   shifted_pos_12 : leftshifter_NbitShifter64_52 port map( shift_in(63) => 
                           positive_inputs_11_63_port, shift_in(62) => 
                           positive_inputs_11_62_port, shift_in(61) => 
                           positive_inputs_11_61_port, shift_in(60) => 
                           positive_inputs_11_60_port, shift_in(59) => 
                           positive_inputs_11_59_port, shift_in(58) => 
                           positive_inputs_11_58_port, shift_in(57) => 
                           positive_inputs_11_57_port, shift_in(56) => 
                           positive_inputs_11_56_port, shift_in(55) => 
                           positive_inputs_11_55_port, shift_in(54) => 
                           positive_inputs_11_54_port, shift_in(53) => 
                           positive_inputs_11_53_port, shift_in(52) => 
                           positive_inputs_11_52_port, shift_in(51) => 
                           positive_inputs_11_51_port, shift_in(50) => 
                           positive_inputs_11_50_port, shift_in(49) => 
                           positive_inputs_11_49_port, shift_in(48) => n62, 
                           shift_in(47) => positive_inputs_11_47_port, 
                           shift_in(46) => positive_inputs_11_46_port, 
                           shift_in(45) => positive_inputs_11_45_port, 
                           shift_in(44) => positive_inputs_11_44_port, 
                           shift_in(43) => positive_inputs_11_43_port, 
                           shift_in(42) => positive_inputs_11_42_port, 
                           shift_in(41) => positive_inputs_11_41_port, 
                           shift_in(40) => positive_inputs_11_40_port, 
                           shift_in(39) => positive_inputs_11_39_port, 
                           shift_in(38) => positive_inputs_11_38_port, 
                           shift_in(37) => positive_inputs_11_37_port, 
                           shift_in(36) => positive_inputs_11_36_port, 
                           shift_in(35) => positive_inputs_11_35_port, 
                           shift_in(34) => positive_inputs_11_34_port, 
                           shift_in(33) => positive_inputs_11_33_port, 
                           shift_in(32) => positive_inputs_11_32_port, 
                           shift_in(31) => positive_inputs_11_31_port, 
                           shift_in(30) => positive_inputs_11_30_port, 
                           shift_in(29) => positive_inputs_11_29_port, 
                           shift_in(28) => positive_inputs_11_28_port, 
                           shift_in(27) => positive_inputs_11_27_port, 
                           shift_in(26) => positive_inputs_11_26_port, 
                           shift_in(25) => positive_inputs_11_25_port, 
                           shift_in(24) => positive_inputs_11_24_port, 
                           shift_in(23) => positive_inputs_11_23_port, 
                           shift_in(22) => positive_inputs_11_22_port, 
                           shift_in(21) => positive_inputs_11_21_port, 
                           shift_in(20) => positive_inputs_11_20_port, 
                           shift_in(19) => positive_inputs_11_19_port, 
                           shift_in(18) => positive_inputs_11_18_port, 
                           shift_in(17) => positive_inputs_11_17_port, 
                           shift_in(16) => positive_inputs_11_16_port, 
                           shift_in(15) => positive_inputs_11_15_port, 
                           shift_in(14) => positive_inputs_11_14_port, 
                           shift_in(13) => positive_inputs_11_13_port, 
                           shift_in(12) => positive_inputs_11_12_port, 
                           shift_in(11) => positive_inputs_11_11_port, 
                           shift_in(10) => positive_inputs_11_10_port, 
                           shift_in(9) => positive_inputs_11_9_port, 
                           shift_in(8) => positive_inputs_11_8_port, 
                           shift_in(7) => positive_inputs_11_7_port, 
                           shift_in(6) => positive_inputs_11_6_port, 
                           shift_in(5) => positive_inputs_11_5_port, 
                           shift_in(4) => positive_inputs_11_4_port, 
                           shift_in(3) => positive_inputs_11_3_port, 
                           shift_in(2) => positive_inputs_11_2_port, 
                           shift_in(1) => positive_inputs_11_1_port, 
                           shift_in(0) => n9, shift_out(63) => 
                           positive_inputs_12_63_port, shift_out(62) => 
                           positive_inputs_12_62_port, shift_out(61) => 
                           positive_inputs_12_61_port, shift_out(60) => 
                           positive_inputs_12_60_port, shift_out(59) => 
                           positive_inputs_12_59_port, shift_out(58) => 
                           positive_inputs_12_58_port, shift_out(57) => 
                           positive_inputs_12_57_port, shift_out(56) => 
                           positive_inputs_12_56_port, shift_out(55) => 
                           positive_inputs_12_55_port, shift_out(54) => 
                           positive_inputs_12_54_port, shift_out(53) => 
                           positive_inputs_12_53_port, shift_out(52) => 
                           positive_inputs_12_52_port, shift_out(51) => 
                           positive_inputs_12_51_port, shift_out(50) => 
                           positive_inputs_12_50_port, shift_out(49) => 
                           positive_inputs_12_49_port, shift_out(48) => 
                           positive_inputs_12_48_port, shift_out(47) => 
                           positive_inputs_12_47_port, shift_out(46) => 
                           positive_inputs_12_46_port, shift_out(45) => 
                           positive_inputs_12_45_port, shift_out(44) => 
                           positive_inputs_12_44_port, shift_out(43) => 
                           positive_inputs_12_43_port, shift_out(42) => 
                           positive_inputs_12_42_port, shift_out(41) => 
                           positive_inputs_12_41_port, shift_out(40) => 
                           positive_inputs_12_40_port, shift_out(39) => 
                           positive_inputs_12_39_port, shift_out(38) => 
                           positive_inputs_12_38_port, shift_out(37) => 
                           positive_inputs_12_37_port, shift_out(36) => 
                           positive_inputs_12_36_port, shift_out(35) => 
                           positive_inputs_12_35_port, shift_out(34) => 
                           positive_inputs_12_34_port, shift_out(33) => 
                           positive_inputs_12_33_port, shift_out(32) => 
                           positive_inputs_12_32_port, shift_out(31) => 
                           positive_inputs_12_31_port, shift_out(30) => 
                           positive_inputs_12_30_port, shift_out(29) => 
                           positive_inputs_12_29_port, shift_out(28) => 
                           positive_inputs_12_28_port, shift_out(27) => 
                           positive_inputs_12_27_port, shift_out(26) => 
                           positive_inputs_12_26_port, shift_out(25) => 
                           positive_inputs_12_25_port, shift_out(24) => 
                           positive_inputs_12_24_port, shift_out(23) => 
                           positive_inputs_12_23_port, shift_out(22) => 
                           positive_inputs_12_22_port, shift_out(21) => 
                           positive_inputs_12_21_port, shift_out(20) => 
                           positive_inputs_12_20_port, shift_out(19) => 
                           positive_inputs_12_19_port, shift_out(18) => 
                           positive_inputs_12_18_port, shift_out(17) => 
                           positive_inputs_12_17_port, shift_out(16) => 
                           positive_inputs_12_16_port, shift_out(15) => 
                           positive_inputs_12_15_port, shift_out(14) => 
                           positive_inputs_12_14_port, shift_out(13) => 
                           positive_inputs_12_13_port, shift_out(12) => 
                           positive_inputs_12_12_port, shift_out(11) => 
                           positive_inputs_12_11_port, shift_out(10) => 
                           positive_inputs_12_10_port, shift_out(9) => 
                           positive_inputs_12_9_port, shift_out(8) => 
                           positive_inputs_12_8_port, shift_out(7) => 
                           positive_inputs_12_7_port, shift_out(6) => 
                           positive_inputs_12_6_port, shift_out(5) => 
                           positive_inputs_12_5_port, shift_out(4) => 
                           positive_inputs_12_4_port, shift_out(3) => 
                           positive_inputs_12_3_port, shift_out(2) => 
                           positive_inputs_12_2_port, shift_out(1) => 
                           positive_inputs_12_1_port, shift_out(0) => n_1012);
   shifted_pos_13 : leftshifter_NbitShifter64_51 port map( shift_in(63) => 
                           positive_inputs_12_63_port, shift_in(62) => 
                           positive_inputs_12_62_port, shift_in(61) => 
                           positive_inputs_12_61_port, shift_in(60) => 
                           positive_inputs_12_60_port, shift_in(59) => 
                           positive_inputs_12_59_port, shift_in(58) => 
                           positive_inputs_12_58_port, shift_in(57) => 
                           positive_inputs_12_57_port, shift_in(56) => 
                           positive_inputs_12_56_port, shift_in(55) => 
                           positive_inputs_12_55_port, shift_in(54) => 
                           positive_inputs_12_54_port, shift_in(53) => 
                           positive_inputs_12_53_port, shift_in(52) => 
                           positive_inputs_12_52_port, shift_in(51) => 
                           positive_inputs_12_51_port, shift_in(50) => 
                           positive_inputs_12_50_port, shift_in(49) => 
                           positive_inputs_12_49_port, shift_in(48) => n61, 
                           shift_in(47) => positive_inputs_12_47_port, 
                           shift_in(46) => positive_inputs_12_46_port, 
                           shift_in(45) => positive_inputs_12_45_port, 
                           shift_in(44) => positive_inputs_12_44_port, 
                           shift_in(43) => positive_inputs_12_43_port, 
                           shift_in(42) => positive_inputs_12_42_port, 
                           shift_in(41) => positive_inputs_12_41_port, 
                           shift_in(40) => positive_inputs_12_40_port, 
                           shift_in(39) => positive_inputs_12_39_port, 
                           shift_in(38) => positive_inputs_12_38_port, 
                           shift_in(37) => positive_inputs_12_37_port, 
                           shift_in(36) => positive_inputs_12_36_port, 
                           shift_in(35) => positive_inputs_12_35_port, 
                           shift_in(34) => positive_inputs_12_34_port, 
                           shift_in(33) => positive_inputs_12_33_port, 
                           shift_in(32) => positive_inputs_12_32_port, 
                           shift_in(31) => positive_inputs_12_31_port, 
                           shift_in(30) => positive_inputs_12_30_port, 
                           shift_in(29) => positive_inputs_12_29_port, 
                           shift_in(28) => positive_inputs_12_28_port, 
                           shift_in(27) => positive_inputs_12_27_port, 
                           shift_in(26) => positive_inputs_12_26_port, 
                           shift_in(25) => positive_inputs_12_25_port, 
                           shift_in(24) => positive_inputs_12_24_port, 
                           shift_in(23) => positive_inputs_12_23_port, 
                           shift_in(22) => positive_inputs_12_22_port, 
                           shift_in(21) => positive_inputs_12_21_port, 
                           shift_in(20) => positive_inputs_12_20_port, 
                           shift_in(19) => positive_inputs_12_19_port, 
                           shift_in(18) => positive_inputs_12_18_port, 
                           shift_in(17) => positive_inputs_12_17_port, 
                           shift_in(16) => positive_inputs_12_16_port, 
                           shift_in(15) => positive_inputs_12_15_port, 
                           shift_in(14) => positive_inputs_12_14_port, 
                           shift_in(13) => positive_inputs_12_13_port, 
                           shift_in(12) => positive_inputs_12_12_port, 
                           shift_in(11) => positive_inputs_12_11_port, 
                           shift_in(10) => positive_inputs_12_10_port, 
                           shift_in(9) => positive_inputs_12_9_port, 
                           shift_in(8) => positive_inputs_12_8_port, 
                           shift_in(7) => positive_inputs_12_7_port, 
                           shift_in(6) => positive_inputs_12_6_port, 
                           shift_in(5) => positive_inputs_12_5_port, 
                           shift_in(4) => positive_inputs_12_4_port, 
                           shift_in(3) => positive_inputs_12_3_port, 
                           shift_in(2) => positive_inputs_12_2_port, 
                           shift_in(1) => positive_inputs_12_1_port, 
                           shift_in(0) => n9, shift_out(63) => 
                           positive_inputs_13_63_port, shift_out(62) => 
                           positive_inputs_13_62_port, shift_out(61) => 
                           positive_inputs_13_61_port, shift_out(60) => 
                           positive_inputs_13_60_port, shift_out(59) => 
                           positive_inputs_13_59_port, shift_out(58) => 
                           positive_inputs_13_58_port, shift_out(57) => 
                           positive_inputs_13_57_port, shift_out(56) => 
                           positive_inputs_13_56_port, shift_out(55) => 
                           positive_inputs_13_55_port, shift_out(54) => 
                           positive_inputs_13_54_port, shift_out(53) => 
                           positive_inputs_13_53_port, shift_out(52) => 
                           positive_inputs_13_52_port, shift_out(51) => 
                           positive_inputs_13_51_port, shift_out(50) => 
                           positive_inputs_13_50_port, shift_out(49) => 
                           positive_inputs_13_49_port, shift_out(48) => 
                           positive_inputs_13_48_port, shift_out(47) => 
                           positive_inputs_13_47_port, shift_out(46) => 
                           positive_inputs_13_46_port, shift_out(45) => 
                           positive_inputs_13_45_port, shift_out(44) => 
                           positive_inputs_13_44_port, shift_out(43) => 
                           positive_inputs_13_43_port, shift_out(42) => 
                           positive_inputs_13_42_port, shift_out(41) => 
                           positive_inputs_13_41_port, shift_out(40) => 
                           positive_inputs_13_40_port, shift_out(39) => 
                           positive_inputs_13_39_port, shift_out(38) => 
                           positive_inputs_13_38_port, shift_out(37) => 
                           positive_inputs_13_37_port, shift_out(36) => 
                           positive_inputs_13_36_port, shift_out(35) => 
                           positive_inputs_13_35_port, shift_out(34) => 
                           positive_inputs_13_34_port, shift_out(33) => 
                           positive_inputs_13_33_port, shift_out(32) => 
                           positive_inputs_13_32_port, shift_out(31) => 
                           positive_inputs_13_31_port, shift_out(30) => 
                           positive_inputs_13_30_port, shift_out(29) => 
                           positive_inputs_13_29_port, shift_out(28) => 
                           positive_inputs_13_28_port, shift_out(27) => 
                           positive_inputs_13_27_port, shift_out(26) => 
                           positive_inputs_13_26_port, shift_out(25) => 
                           positive_inputs_13_25_port, shift_out(24) => 
                           positive_inputs_13_24_port, shift_out(23) => 
                           positive_inputs_13_23_port, shift_out(22) => 
                           positive_inputs_13_22_port, shift_out(21) => 
                           positive_inputs_13_21_port, shift_out(20) => 
                           positive_inputs_13_20_port, shift_out(19) => 
                           positive_inputs_13_19_port, shift_out(18) => 
                           positive_inputs_13_18_port, shift_out(17) => 
                           positive_inputs_13_17_port, shift_out(16) => 
                           positive_inputs_13_16_port, shift_out(15) => 
                           positive_inputs_13_15_port, shift_out(14) => 
                           positive_inputs_13_14_port, shift_out(13) => 
                           positive_inputs_13_13_port, shift_out(12) => 
                           positive_inputs_13_12_port, shift_out(11) => 
                           positive_inputs_13_11_port, shift_out(10) => 
                           positive_inputs_13_10_port, shift_out(9) => 
                           positive_inputs_13_9_port, shift_out(8) => 
                           positive_inputs_13_8_port, shift_out(7) => 
                           positive_inputs_13_7_port, shift_out(6) => 
                           positive_inputs_13_6_port, shift_out(5) => 
                           positive_inputs_13_5_port, shift_out(4) => 
                           positive_inputs_13_4_port, shift_out(3) => 
                           positive_inputs_13_3_port, shift_out(2) => 
                           positive_inputs_13_2_port, shift_out(1) => 
                           positive_inputs_13_1_port, shift_out(0) => n_1013);
   shifted_pos_14 : leftshifter_NbitShifter64_50 port map( shift_in(63) => 
                           positive_inputs_13_63_port, shift_in(62) => 
                           positive_inputs_13_62_port, shift_in(61) => 
                           positive_inputs_13_61_port, shift_in(60) => 
                           positive_inputs_13_60_port, shift_in(59) => 
                           positive_inputs_13_59_port, shift_in(58) => 
                           positive_inputs_13_58_port, shift_in(57) => 
                           positive_inputs_13_57_port, shift_in(56) => 
                           positive_inputs_13_56_port, shift_in(55) => 
                           positive_inputs_13_55_port, shift_in(54) => 
                           positive_inputs_13_54_port, shift_in(53) => 
                           positive_inputs_13_53_port, shift_in(52) => 
                           positive_inputs_13_52_port, shift_in(51) => 
                           positive_inputs_13_51_port, shift_in(50) => 
                           positive_inputs_13_50_port, shift_in(49) => 
                           positive_inputs_13_49_port, shift_in(48) => n60, 
                           shift_in(47) => positive_inputs_13_47_port, 
                           shift_in(46) => positive_inputs_13_46_port, 
                           shift_in(45) => positive_inputs_13_45_port, 
                           shift_in(44) => positive_inputs_13_44_port, 
                           shift_in(43) => positive_inputs_13_43_port, 
                           shift_in(42) => positive_inputs_13_42_port, 
                           shift_in(41) => positive_inputs_13_41_port, 
                           shift_in(40) => positive_inputs_13_40_port, 
                           shift_in(39) => positive_inputs_13_39_port, 
                           shift_in(38) => positive_inputs_13_38_port, 
                           shift_in(37) => positive_inputs_13_37_port, 
                           shift_in(36) => positive_inputs_13_36_port, 
                           shift_in(35) => positive_inputs_13_35_port, 
                           shift_in(34) => positive_inputs_13_34_port, 
                           shift_in(33) => positive_inputs_13_33_port, 
                           shift_in(32) => positive_inputs_13_32_port, 
                           shift_in(31) => positive_inputs_13_31_port, 
                           shift_in(30) => positive_inputs_13_30_port, 
                           shift_in(29) => positive_inputs_13_29_port, 
                           shift_in(28) => positive_inputs_13_28_port, 
                           shift_in(27) => positive_inputs_13_27_port, 
                           shift_in(26) => positive_inputs_13_26_port, 
                           shift_in(25) => positive_inputs_13_25_port, 
                           shift_in(24) => positive_inputs_13_24_port, 
                           shift_in(23) => positive_inputs_13_23_port, 
                           shift_in(22) => positive_inputs_13_22_port, 
                           shift_in(21) => positive_inputs_13_21_port, 
                           shift_in(20) => positive_inputs_13_20_port, 
                           shift_in(19) => positive_inputs_13_19_port, 
                           shift_in(18) => positive_inputs_13_18_port, 
                           shift_in(17) => positive_inputs_13_17_port, 
                           shift_in(16) => positive_inputs_13_16_port, 
                           shift_in(15) => positive_inputs_13_15_port, 
                           shift_in(14) => positive_inputs_13_14_port, 
                           shift_in(13) => positive_inputs_13_13_port, 
                           shift_in(12) => positive_inputs_13_12_port, 
                           shift_in(11) => positive_inputs_13_11_port, 
                           shift_in(10) => positive_inputs_13_10_port, 
                           shift_in(9) => positive_inputs_13_9_port, 
                           shift_in(8) => positive_inputs_13_8_port, 
                           shift_in(7) => positive_inputs_13_7_port, 
                           shift_in(6) => positive_inputs_13_6_port, 
                           shift_in(5) => positive_inputs_13_5_port, 
                           shift_in(4) => positive_inputs_13_4_port, 
                           shift_in(3) => positive_inputs_13_3_port, 
                           shift_in(2) => positive_inputs_13_2_port, 
                           shift_in(1) => positive_inputs_13_1_port, 
                           shift_in(0) => n9, shift_out(63) => 
                           positive_inputs_14_63_port, shift_out(62) => 
                           positive_inputs_14_62_port, shift_out(61) => 
                           positive_inputs_14_61_port, shift_out(60) => 
                           positive_inputs_14_60_port, shift_out(59) => 
                           positive_inputs_14_59_port, shift_out(58) => 
                           positive_inputs_14_58_port, shift_out(57) => 
                           positive_inputs_14_57_port, shift_out(56) => 
                           positive_inputs_14_56_port, shift_out(55) => 
                           positive_inputs_14_55_port, shift_out(54) => 
                           positive_inputs_14_54_port, shift_out(53) => 
                           positive_inputs_14_53_port, shift_out(52) => 
                           positive_inputs_14_52_port, shift_out(51) => 
                           positive_inputs_14_51_port, shift_out(50) => 
                           positive_inputs_14_50_port, shift_out(49) => 
                           positive_inputs_14_49_port, shift_out(48) => 
                           positive_inputs_14_48_port, shift_out(47) => 
                           positive_inputs_14_47_port, shift_out(46) => 
                           positive_inputs_14_46_port, shift_out(45) => 
                           positive_inputs_14_45_port, shift_out(44) => 
                           positive_inputs_14_44_port, shift_out(43) => 
                           positive_inputs_14_43_port, shift_out(42) => 
                           positive_inputs_14_42_port, shift_out(41) => 
                           positive_inputs_14_41_port, shift_out(40) => 
                           positive_inputs_14_40_port, shift_out(39) => 
                           positive_inputs_14_39_port, shift_out(38) => 
                           positive_inputs_14_38_port, shift_out(37) => 
                           positive_inputs_14_37_port, shift_out(36) => 
                           positive_inputs_14_36_port, shift_out(35) => 
                           positive_inputs_14_35_port, shift_out(34) => 
                           positive_inputs_14_34_port, shift_out(33) => 
                           positive_inputs_14_33_port, shift_out(32) => 
                           positive_inputs_14_32_port, shift_out(31) => 
                           positive_inputs_14_31_port, shift_out(30) => 
                           positive_inputs_14_30_port, shift_out(29) => 
                           positive_inputs_14_29_port, shift_out(28) => 
                           positive_inputs_14_28_port, shift_out(27) => 
                           positive_inputs_14_27_port, shift_out(26) => 
                           positive_inputs_14_26_port, shift_out(25) => 
                           positive_inputs_14_25_port, shift_out(24) => 
                           positive_inputs_14_24_port, shift_out(23) => 
                           positive_inputs_14_23_port, shift_out(22) => 
                           positive_inputs_14_22_port, shift_out(21) => 
                           positive_inputs_14_21_port, shift_out(20) => 
                           positive_inputs_14_20_port, shift_out(19) => 
                           positive_inputs_14_19_port, shift_out(18) => 
                           positive_inputs_14_18_port, shift_out(17) => 
                           positive_inputs_14_17_port, shift_out(16) => 
                           positive_inputs_14_16_port, shift_out(15) => 
                           positive_inputs_14_15_port, shift_out(14) => 
                           positive_inputs_14_14_port, shift_out(13) => 
                           positive_inputs_14_13_port, shift_out(12) => 
                           positive_inputs_14_12_port, shift_out(11) => 
                           positive_inputs_14_11_port, shift_out(10) => 
                           positive_inputs_14_10_port, shift_out(9) => 
                           positive_inputs_14_9_port, shift_out(8) => 
                           positive_inputs_14_8_port, shift_out(7) => 
                           positive_inputs_14_7_port, shift_out(6) => 
                           positive_inputs_14_6_port, shift_out(5) => 
                           positive_inputs_14_5_port, shift_out(4) => 
                           positive_inputs_14_4_port, shift_out(3) => 
                           positive_inputs_14_3_port, shift_out(2) => 
                           positive_inputs_14_2_port, shift_out(1) => 
                           positive_inputs_14_1_port, shift_out(0) => n_1014);
   shifted_pos_15 : leftshifter_NbitShifter64_49 port map( shift_in(63) => 
                           positive_inputs_14_63_port, shift_in(62) => 
                           positive_inputs_14_62_port, shift_in(61) => 
                           positive_inputs_14_61_port, shift_in(60) => 
                           positive_inputs_14_60_port, shift_in(59) => 
                           positive_inputs_14_59_port, shift_in(58) => 
                           positive_inputs_14_58_port, shift_in(57) => 
                           positive_inputs_14_57_port, shift_in(56) => 
                           positive_inputs_14_56_port, shift_in(55) => 
                           positive_inputs_14_55_port, shift_in(54) => 
                           positive_inputs_14_54_port, shift_in(53) => 
                           positive_inputs_14_53_port, shift_in(52) => 
                           positive_inputs_14_52_port, shift_in(51) => 
                           positive_inputs_14_51_port, shift_in(50) => 
                           positive_inputs_14_50_port, shift_in(49) => 
                           positive_inputs_14_49_port, shift_in(48) => n59, 
                           shift_in(47) => positive_inputs_14_47_port, 
                           shift_in(46) => positive_inputs_14_46_port, 
                           shift_in(45) => positive_inputs_14_45_port, 
                           shift_in(44) => positive_inputs_14_44_port, 
                           shift_in(43) => positive_inputs_14_43_port, 
                           shift_in(42) => positive_inputs_14_42_port, 
                           shift_in(41) => positive_inputs_14_41_port, 
                           shift_in(40) => positive_inputs_14_40_port, 
                           shift_in(39) => positive_inputs_14_39_port, 
                           shift_in(38) => positive_inputs_14_38_port, 
                           shift_in(37) => positive_inputs_14_37_port, 
                           shift_in(36) => positive_inputs_14_36_port, 
                           shift_in(35) => positive_inputs_14_35_port, 
                           shift_in(34) => positive_inputs_14_34_port, 
                           shift_in(33) => positive_inputs_14_33_port, 
                           shift_in(32) => positive_inputs_14_32_port, 
                           shift_in(31) => positive_inputs_14_31_port, 
                           shift_in(30) => positive_inputs_14_30_port, 
                           shift_in(29) => positive_inputs_14_29_port, 
                           shift_in(28) => positive_inputs_14_28_port, 
                           shift_in(27) => positive_inputs_14_27_port, 
                           shift_in(26) => positive_inputs_14_26_port, 
                           shift_in(25) => positive_inputs_14_25_port, 
                           shift_in(24) => positive_inputs_14_24_port, 
                           shift_in(23) => positive_inputs_14_23_port, 
                           shift_in(22) => positive_inputs_14_22_port, 
                           shift_in(21) => positive_inputs_14_21_port, 
                           shift_in(20) => positive_inputs_14_20_port, 
                           shift_in(19) => positive_inputs_14_19_port, 
                           shift_in(18) => positive_inputs_14_18_port, 
                           shift_in(17) => positive_inputs_14_17_port, 
                           shift_in(16) => positive_inputs_14_16_port, 
                           shift_in(15) => positive_inputs_14_15_port, 
                           shift_in(14) => positive_inputs_14_14_port, 
                           shift_in(13) => positive_inputs_14_13_port, 
                           shift_in(12) => positive_inputs_14_12_port, 
                           shift_in(11) => positive_inputs_14_11_port, 
                           shift_in(10) => positive_inputs_14_10_port, 
                           shift_in(9) => positive_inputs_14_9_port, 
                           shift_in(8) => positive_inputs_14_8_port, 
                           shift_in(7) => positive_inputs_14_7_port, 
                           shift_in(6) => positive_inputs_14_6_port, 
                           shift_in(5) => positive_inputs_14_5_port, 
                           shift_in(4) => positive_inputs_14_4_port, 
                           shift_in(3) => positive_inputs_14_3_port, 
                           shift_in(2) => positive_inputs_14_2_port, 
                           shift_in(1) => positive_inputs_14_1_port, 
                           shift_in(0) => n9, shift_out(63) => 
                           positive_inputs_15_63_port, shift_out(62) => 
                           positive_inputs_15_62_port, shift_out(61) => 
                           positive_inputs_15_61_port, shift_out(60) => 
                           positive_inputs_15_60_port, shift_out(59) => 
                           positive_inputs_15_59_port, shift_out(58) => 
                           positive_inputs_15_58_port, shift_out(57) => 
                           positive_inputs_15_57_port, shift_out(56) => 
                           positive_inputs_15_56_port, shift_out(55) => 
                           positive_inputs_15_55_port, shift_out(54) => 
                           positive_inputs_15_54_port, shift_out(53) => 
                           positive_inputs_15_53_port, shift_out(52) => 
                           positive_inputs_15_52_port, shift_out(51) => 
                           positive_inputs_15_51_port, shift_out(50) => 
                           positive_inputs_15_50_port, shift_out(49) => 
                           positive_inputs_15_49_port, shift_out(48) => 
                           positive_inputs_15_48_port, shift_out(47) => 
                           positive_inputs_15_47_port, shift_out(46) => 
                           positive_inputs_15_46_port, shift_out(45) => 
                           positive_inputs_15_45_port, shift_out(44) => 
                           positive_inputs_15_44_port, shift_out(43) => 
                           positive_inputs_15_43_port, shift_out(42) => 
                           positive_inputs_15_42_port, shift_out(41) => 
                           positive_inputs_15_41_port, shift_out(40) => 
                           positive_inputs_15_40_port, shift_out(39) => 
                           positive_inputs_15_39_port, shift_out(38) => 
                           positive_inputs_15_38_port, shift_out(37) => 
                           positive_inputs_15_37_port, shift_out(36) => 
                           positive_inputs_15_36_port, shift_out(35) => 
                           positive_inputs_15_35_port, shift_out(34) => 
                           positive_inputs_15_34_port, shift_out(33) => 
                           positive_inputs_15_33_port, shift_out(32) => 
                           positive_inputs_15_32_port, shift_out(31) => 
                           positive_inputs_15_31_port, shift_out(30) => 
                           positive_inputs_15_30_port, shift_out(29) => 
                           positive_inputs_15_29_port, shift_out(28) => 
                           positive_inputs_15_28_port, shift_out(27) => 
                           positive_inputs_15_27_port, shift_out(26) => 
                           positive_inputs_15_26_port, shift_out(25) => 
                           positive_inputs_15_25_port, shift_out(24) => 
                           positive_inputs_15_24_port, shift_out(23) => 
                           positive_inputs_15_23_port, shift_out(22) => 
                           positive_inputs_15_22_port, shift_out(21) => 
                           positive_inputs_15_21_port, shift_out(20) => 
                           positive_inputs_15_20_port, shift_out(19) => 
                           positive_inputs_15_19_port, shift_out(18) => 
                           positive_inputs_15_18_port, shift_out(17) => 
                           positive_inputs_15_17_port, shift_out(16) => 
                           positive_inputs_15_16_port, shift_out(15) => 
                           positive_inputs_15_15_port, shift_out(14) => 
                           positive_inputs_15_14_port, shift_out(13) => 
                           positive_inputs_15_13_port, shift_out(12) => 
                           positive_inputs_15_12_port, shift_out(11) => 
                           positive_inputs_15_11_port, shift_out(10) => 
                           positive_inputs_15_10_port, shift_out(9) => 
                           positive_inputs_15_9_port, shift_out(8) => 
                           positive_inputs_15_8_port, shift_out(7) => 
                           positive_inputs_15_7_port, shift_out(6) => 
                           positive_inputs_15_6_port, shift_out(5) => 
                           positive_inputs_15_5_port, shift_out(4) => 
                           positive_inputs_15_4_port, shift_out(3) => 
                           positive_inputs_15_3_port, shift_out(2) => 
                           positive_inputs_15_2_port, shift_out(1) => 
                           positive_inputs_15_1_port, shift_out(0) => n_1015);
   shifted_pos_16 : leftshifter_NbitShifter64_48 port map( shift_in(63) => 
                           positive_inputs_15_63_port, shift_in(62) => 
                           positive_inputs_15_62_port, shift_in(61) => 
                           positive_inputs_15_61_port, shift_in(60) => 
                           positive_inputs_15_60_port, shift_in(59) => 
                           positive_inputs_15_59_port, shift_in(58) => 
                           positive_inputs_15_58_port, shift_in(57) => 
                           positive_inputs_15_57_port, shift_in(56) => 
                           positive_inputs_15_56_port, shift_in(55) => 
                           positive_inputs_15_55_port, shift_in(54) => 
                           positive_inputs_15_54_port, shift_in(53) => 
                           positive_inputs_15_53_port, shift_in(52) => 
                           positive_inputs_15_52_port, shift_in(51) => 
                           positive_inputs_15_51_port, shift_in(50) => 
                           positive_inputs_15_50_port, shift_in(49) => 
                           positive_inputs_15_49_port, shift_in(48) => n58, 
                           shift_in(47) => positive_inputs_15_47_port, 
                           shift_in(46) => positive_inputs_15_46_port, 
                           shift_in(45) => positive_inputs_15_45_port, 
                           shift_in(44) => positive_inputs_15_44_port, 
                           shift_in(43) => positive_inputs_15_43_port, 
                           shift_in(42) => positive_inputs_15_42_port, 
                           shift_in(41) => positive_inputs_15_41_port, 
                           shift_in(40) => positive_inputs_15_40_port, 
                           shift_in(39) => positive_inputs_15_39_port, 
                           shift_in(38) => positive_inputs_15_38_port, 
                           shift_in(37) => positive_inputs_15_37_port, 
                           shift_in(36) => positive_inputs_15_36_port, 
                           shift_in(35) => positive_inputs_15_35_port, 
                           shift_in(34) => positive_inputs_15_34_port, 
                           shift_in(33) => positive_inputs_15_33_port, 
                           shift_in(32) => positive_inputs_15_32_port, 
                           shift_in(31) => positive_inputs_15_31_port, 
                           shift_in(30) => positive_inputs_15_30_port, 
                           shift_in(29) => positive_inputs_15_29_port, 
                           shift_in(28) => positive_inputs_15_28_port, 
                           shift_in(27) => positive_inputs_15_27_port, 
                           shift_in(26) => positive_inputs_15_26_port, 
                           shift_in(25) => positive_inputs_15_25_port, 
                           shift_in(24) => positive_inputs_15_24_port, 
                           shift_in(23) => positive_inputs_15_23_port, 
                           shift_in(22) => positive_inputs_15_22_port, 
                           shift_in(21) => positive_inputs_15_21_port, 
                           shift_in(20) => positive_inputs_15_20_port, 
                           shift_in(19) => positive_inputs_15_19_port, 
                           shift_in(18) => positive_inputs_15_18_port, 
                           shift_in(17) => positive_inputs_15_17_port, 
                           shift_in(16) => positive_inputs_15_16_port, 
                           shift_in(15) => positive_inputs_15_15_port, 
                           shift_in(14) => positive_inputs_15_14_port, 
                           shift_in(13) => positive_inputs_15_13_port, 
                           shift_in(12) => positive_inputs_15_12_port, 
                           shift_in(11) => positive_inputs_15_11_port, 
                           shift_in(10) => positive_inputs_15_10_port, 
                           shift_in(9) => positive_inputs_15_9_port, 
                           shift_in(8) => positive_inputs_15_8_port, 
                           shift_in(7) => positive_inputs_15_7_port, 
                           shift_in(6) => positive_inputs_15_6_port, 
                           shift_in(5) => positive_inputs_15_5_port, 
                           shift_in(4) => positive_inputs_15_4_port, 
                           shift_in(3) => positive_inputs_15_3_port, 
                           shift_in(2) => positive_inputs_15_2_port, 
                           shift_in(1) => positive_inputs_15_1_port, 
                           shift_in(0) => n9, shift_out(63) => 
                           positive_inputs_16_63_port, shift_out(62) => 
                           positive_inputs_16_62_port, shift_out(61) => 
                           positive_inputs_16_61_port, shift_out(60) => 
                           positive_inputs_16_60_port, shift_out(59) => 
                           positive_inputs_16_59_port, shift_out(58) => 
                           positive_inputs_16_58_port, shift_out(57) => 
                           positive_inputs_16_57_port, shift_out(56) => 
                           positive_inputs_16_56_port, shift_out(55) => 
                           positive_inputs_16_55_port, shift_out(54) => 
                           positive_inputs_16_54_port, shift_out(53) => 
                           positive_inputs_16_53_port, shift_out(52) => 
                           positive_inputs_16_52_port, shift_out(51) => 
                           positive_inputs_16_51_port, shift_out(50) => 
                           positive_inputs_16_50_port, shift_out(49) => 
                           positive_inputs_16_49_port, shift_out(48) => 
                           positive_inputs_16_48_port, shift_out(47) => 
                           positive_inputs_16_47_port, shift_out(46) => 
                           positive_inputs_16_46_port, shift_out(45) => 
                           positive_inputs_16_45_port, shift_out(44) => 
                           positive_inputs_16_44_port, shift_out(43) => 
                           positive_inputs_16_43_port, shift_out(42) => 
                           positive_inputs_16_42_port, shift_out(41) => 
                           positive_inputs_16_41_port, shift_out(40) => 
                           positive_inputs_16_40_port, shift_out(39) => 
                           positive_inputs_16_39_port, shift_out(38) => 
                           positive_inputs_16_38_port, shift_out(37) => 
                           positive_inputs_16_37_port, shift_out(36) => 
                           positive_inputs_16_36_port, shift_out(35) => 
                           positive_inputs_16_35_port, shift_out(34) => 
                           positive_inputs_16_34_port, shift_out(33) => 
                           positive_inputs_16_33_port, shift_out(32) => 
                           positive_inputs_16_32_port, shift_out(31) => 
                           positive_inputs_16_31_port, shift_out(30) => 
                           positive_inputs_16_30_port, shift_out(29) => 
                           positive_inputs_16_29_port, shift_out(28) => 
                           positive_inputs_16_28_port, shift_out(27) => 
                           positive_inputs_16_27_port, shift_out(26) => 
                           positive_inputs_16_26_port, shift_out(25) => 
                           positive_inputs_16_25_port, shift_out(24) => 
                           positive_inputs_16_24_port, shift_out(23) => 
                           positive_inputs_16_23_port, shift_out(22) => 
                           positive_inputs_16_22_port, shift_out(21) => 
                           positive_inputs_16_21_port, shift_out(20) => 
                           positive_inputs_16_20_port, shift_out(19) => 
                           positive_inputs_16_19_port, shift_out(18) => 
                           positive_inputs_16_18_port, shift_out(17) => 
                           positive_inputs_16_17_port, shift_out(16) => 
                           positive_inputs_16_16_port, shift_out(15) => 
                           positive_inputs_16_15_port, shift_out(14) => 
                           positive_inputs_16_14_port, shift_out(13) => 
                           positive_inputs_16_13_port, shift_out(12) => 
                           positive_inputs_16_12_port, shift_out(11) => 
                           positive_inputs_16_11_port, shift_out(10) => 
                           positive_inputs_16_10_port, shift_out(9) => 
                           positive_inputs_16_9_port, shift_out(8) => 
                           positive_inputs_16_8_port, shift_out(7) => 
                           positive_inputs_16_7_port, shift_out(6) => 
                           positive_inputs_16_6_port, shift_out(5) => 
                           positive_inputs_16_5_port, shift_out(4) => 
                           positive_inputs_16_4_port, shift_out(3) => 
                           positive_inputs_16_3_port, shift_out(2) => 
                           positive_inputs_16_2_port, shift_out(1) => 
                           positive_inputs_16_1_port, shift_out(0) => n_1016);
   shifted_pos_17 : leftshifter_NbitShifter64_47 port map( shift_in(63) => 
                           positive_inputs_16_63_port, shift_in(62) => 
                           positive_inputs_16_62_port, shift_in(61) => 
                           positive_inputs_16_61_port, shift_in(60) => 
                           positive_inputs_16_60_port, shift_in(59) => 
                           positive_inputs_16_59_port, shift_in(58) => 
                           positive_inputs_16_58_port, shift_in(57) => 
                           positive_inputs_16_57_port, shift_in(56) => 
                           positive_inputs_16_56_port, shift_in(55) => 
                           positive_inputs_16_55_port, shift_in(54) => 
                           positive_inputs_16_54_port, shift_in(53) => 
                           positive_inputs_16_53_port, shift_in(52) => 
                           positive_inputs_16_52_port, shift_in(51) => 
                           positive_inputs_16_51_port, shift_in(50) => 
                           positive_inputs_16_50_port, shift_in(49) => 
                           positive_inputs_16_49_port, shift_in(48) => n57, 
                           shift_in(47) => n56, shift_in(46) => n215, 
                           shift_in(45) => n213, shift_in(44) => n211, 
                           shift_in(43) => n209, shift_in(42) => n207, 
                           shift_in(41) => n205, shift_in(40) => n203, 
                           shift_in(39) => n201, shift_in(38) => n199, 
                           shift_in(37) => n197, shift_in(36) => n195, 
                           shift_in(35) => n193, shift_in(34) => n191, 
                           shift_in(33) => n189, shift_in(32) => n187, 
                           shift_in(31) => n185, shift_in(30) => n183, 
                           shift_in(29) => n181, shift_in(28) => n179, 
                           shift_in(27) => n177, shift_in(26) => n175, 
                           shift_in(25) => n173, shift_in(24) => n171, 
                           shift_in(23) => n169, shift_in(22) => n167, 
                           shift_in(21) => n165, shift_in(20) => n163, 
                           shift_in(19) => n161, shift_in(18) => n159, 
                           shift_in(17) => n157, shift_in(16) => n155, 
                           shift_in(15) => positive_inputs_16_15_port, 
                           shift_in(14) => positive_inputs_16_14_port, 
                           shift_in(13) => positive_inputs_16_13_port, 
                           shift_in(12) => positive_inputs_16_12_port, 
                           shift_in(11) => positive_inputs_16_11_port, 
                           shift_in(10) => positive_inputs_16_10_port, 
                           shift_in(9) => positive_inputs_16_9_port, 
                           shift_in(8) => positive_inputs_16_8_port, 
                           shift_in(7) => positive_inputs_16_7_port, 
                           shift_in(6) => positive_inputs_16_6_port, 
                           shift_in(5) => positive_inputs_16_5_port, 
                           shift_in(4) => positive_inputs_16_4_port, 
                           shift_in(3) => positive_inputs_16_3_port, 
                           shift_in(2) => positive_inputs_16_2_port, 
                           shift_in(1) => positive_inputs_16_1_port, 
                           shift_in(0) => n9, shift_out(63) => 
                           positive_inputs_17_63_port, shift_out(62) => 
                           positive_inputs_17_62_port, shift_out(61) => 
                           positive_inputs_17_61_port, shift_out(60) => 
                           positive_inputs_17_60_port, shift_out(59) => 
                           positive_inputs_17_59_port, shift_out(58) => 
                           positive_inputs_17_58_port, shift_out(57) => 
                           positive_inputs_17_57_port, shift_out(56) => 
                           positive_inputs_17_56_port, shift_out(55) => 
                           positive_inputs_17_55_port, shift_out(54) => 
                           positive_inputs_17_54_port, shift_out(53) => 
                           positive_inputs_17_53_port, shift_out(52) => 
                           positive_inputs_17_52_port, shift_out(51) => 
                           positive_inputs_17_51_port, shift_out(50) => 
                           positive_inputs_17_50_port, shift_out(49) => 
                           positive_inputs_17_49_port, shift_out(48) => 
                           positive_inputs_17_48_port, shift_out(47) => 
                           positive_inputs_17_47_port, shift_out(46) => 
                           positive_inputs_17_46_port, shift_out(45) => 
                           positive_inputs_17_45_port, shift_out(44) => 
                           positive_inputs_17_44_port, shift_out(43) => 
                           positive_inputs_17_43_port, shift_out(42) => 
                           positive_inputs_17_42_port, shift_out(41) => 
                           positive_inputs_17_41_port, shift_out(40) => 
                           positive_inputs_17_40_port, shift_out(39) => 
                           positive_inputs_17_39_port, shift_out(38) => 
                           positive_inputs_17_38_port, shift_out(37) => 
                           positive_inputs_17_37_port, shift_out(36) => 
                           positive_inputs_17_36_port, shift_out(35) => 
                           positive_inputs_17_35_port, shift_out(34) => 
                           positive_inputs_17_34_port, shift_out(33) => 
                           positive_inputs_17_33_port, shift_out(32) => 
                           positive_inputs_17_32_port, shift_out(31) => 
                           positive_inputs_17_31_port, shift_out(30) => 
                           positive_inputs_17_30_port, shift_out(29) => 
                           positive_inputs_17_29_port, shift_out(28) => 
                           positive_inputs_17_28_port, shift_out(27) => 
                           positive_inputs_17_27_port, shift_out(26) => 
                           positive_inputs_17_26_port, shift_out(25) => 
                           positive_inputs_17_25_port, shift_out(24) => 
                           positive_inputs_17_24_port, shift_out(23) => 
                           positive_inputs_17_23_port, shift_out(22) => 
                           positive_inputs_17_22_port, shift_out(21) => 
                           positive_inputs_17_21_port, shift_out(20) => 
                           positive_inputs_17_20_port, shift_out(19) => 
                           positive_inputs_17_19_port, shift_out(18) => 
                           positive_inputs_17_18_port, shift_out(17) => 
                           positive_inputs_17_17_port, shift_out(16) => 
                           positive_inputs_17_16_port, shift_out(15) => 
                           positive_inputs_17_15_port, shift_out(14) => 
                           positive_inputs_17_14_port, shift_out(13) => 
                           positive_inputs_17_13_port, shift_out(12) => 
                           positive_inputs_17_12_port, shift_out(11) => 
                           positive_inputs_17_11_port, shift_out(10) => 
                           positive_inputs_17_10_port, shift_out(9) => 
                           positive_inputs_17_9_port, shift_out(8) => 
                           positive_inputs_17_8_port, shift_out(7) => 
                           positive_inputs_17_7_port, shift_out(6) => 
                           positive_inputs_17_6_port, shift_out(5) => 
                           positive_inputs_17_5_port, shift_out(4) => 
                           positive_inputs_17_4_port, shift_out(3) => 
                           positive_inputs_17_3_port, shift_out(2) => 
                           positive_inputs_17_2_port, shift_out(1) => 
                           positive_inputs_17_1_port, shift_out(0) => n_1017);
   shifted_pos_18 : leftshifter_NbitShifter64_46 port map( shift_in(63) => 
                           positive_inputs_17_63_port, shift_in(62) => 
                           positive_inputs_17_62_port, shift_in(61) => 
                           positive_inputs_17_61_port, shift_in(60) => 
                           positive_inputs_17_60_port, shift_in(59) => 
                           positive_inputs_17_59_port, shift_in(58) => 
                           positive_inputs_17_58_port, shift_in(57) => 
                           positive_inputs_17_57_port, shift_in(56) => 
                           positive_inputs_17_56_port, shift_in(55) => 
                           positive_inputs_17_55_port, shift_in(54) => 
                           positive_inputs_17_54_port, shift_in(53) => 
                           positive_inputs_17_53_port, shift_in(52) => 
                           positive_inputs_17_52_port, shift_in(51) => 
                           positive_inputs_17_51_port, shift_in(50) => 
                           positive_inputs_17_50_port, shift_in(49) => 
                           positive_inputs_17_49_port, shift_in(48) => 
                           positive_inputs_17_48_port, shift_in(47) => 
                           positive_inputs_17_47_port, shift_in(46) => 
                           positive_inputs_17_46_port, shift_in(45) => 
                           positive_inputs_17_45_port, shift_in(44) => 
                           positive_inputs_17_44_port, shift_in(43) => 
                           positive_inputs_17_43_port, shift_in(42) => 
                           positive_inputs_17_42_port, shift_in(41) => 
                           positive_inputs_17_41_port, shift_in(40) => 
                           positive_inputs_17_40_port, shift_in(39) => 
                           positive_inputs_17_39_port, shift_in(38) => 
                           positive_inputs_17_38_port, shift_in(37) => 
                           positive_inputs_17_37_port, shift_in(36) => 
                           positive_inputs_17_36_port, shift_in(35) => 
                           positive_inputs_17_35_port, shift_in(34) => 
                           positive_inputs_17_34_port, shift_in(33) => 
                           positive_inputs_17_33_port, shift_in(32) => 
                           positive_inputs_17_32_port, shift_in(31) => 
                           positive_inputs_17_31_port, shift_in(30) => 
                           positive_inputs_17_30_port, shift_in(29) => 
                           positive_inputs_17_29_port, shift_in(28) => 
                           positive_inputs_17_28_port, shift_in(27) => 
                           positive_inputs_17_27_port, shift_in(26) => 
                           positive_inputs_17_26_port, shift_in(25) => 
                           positive_inputs_17_25_port, shift_in(24) => 
                           positive_inputs_17_24_port, shift_in(23) => 
                           positive_inputs_17_23_port, shift_in(22) => 
                           positive_inputs_17_22_port, shift_in(21) => 
                           positive_inputs_17_21_port, shift_in(20) => 
                           positive_inputs_17_20_port, shift_in(19) => 
                           positive_inputs_17_19_port, shift_in(18) => 
                           positive_inputs_17_18_port, shift_in(17) => 
                           positive_inputs_17_17_port, shift_in(16) => 
                           positive_inputs_17_16_port, shift_in(15) => 
                           positive_inputs_17_15_port, shift_in(14) => 
                           positive_inputs_17_14_port, shift_in(13) => 
                           positive_inputs_17_13_port, shift_in(12) => 
                           positive_inputs_17_12_port, shift_in(11) => 
                           positive_inputs_17_11_port, shift_in(10) => 
                           positive_inputs_17_10_port, shift_in(9) => 
                           positive_inputs_17_9_port, shift_in(8) => 
                           positive_inputs_17_8_port, shift_in(7) => 
                           positive_inputs_17_7_port, shift_in(6) => 
                           positive_inputs_17_6_port, shift_in(5) => 
                           positive_inputs_17_5_port, shift_in(4) => 
                           positive_inputs_17_4_port, shift_in(3) => 
                           positive_inputs_17_3_port, shift_in(2) => 
                           positive_inputs_17_2_port, shift_in(1) => 
                           positive_inputs_17_1_port, shift_in(0) => n9, 
                           shift_out(63) => positive_inputs_18_63_port, 
                           shift_out(62) => positive_inputs_18_62_port, 
                           shift_out(61) => positive_inputs_18_61_port, 
                           shift_out(60) => positive_inputs_18_60_port, 
                           shift_out(59) => positive_inputs_18_59_port, 
                           shift_out(58) => positive_inputs_18_58_port, 
                           shift_out(57) => positive_inputs_18_57_port, 
                           shift_out(56) => positive_inputs_18_56_port, 
                           shift_out(55) => positive_inputs_18_55_port, 
                           shift_out(54) => positive_inputs_18_54_port, 
                           shift_out(53) => positive_inputs_18_53_port, 
                           shift_out(52) => positive_inputs_18_52_port, 
                           shift_out(51) => positive_inputs_18_51_port, 
                           shift_out(50) => positive_inputs_18_50_port, 
                           shift_out(49) => positive_inputs_18_49_port, 
                           shift_out(48) => positive_inputs_18_48_port, 
                           shift_out(47) => positive_inputs_18_47_port, 
                           shift_out(46) => positive_inputs_18_46_port, 
                           shift_out(45) => positive_inputs_18_45_port, 
                           shift_out(44) => positive_inputs_18_44_port, 
                           shift_out(43) => positive_inputs_18_43_port, 
                           shift_out(42) => positive_inputs_18_42_port, 
                           shift_out(41) => positive_inputs_18_41_port, 
                           shift_out(40) => positive_inputs_18_40_port, 
                           shift_out(39) => positive_inputs_18_39_port, 
                           shift_out(38) => positive_inputs_18_38_port, 
                           shift_out(37) => positive_inputs_18_37_port, 
                           shift_out(36) => positive_inputs_18_36_port, 
                           shift_out(35) => positive_inputs_18_35_port, 
                           shift_out(34) => positive_inputs_18_34_port, 
                           shift_out(33) => positive_inputs_18_33_port, 
                           shift_out(32) => positive_inputs_18_32_port, 
                           shift_out(31) => positive_inputs_18_31_port, 
                           shift_out(30) => positive_inputs_18_30_port, 
                           shift_out(29) => positive_inputs_18_29_port, 
                           shift_out(28) => positive_inputs_18_28_port, 
                           shift_out(27) => positive_inputs_18_27_port, 
                           shift_out(26) => positive_inputs_18_26_port, 
                           shift_out(25) => positive_inputs_18_25_port, 
                           shift_out(24) => positive_inputs_18_24_port, 
                           shift_out(23) => positive_inputs_18_23_port, 
                           shift_out(22) => positive_inputs_18_22_port, 
                           shift_out(21) => positive_inputs_18_21_port, 
                           shift_out(20) => positive_inputs_18_20_port, 
                           shift_out(19) => positive_inputs_18_19_port, 
                           shift_out(18) => positive_inputs_18_18_port, 
                           shift_out(17) => positive_inputs_18_17_port, 
                           shift_out(16) => positive_inputs_18_16_port, 
                           shift_out(15) => positive_inputs_18_15_port, 
                           shift_out(14) => positive_inputs_18_14_port, 
                           shift_out(13) => positive_inputs_18_13_port, 
                           shift_out(12) => positive_inputs_18_12_port, 
                           shift_out(11) => positive_inputs_18_11_port, 
                           shift_out(10) => positive_inputs_18_10_port, 
                           shift_out(9) => positive_inputs_18_9_port, 
                           shift_out(8) => positive_inputs_18_8_port, 
                           shift_out(7) => positive_inputs_18_7_port, 
                           shift_out(6) => positive_inputs_18_6_port, 
                           shift_out(5) => positive_inputs_18_5_port, 
                           shift_out(4) => positive_inputs_18_4_port, 
                           shift_out(3) => positive_inputs_18_3_port, 
                           shift_out(2) => positive_inputs_18_2_port, 
                           shift_out(1) => positive_inputs_18_1_port, 
                           shift_out(0) => n_1018);
   shifted_pos_19 : leftshifter_NbitShifter64_45 port map( shift_in(63) => 
                           positive_inputs_18_63_port, shift_in(62) => 
                           positive_inputs_18_62_port, shift_in(61) => 
                           positive_inputs_18_61_port, shift_in(60) => 
                           positive_inputs_18_60_port, shift_in(59) => 
                           positive_inputs_18_59_port, shift_in(58) => 
                           positive_inputs_18_58_port, shift_in(57) => 
                           positive_inputs_18_57_port, shift_in(56) => 
                           positive_inputs_18_56_port, shift_in(55) => 
                           positive_inputs_18_55_port, shift_in(54) => 
                           positive_inputs_18_54_port, shift_in(53) => 
                           positive_inputs_18_53_port, shift_in(52) => 
                           positive_inputs_18_52_port, shift_in(51) => 
                           positive_inputs_18_51_port, shift_in(50) => 
                           positive_inputs_18_50_port, shift_in(49) => 
                           positive_inputs_18_49_port, shift_in(48) => 
                           positive_inputs_18_48_port, shift_in(47) => 
                           positive_inputs_18_47_port, shift_in(46) => 
                           positive_inputs_18_46_port, shift_in(45) => 
                           positive_inputs_18_45_port, shift_in(44) => 
                           positive_inputs_18_44_port, shift_in(43) => 
                           positive_inputs_18_43_port, shift_in(42) => 
                           positive_inputs_18_42_port, shift_in(41) => 
                           positive_inputs_18_41_port, shift_in(40) => 
                           positive_inputs_18_40_port, shift_in(39) => 
                           positive_inputs_18_39_port, shift_in(38) => 
                           positive_inputs_18_38_port, shift_in(37) => 
                           positive_inputs_18_37_port, shift_in(36) => 
                           positive_inputs_18_36_port, shift_in(35) => 
                           positive_inputs_18_35_port, shift_in(34) => 
                           positive_inputs_18_34_port, shift_in(33) => 
                           positive_inputs_18_33_port, shift_in(32) => 
                           positive_inputs_18_32_port, shift_in(31) => 
                           positive_inputs_18_31_port, shift_in(30) => 
                           positive_inputs_18_30_port, shift_in(29) => 
                           positive_inputs_18_29_port, shift_in(28) => 
                           positive_inputs_18_28_port, shift_in(27) => 
                           positive_inputs_18_27_port, shift_in(26) => 
                           positive_inputs_18_26_port, shift_in(25) => 
                           positive_inputs_18_25_port, shift_in(24) => 
                           positive_inputs_18_24_port, shift_in(23) => 
                           positive_inputs_18_23_port, shift_in(22) => 
                           positive_inputs_18_22_port, shift_in(21) => 
                           positive_inputs_18_21_port, shift_in(20) => 
                           positive_inputs_18_20_port, shift_in(19) => 
                           positive_inputs_18_19_port, shift_in(18) => 
                           positive_inputs_18_18_port, shift_in(17) => 
                           positive_inputs_18_17_port, shift_in(16) => 
                           positive_inputs_18_16_port, shift_in(15) => 
                           positive_inputs_18_15_port, shift_in(14) => 
                           positive_inputs_18_14_port, shift_in(13) => 
                           positive_inputs_18_13_port, shift_in(12) => 
                           positive_inputs_18_12_port, shift_in(11) => 
                           positive_inputs_18_11_port, shift_in(10) => 
                           positive_inputs_18_10_port, shift_in(9) => 
                           positive_inputs_18_9_port, shift_in(8) => 
                           positive_inputs_18_8_port, shift_in(7) => 
                           positive_inputs_18_7_port, shift_in(6) => 
                           positive_inputs_18_6_port, shift_in(5) => 
                           positive_inputs_18_5_port, shift_in(4) => 
                           positive_inputs_18_4_port, shift_in(3) => 
                           positive_inputs_18_3_port, shift_in(2) => 
                           positive_inputs_18_2_port, shift_in(1) => 
                           positive_inputs_18_1_port, shift_in(0) => n9, 
                           shift_out(63) => positive_inputs_19_63_port, 
                           shift_out(62) => positive_inputs_19_62_port, 
                           shift_out(61) => positive_inputs_19_61_port, 
                           shift_out(60) => positive_inputs_19_60_port, 
                           shift_out(59) => positive_inputs_19_59_port, 
                           shift_out(58) => positive_inputs_19_58_port, 
                           shift_out(57) => positive_inputs_19_57_port, 
                           shift_out(56) => positive_inputs_19_56_port, 
                           shift_out(55) => positive_inputs_19_55_port, 
                           shift_out(54) => positive_inputs_19_54_port, 
                           shift_out(53) => positive_inputs_19_53_port, 
                           shift_out(52) => positive_inputs_19_52_port, 
                           shift_out(51) => positive_inputs_19_51_port, 
                           shift_out(50) => positive_inputs_19_50_port, 
                           shift_out(49) => positive_inputs_19_49_port, 
                           shift_out(48) => positive_inputs_19_48_port, 
                           shift_out(47) => positive_inputs_19_47_port, 
                           shift_out(46) => positive_inputs_19_46_port, 
                           shift_out(45) => positive_inputs_19_45_port, 
                           shift_out(44) => positive_inputs_19_44_port, 
                           shift_out(43) => positive_inputs_19_43_port, 
                           shift_out(42) => positive_inputs_19_42_port, 
                           shift_out(41) => positive_inputs_19_41_port, 
                           shift_out(40) => positive_inputs_19_40_port, 
                           shift_out(39) => positive_inputs_19_39_port, 
                           shift_out(38) => positive_inputs_19_38_port, 
                           shift_out(37) => positive_inputs_19_37_port, 
                           shift_out(36) => positive_inputs_19_36_port, 
                           shift_out(35) => positive_inputs_19_35_port, 
                           shift_out(34) => positive_inputs_19_34_port, 
                           shift_out(33) => positive_inputs_19_33_port, 
                           shift_out(32) => positive_inputs_19_32_port, 
                           shift_out(31) => positive_inputs_19_31_port, 
                           shift_out(30) => positive_inputs_19_30_port, 
                           shift_out(29) => positive_inputs_19_29_port, 
                           shift_out(28) => positive_inputs_19_28_port, 
                           shift_out(27) => positive_inputs_19_27_port, 
                           shift_out(26) => positive_inputs_19_26_port, 
                           shift_out(25) => positive_inputs_19_25_port, 
                           shift_out(24) => positive_inputs_19_24_port, 
                           shift_out(23) => positive_inputs_19_23_port, 
                           shift_out(22) => positive_inputs_19_22_port, 
                           shift_out(21) => positive_inputs_19_21_port, 
                           shift_out(20) => positive_inputs_19_20_port, 
                           shift_out(19) => positive_inputs_19_19_port, 
                           shift_out(18) => positive_inputs_19_18_port, 
                           shift_out(17) => positive_inputs_19_17_port, 
                           shift_out(16) => positive_inputs_19_16_port, 
                           shift_out(15) => positive_inputs_19_15_port, 
                           shift_out(14) => positive_inputs_19_14_port, 
                           shift_out(13) => positive_inputs_19_13_port, 
                           shift_out(12) => positive_inputs_19_12_port, 
                           shift_out(11) => positive_inputs_19_11_port, 
                           shift_out(10) => positive_inputs_19_10_port, 
                           shift_out(9) => positive_inputs_19_9_port, 
                           shift_out(8) => positive_inputs_19_8_port, 
                           shift_out(7) => positive_inputs_19_7_port, 
                           shift_out(6) => positive_inputs_19_6_port, 
                           shift_out(5) => positive_inputs_19_5_port, 
                           shift_out(4) => positive_inputs_19_4_port, 
                           shift_out(3) => positive_inputs_19_3_port, 
                           shift_out(2) => positive_inputs_19_2_port, 
                           shift_out(1) => positive_inputs_19_1_port, 
                           shift_out(0) => n_1019);
   shifted_pos_20 : leftshifter_NbitShifter64_44 port map( shift_in(63) => 
                           positive_inputs_19_63_port, shift_in(62) => 
                           positive_inputs_19_62_port, shift_in(61) => 
                           positive_inputs_19_61_port, shift_in(60) => 
                           positive_inputs_19_60_port, shift_in(59) => 
                           positive_inputs_19_59_port, shift_in(58) => 
                           positive_inputs_19_58_port, shift_in(57) => 
                           positive_inputs_19_57_port, shift_in(56) => 
                           positive_inputs_19_56_port, shift_in(55) => 
                           positive_inputs_19_55_port, shift_in(54) => 
                           positive_inputs_19_54_port, shift_in(53) => 
                           positive_inputs_19_53_port, shift_in(52) => 
                           positive_inputs_19_52_port, shift_in(51) => 
                           positive_inputs_19_51_port, shift_in(50) => 
                           positive_inputs_19_50_port, shift_in(49) => 
                           positive_inputs_19_49_port, shift_in(48) => 
                           positive_inputs_19_48_port, shift_in(47) => 
                           positive_inputs_19_47_port, shift_in(46) => 
                           positive_inputs_19_46_port, shift_in(45) => 
                           positive_inputs_19_45_port, shift_in(44) => 
                           positive_inputs_19_44_port, shift_in(43) => 
                           positive_inputs_19_43_port, shift_in(42) => 
                           positive_inputs_19_42_port, shift_in(41) => 
                           positive_inputs_19_41_port, shift_in(40) => 
                           positive_inputs_19_40_port, shift_in(39) => 
                           positive_inputs_19_39_port, shift_in(38) => 
                           positive_inputs_19_38_port, shift_in(37) => 
                           positive_inputs_19_37_port, shift_in(36) => 
                           positive_inputs_19_36_port, shift_in(35) => 
                           positive_inputs_19_35_port, shift_in(34) => 
                           positive_inputs_19_34_port, shift_in(33) => 
                           positive_inputs_19_33_port, shift_in(32) => 
                           positive_inputs_19_32_port, shift_in(31) => 
                           positive_inputs_19_31_port, shift_in(30) => 
                           positive_inputs_19_30_port, shift_in(29) => 
                           positive_inputs_19_29_port, shift_in(28) => 
                           positive_inputs_19_28_port, shift_in(27) => 
                           positive_inputs_19_27_port, shift_in(26) => 
                           positive_inputs_19_26_port, shift_in(25) => 
                           positive_inputs_19_25_port, shift_in(24) => 
                           positive_inputs_19_24_port, shift_in(23) => 
                           positive_inputs_19_23_port, shift_in(22) => 
                           positive_inputs_19_22_port, shift_in(21) => 
                           positive_inputs_19_21_port, shift_in(20) => 
                           positive_inputs_19_20_port, shift_in(19) => 
                           positive_inputs_19_19_port, shift_in(18) => 
                           positive_inputs_19_18_port, shift_in(17) => 
                           positive_inputs_19_17_port, shift_in(16) => 
                           positive_inputs_19_16_port, shift_in(15) => 
                           positive_inputs_19_15_port, shift_in(14) => 
                           positive_inputs_19_14_port, shift_in(13) => 
                           positive_inputs_19_13_port, shift_in(12) => 
                           positive_inputs_19_12_port, shift_in(11) => 
                           positive_inputs_19_11_port, shift_in(10) => 
                           positive_inputs_19_10_port, shift_in(9) => 
                           positive_inputs_19_9_port, shift_in(8) => 
                           positive_inputs_19_8_port, shift_in(7) => 
                           positive_inputs_19_7_port, shift_in(6) => 
                           positive_inputs_19_6_port, shift_in(5) => 
                           positive_inputs_19_5_port, shift_in(4) => 
                           positive_inputs_19_4_port, shift_in(3) => 
                           positive_inputs_19_3_port, shift_in(2) => 
                           positive_inputs_19_2_port, shift_in(1) => 
                           positive_inputs_19_1_port, shift_in(0) => n9, 
                           shift_out(63) => positive_inputs_20_63_port, 
                           shift_out(62) => positive_inputs_20_62_port, 
                           shift_out(61) => positive_inputs_20_61_port, 
                           shift_out(60) => positive_inputs_20_60_port, 
                           shift_out(59) => positive_inputs_20_59_port, 
                           shift_out(58) => positive_inputs_20_58_port, 
                           shift_out(57) => positive_inputs_20_57_port, 
                           shift_out(56) => positive_inputs_20_56_port, 
                           shift_out(55) => positive_inputs_20_55_port, 
                           shift_out(54) => positive_inputs_20_54_port, 
                           shift_out(53) => positive_inputs_20_53_port, 
                           shift_out(52) => positive_inputs_20_52_port, 
                           shift_out(51) => positive_inputs_20_51_port, 
                           shift_out(50) => positive_inputs_20_50_port, 
                           shift_out(49) => positive_inputs_20_49_port, 
                           shift_out(48) => positive_inputs_20_48_port, 
                           shift_out(47) => positive_inputs_20_47_port, 
                           shift_out(46) => positive_inputs_20_46_port, 
                           shift_out(45) => positive_inputs_20_45_port, 
                           shift_out(44) => positive_inputs_20_44_port, 
                           shift_out(43) => positive_inputs_20_43_port, 
                           shift_out(42) => positive_inputs_20_42_port, 
                           shift_out(41) => positive_inputs_20_41_port, 
                           shift_out(40) => positive_inputs_20_40_port, 
                           shift_out(39) => positive_inputs_20_39_port, 
                           shift_out(38) => positive_inputs_20_38_port, 
                           shift_out(37) => positive_inputs_20_37_port, 
                           shift_out(36) => positive_inputs_20_36_port, 
                           shift_out(35) => positive_inputs_20_35_port, 
                           shift_out(34) => positive_inputs_20_34_port, 
                           shift_out(33) => positive_inputs_20_33_port, 
                           shift_out(32) => positive_inputs_20_32_port, 
                           shift_out(31) => positive_inputs_20_31_port, 
                           shift_out(30) => positive_inputs_20_30_port, 
                           shift_out(29) => positive_inputs_20_29_port, 
                           shift_out(28) => positive_inputs_20_28_port, 
                           shift_out(27) => positive_inputs_20_27_port, 
                           shift_out(26) => positive_inputs_20_26_port, 
                           shift_out(25) => positive_inputs_20_25_port, 
                           shift_out(24) => positive_inputs_20_24_port, 
                           shift_out(23) => positive_inputs_20_23_port, 
                           shift_out(22) => positive_inputs_20_22_port, 
                           shift_out(21) => positive_inputs_20_21_port, 
                           shift_out(20) => positive_inputs_20_20_port, 
                           shift_out(19) => positive_inputs_20_19_port, 
                           shift_out(18) => positive_inputs_20_18_port, 
                           shift_out(17) => positive_inputs_20_17_port, 
                           shift_out(16) => positive_inputs_20_16_port, 
                           shift_out(15) => positive_inputs_20_15_port, 
                           shift_out(14) => positive_inputs_20_14_port, 
                           shift_out(13) => positive_inputs_20_13_port, 
                           shift_out(12) => positive_inputs_20_12_port, 
                           shift_out(11) => positive_inputs_20_11_port, 
                           shift_out(10) => positive_inputs_20_10_port, 
                           shift_out(9) => positive_inputs_20_9_port, 
                           shift_out(8) => positive_inputs_20_8_port, 
                           shift_out(7) => positive_inputs_20_7_port, 
                           shift_out(6) => positive_inputs_20_6_port, 
                           shift_out(5) => positive_inputs_20_5_port, 
                           shift_out(4) => positive_inputs_20_4_port, 
                           shift_out(3) => positive_inputs_20_3_port, 
                           shift_out(2) => positive_inputs_20_2_port, 
                           shift_out(1) => positive_inputs_20_1_port, 
                           shift_out(0) => n_1020);
   shifted_pos_21 : leftshifter_NbitShifter64_43 port map( shift_in(63) => 
                           positive_inputs_20_63_port, shift_in(62) => 
                           positive_inputs_20_62_port, shift_in(61) => 
                           positive_inputs_20_61_port, shift_in(60) => 
                           positive_inputs_20_60_port, shift_in(59) => 
                           positive_inputs_20_59_port, shift_in(58) => 
                           positive_inputs_20_58_port, shift_in(57) => 
                           positive_inputs_20_57_port, shift_in(56) => 
                           positive_inputs_20_56_port, shift_in(55) => 
                           positive_inputs_20_55_port, shift_in(54) => 
                           positive_inputs_20_54_port, shift_in(53) => 
                           positive_inputs_20_53_port, shift_in(52) => 
                           positive_inputs_20_52_port, shift_in(51) => 
                           positive_inputs_20_51_port, shift_in(50) => 
                           positive_inputs_20_50_port, shift_in(49) => 
                           positive_inputs_20_49_port, shift_in(48) => 
                           positive_inputs_20_48_port, shift_in(47) => 
                           positive_inputs_20_47_port, shift_in(46) => 
                           positive_inputs_20_46_port, shift_in(45) => 
                           positive_inputs_20_45_port, shift_in(44) => 
                           positive_inputs_20_44_port, shift_in(43) => 
                           positive_inputs_20_43_port, shift_in(42) => 
                           positive_inputs_20_42_port, shift_in(41) => 
                           positive_inputs_20_41_port, shift_in(40) => 
                           positive_inputs_20_40_port, shift_in(39) => 
                           positive_inputs_20_39_port, shift_in(38) => 
                           positive_inputs_20_38_port, shift_in(37) => 
                           positive_inputs_20_37_port, shift_in(36) => 
                           positive_inputs_20_36_port, shift_in(35) => 
                           positive_inputs_20_35_port, shift_in(34) => 
                           positive_inputs_20_34_port, shift_in(33) => 
                           positive_inputs_20_33_port, shift_in(32) => 
                           positive_inputs_20_32_port, shift_in(31) => 
                           positive_inputs_20_31_port, shift_in(30) => 
                           positive_inputs_20_30_port, shift_in(29) => 
                           positive_inputs_20_29_port, shift_in(28) => 
                           positive_inputs_20_28_port, shift_in(27) => 
                           positive_inputs_20_27_port, shift_in(26) => 
                           positive_inputs_20_26_port, shift_in(25) => 
                           positive_inputs_20_25_port, shift_in(24) => 
                           positive_inputs_20_24_port, shift_in(23) => 
                           positive_inputs_20_23_port, shift_in(22) => 
                           positive_inputs_20_22_port, shift_in(21) => 
                           positive_inputs_20_21_port, shift_in(20) => 
                           positive_inputs_20_20_port, shift_in(19) => 
                           positive_inputs_20_19_port, shift_in(18) => 
                           positive_inputs_20_18_port, shift_in(17) => 
                           positive_inputs_20_17_port, shift_in(16) => 
                           positive_inputs_20_16_port, shift_in(15) => 
                           positive_inputs_20_15_port, shift_in(14) => 
                           positive_inputs_20_14_port, shift_in(13) => 
                           positive_inputs_20_13_port, shift_in(12) => 
                           positive_inputs_20_12_port, shift_in(11) => 
                           positive_inputs_20_11_port, shift_in(10) => 
                           positive_inputs_20_10_port, shift_in(9) => 
                           positive_inputs_20_9_port, shift_in(8) => 
                           positive_inputs_20_8_port, shift_in(7) => 
                           positive_inputs_20_7_port, shift_in(6) => 
                           positive_inputs_20_6_port, shift_in(5) => 
                           positive_inputs_20_5_port, shift_in(4) => 
                           positive_inputs_20_4_port, shift_in(3) => 
                           positive_inputs_20_3_port, shift_in(2) => 
                           positive_inputs_20_2_port, shift_in(1) => 
                           positive_inputs_20_1_port, shift_in(0) => n9, 
                           shift_out(63) => positive_inputs_21_63_port, 
                           shift_out(62) => positive_inputs_21_62_port, 
                           shift_out(61) => positive_inputs_21_61_port, 
                           shift_out(60) => positive_inputs_21_60_port, 
                           shift_out(59) => positive_inputs_21_59_port, 
                           shift_out(58) => positive_inputs_21_58_port, 
                           shift_out(57) => positive_inputs_21_57_port, 
                           shift_out(56) => positive_inputs_21_56_port, 
                           shift_out(55) => positive_inputs_21_55_port, 
                           shift_out(54) => positive_inputs_21_54_port, 
                           shift_out(53) => positive_inputs_21_53_port, 
                           shift_out(52) => positive_inputs_21_52_port, 
                           shift_out(51) => positive_inputs_21_51_port, 
                           shift_out(50) => positive_inputs_21_50_port, 
                           shift_out(49) => positive_inputs_21_49_port, 
                           shift_out(48) => positive_inputs_21_48_port, 
                           shift_out(47) => positive_inputs_21_47_port, 
                           shift_out(46) => positive_inputs_21_46_port, 
                           shift_out(45) => positive_inputs_21_45_port, 
                           shift_out(44) => positive_inputs_21_44_port, 
                           shift_out(43) => positive_inputs_21_43_port, 
                           shift_out(42) => positive_inputs_21_42_port, 
                           shift_out(41) => positive_inputs_21_41_port, 
                           shift_out(40) => positive_inputs_21_40_port, 
                           shift_out(39) => positive_inputs_21_39_port, 
                           shift_out(38) => positive_inputs_21_38_port, 
                           shift_out(37) => positive_inputs_21_37_port, 
                           shift_out(36) => positive_inputs_21_36_port, 
                           shift_out(35) => positive_inputs_21_35_port, 
                           shift_out(34) => positive_inputs_21_34_port, 
                           shift_out(33) => positive_inputs_21_33_port, 
                           shift_out(32) => positive_inputs_21_32_port, 
                           shift_out(31) => positive_inputs_21_31_port, 
                           shift_out(30) => positive_inputs_21_30_port, 
                           shift_out(29) => positive_inputs_21_29_port, 
                           shift_out(28) => positive_inputs_21_28_port, 
                           shift_out(27) => positive_inputs_21_27_port, 
                           shift_out(26) => positive_inputs_21_26_port, 
                           shift_out(25) => positive_inputs_21_25_port, 
                           shift_out(24) => positive_inputs_21_24_port, 
                           shift_out(23) => positive_inputs_21_23_port, 
                           shift_out(22) => positive_inputs_21_22_port, 
                           shift_out(21) => positive_inputs_21_21_port, 
                           shift_out(20) => positive_inputs_21_20_port, 
                           shift_out(19) => positive_inputs_21_19_port, 
                           shift_out(18) => positive_inputs_21_18_port, 
                           shift_out(17) => positive_inputs_21_17_port, 
                           shift_out(16) => positive_inputs_21_16_port, 
                           shift_out(15) => positive_inputs_21_15_port, 
                           shift_out(14) => positive_inputs_21_14_port, 
                           shift_out(13) => positive_inputs_21_13_port, 
                           shift_out(12) => positive_inputs_21_12_port, 
                           shift_out(11) => positive_inputs_21_11_port, 
                           shift_out(10) => positive_inputs_21_10_port, 
                           shift_out(9) => positive_inputs_21_9_port, 
                           shift_out(8) => positive_inputs_21_8_port, 
                           shift_out(7) => positive_inputs_21_7_port, 
                           shift_out(6) => positive_inputs_21_6_port, 
                           shift_out(5) => positive_inputs_21_5_port, 
                           shift_out(4) => positive_inputs_21_4_port, 
                           shift_out(3) => positive_inputs_21_3_port, 
                           shift_out(2) => positive_inputs_21_2_port, 
                           shift_out(1) => positive_inputs_21_1_port, 
                           shift_out(0) => n_1021);
   shifted_pos_22 : leftshifter_NbitShifter64_42 port map( shift_in(63) => 
                           positive_inputs_21_63_port, shift_in(62) => 
                           positive_inputs_21_62_port, shift_in(61) => 
                           positive_inputs_21_61_port, shift_in(60) => 
                           positive_inputs_21_60_port, shift_in(59) => 
                           positive_inputs_21_59_port, shift_in(58) => 
                           positive_inputs_21_58_port, shift_in(57) => 
                           positive_inputs_21_57_port, shift_in(56) => 
                           positive_inputs_21_56_port, shift_in(55) => 
                           positive_inputs_21_55_port, shift_in(54) => 
                           positive_inputs_21_54_port, shift_in(53) => 
                           positive_inputs_21_53_port, shift_in(52) => 
                           positive_inputs_21_52_port, shift_in(51) => 
                           positive_inputs_21_51_port, shift_in(50) => 
                           positive_inputs_21_50_port, shift_in(49) => 
                           positive_inputs_21_49_port, shift_in(48) => 
                           positive_inputs_21_48_port, shift_in(47) => 
                           positive_inputs_21_47_port, shift_in(46) => 
                           positive_inputs_21_46_port, shift_in(45) => 
                           positive_inputs_21_45_port, shift_in(44) => 
                           positive_inputs_21_44_port, shift_in(43) => 
                           positive_inputs_21_43_port, shift_in(42) => 
                           positive_inputs_21_42_port, shift_in(41) => 
                           positive_inputs_21_41_port, shift_in(40) => 
                           positive_inputs_21_40_port, shift_in(39) => 
                           positive_inputs_21_39_port, shift_in(38) => 
                           positive_inputs_21_38_port, shift_in(37) => 
                           positive_inputs_21_37_port, shift_in(36) => 
                           positive_inputs_21_36_port, shift_in(35) => 
                           positive_inputs_21_35_port, shift_in(34) => 
                           positive_inputs_21_34_port, shift_in(33) => 
                           positive_inputs_21_33_port, shift_in(32) => 
                           positive_inputs_21_32_port, shift_in(31) => 
                           positive_inputs_21_31_port, shift_in(30) => 
                           positive_inputs_21_30_port, shift_in(29) => 
                           positive_inputs_21_29_port, shift_in(28) => 
                           positive_inputs_21_28_port, shift_in(27) => 
                           positive_inputs_21_27_port, shift_in(26) => 
                           positive_inputs_21_26_port, shift_in(25) => 
                           positive_inputs_21_25_port, shift_in(24) => 
                           positive_inputs_21_24_port, shift_in(23) => 
                           positive_inputs_21_23_port, shift_in(22) => 
                           positive_inputs_21_22_port, shift_in(21) => 
                           positive_inputs_21_21_port, shift_in(20) => 
                           positive_inputs_21_20_port, shift_in(19) => 
                           positive_inputs_21_19_port, shift_in(18) => 
                           positive_inputs_21_18_port, shift_in(17) => 
                           positive_inputs_21_17_port, shift_in(16) => 
                           positive_inputs_21_16_port, shift_in(15) => 
                           positive_inputs_21_15_port, shift_in(14) => 
                           positive_inputs_21_14_port, shift_in(13) => 
                           positive_inputs_21_13_port, shift_in(12) => 
                           positive_inputs_21_12_port, shift_in(11) => 
                           positive_inputs_21_11_port, shift_in(10) => 
                           positive_inputs_21_10_port, shift_in(9) => 
                           positive_inputs_21_9_port, shift_in(8) => 
                           positive_inputs_21_8_port, shift_in(7) => 
                           positive_inputs_21_7_port, shift_in(6) => 
                           positive_inputs_21_6_port, shift_in(5) => 
                           positive_inputs_21_5_port, shift_in(4) => 
                           positive_inputs_21_4_port, shift_in(3) => 
                           positive_inputs_21_3_port, shift_in(2) => 
                           positive_inputs_21_2_port, shift_in(1) => 
                           positive_inputs_21_1_port, shift_in(0) => n9, 
                           shift_out(63) => positive_inputs_22_63_port, 
                           shift_out(62) => positive_inputs_22_62_port, 
                           shift_out(61) => positive_inputs_22_61_port, 
                           shift_out(60) => positive_inputs_22_60_port, 
                           shift_out(59) => positive_inputs_22_59_port, 
                           shift_out(58) => positive_inputs_22_58_port, 
                           shift_out(57) => positive_inputs_22_57_port, 
                           shift_out(56) => positive_inputs_22_56_port, 
                           shift_out(55) => positive_inputs_22_55_port, 
                           shift_out(54) => positive_inputs_22_54_port, 
                           shift_out(53) => positive_inputs_22_53_port, 
                           shift_out(52) => positive_inputs_22_52_port, 
                           shift_out(51) => positive_inputs_22_51_port, 
                           shift_out(50) => positive_inputs_22_50_port, 
                           shift_out(49) => positive_inputs_22_49_port, 
                           shift_out(48) => positive_inputs_22_48_port, 
                           shift_out(47) => positive_inputs_22_47_port, 
                           shift_out(46) => positive_inputs_22_46_port, 
                           shift_out(45) => positive_inputs_22_45_port, 
                           shift_out(44) => positive_inputs_22_44_port, 
                           shift_out(43) => positive_inputs_22_43_port, 
                           shift_out(42) => positive_inputs_22_42_port, 
                           shift_out(41) => positive_inputs_22_41_port, 
                           shift_out(40) => positive_inputs_22_40_port, 
                           shift_out(39) => positive_inputs_22_39_port, 
                           shift_out(38) => positive_inputs_22_38_port, 
                           shift_out(37) => positive_inputs_22_37_port, 
                           shift_out(36) => positive_inputs_22_36_port, 
                           shift_out(35) => positive_inputs_22_35_port, 
                           shift_out(34) => positive_inputs_22_34_port, 
                           shift_out(33) => positive_inputs_22_33_port, 
                           shift_out(32) => positive_inputs_22_32_port, 
                           shift_out(31) => positive_inputs_22_31_port, 
                           shift_out(30) => positive_inputs_22_30_port, 
                           shift_out(29) => positive_inputs_22_29_port, 
                           shift_out(28) => positive_inputs_22_28_port, 
                           shift_out(27) => positive_inputs_22_27_port, 
                           shift_out(26) => positive_inputs_22_26_port, 
                           shift_out(25) => positive_inputs_22_25_port, 
                           shift_out(24) => positive_inputs_22_24_port, 
                           shift_out(23) => positive_inputs_22_23_port, 
                           shift_out(22) => positive_inputs_22_22_port, 
                           shift_out(21) => positive_inputs_22_21_port, 
                           shift_out(20) => positive_inputs_22_20_port, 
                           shift_out(19) => positive_inputs_22_19_port, 
                           shift_out(18) => positive_inputs_22_18_port, 
                           shift_out(17) => positive_inputs_22_17_port, 
                           shift_out(16) => positive_inputs_22_16_port, 
                           shift_out(15) => positive_inputs_22_15_port, 
                           shift_out(14) => positive_inputs_22_14_port, 
                           shift_out(13) => positive_inputs_22_13_port, 
                           shift_out(12) => positive_inputs_22_12_port, 
                           shift_out(11) => positive_inputs_22_11_port, 
                           shift_out(10) => positive_inputs_22_10_port, 
                           shift_out(9) => positive_inputs_22_9_port, 
                           shift_out(8) => positive_inputs_22_8_port, 
                           shift_out(7) => positive_inputs_22_7_port, 
                           shift_out(6) => positive_inputs_22_6_port, 
                           shift_out(5) => positive_inputs_22_5_port, 
                           shift_out(4) => positive_inputs_22_4_port, 
                           shift_out(3) => positive_inputs_22_3_port, 
                           shift_out(2) => positive_inputs_22_2_port, 
                           shift_out(1) => positive_inputs_22_1_port, 
                           shift_out(0) => n_1022);
   shifted_pos_23 : leftshifter_NbitShifter64_41 port map( shift_in(63) => 
                           positive_inputs_22_63_port, shift_in(62) => 
                           positive_inputs_22_62_port, shift_in(61) => 
                           positive_inputs_22_61_port, shift_in(60) => 
                           positive_inputs_22_60_port, shift_in(59) => 
                           positive_inputs_22_59_port, shift_in(58) => 
                           positive_inputs_22_58_port, shift_in(57) => 
                           positive_inputs_22_57_port, shift_in(56) => 
                           positive_inputs_22_56_port, shift_in(55) => 
                           positive_inputs_22_55_port, shift_in(54) => 
                           positive_inputs_22_54_port, shift_in(53) => 
                           positive_inputs_22_53_port, shift_in(52) => 
                           positive_inputs_22_52_port, shift_in(51) => 
                           positive_inputs_22_51_port, shift_in(50) => 
                           positive_inputs_22_50_port, shift_in(49) => 
                           positive_inputs_22_49_port, shift_in(48) => 
                           positive_inputs_22_48_port, shift_in(47) => 
                           positive_inputs_22_47_port, shift_in(46) => 
                           positive_inputs_22_46_port, shift_in(45) => 
                           positive_inputs_22_45_port, shift_in(44) => 
                           positive_inputs_22_44_port, shift_in(43) => 
                           positive_inputs_22_43_port, shift_in(42) => 
                           positive_inputs_22_42_port, shift_in(41) => 
                           positive_inputs_22_41_port, shift_in(40) => 
                           positive_inputs_22_40_port, shift_in(39) => 
                           positive_inputs_22_39_port, shift_in(38) => 
                           positive_inputs_22_38_port, shift_in(37) => 
                           positive_inputs_22_37_port, shift_in(36) => 
                           positive_inputs_22_36_port, shift_in(35) => 
                           positive_inputs_22_35_port, shift_in(34) => 
                           positive_inputs_22_34_port, shift_in(33) => 
                           positive_inputs_22_33_port, shift_in(32) => 
                           positive_inputs_22_32_port, shift_in(31) => 
                           positive_inputs_22_31_port, shift_in(30) => 
                           positive_inputs_22_30_port, shift_in(29) => 
                           positive_inputs_22_29_port, shift_in(28) => 
                           positive_inputs_22_28_port, shift_in(27) => 
                           positive_inputs_22_27_port, shift_in(26) => 
                           positive_inputs_22_26_port, shift_in(25) => 
                           positive_inputs_22_25_port, shift_in(24) => 
                           positive_inputs_22_24_port, shift_in(23) => 
                           positive_inputs_22_23_port, shift_in(22) => 
                           positive_inputs_22_22_port, shift_in(21) => 
                           positive_inputs_22_21_port, shift_in(20) => 
                           positive_inputs_22_20_port, shift_in(19) => 
                           positive_inputs_22_19_port, shift_in(18) => 
                           positive_inputs_22_18_port, shift_in(17) => 
                           positive_inputs_22_17_port, shift_in(16) => 
                           positive_inputs_22_16_port, shift_in(15) => 
                           positive_inputs_22_15_port, shift_in(14) => 
                           positive_inputs_22_14_port, shift_in(13) => 
                           positive_inputs_22_13_port, shift_in(12) => 
                           positive_inputs_22_12_port, shift_in(11) => 
                           positive_inputs_22_11_port, shift_in(10) => 
                           positive_inputs_22_10_port, shift_in(9) => 
                           positive_inputs_22_9_port, shift_in(8) => 
                           positive_inputs_22_8_port, shift_in(7) => 
                           positive_inputs_22_7_port, shift_in(6) => 
                           positive_inputs_22_6_port, shift_in(5) => 
                           positive_inputs_22_5_port, shift_in(4) => 
                           positive_inputs_22_4_port, shift_in(3) => 
                           positive_inputs_22_3_port, shift_in(2) => 
                           positive_inputs_22_2_port, shift_in(1) => 
                           positive_inputs_22_1_port, shift_in(0) => n9, 
                           shift_out(63) => positive_inputs_23_63_port, 
                           shift_out(62) => positive_inputs_23_62_port, 
                           shift_out(61) => positive_inputs_23_61_port, 
                           shift_out(60) => positive_inputs_23_60_port, 
                           shift_out(59) => positive_inputs_23_59_port, 
                           shift_out(58) => positive_inputs_23_58_port, 
                           shift_out(57) => positive_inputs_23_57_port, 
                           shift_out(56) => positive_inputs_23_56_port, 
                           shift_out(55) => positive_inputs_23_55_port, 
                           shift_out(54) => positive_inputs_23_54_port, 
                           shift_out(53) => positive_inputs_23_53_port, 
                           shift_out(52) => positive_inputs_23_52_port, 
                           shift_out(51) => positive_inputs_23_51_port, 
                           shift_out(50) => positive_inputs_23_50_port, 
                           shift_out(49) => positive_inputs_23_49_port, 
                           shift_out(48) => positive_inputs_23_48_port, 
                           shift_out(47) => positive_inputs_23_47_port, 
                           shift_out(46) => positive_inputs_23_46_port, 
                           shift_out(45) => positive_inputs_23_45_port, 
                           shift_out(44) => positive_inputs_23_44_port, 
                           shift_out(43) => positive_inputs_23_43_port, 
                           shift_out(42) => positive_inputs_23_42_port, 
                           shift_out(41) => positive_inputs_23_41_port, 
                           shift_out(40) => positive_inputs_23_40_port, 
                           shift_out(39) => positive_inputs_23_39_port, 
                           shift_out(38) => positive_inputs_23_38_port, 
                           shift_out(37) => positive_inputs_23_37_port, 
                           shift_out(36) => positive_inputs_23_36_port, 
                           shift_out(35) => positive_inputs_23_35_port, 
                           shift_out(34) => positive_inputs_23_34_port, 
                           shift_out(33) => positive_inputs_23_33_port, 
                           shift_out(32) => positive_inputs_23_32_port, 
                           shift_out(31) => positive_inputs_23_31_port, 
                           shift_out(30) => positive_inputs_23_30_port, 
                           shift_out(29) => positive_inputs_23_29_port, 
                           shift_out(28) => positive_inputs_23_28_port, 
                           shift_out(27) => positive_inputs_23_27_port, 
                           shift_out(26) => positive_inputs_23_26_port, 
                           shift_out(25) => positive_inputs_23_25_port, 
                           shift_out(24) => positive_inputs_23_24_port, 
                           shift_out(23) => positive_inputs_23_23_port, 
                           shift_out(22) => positive_inputs_23_22_port, 
                           shift_out(21) => positive_inputs_23_21_port, 
                           shift_out(20) => positive_inputs_23_20_port, 
                           shift_out(19) => positive_inputs_23_19_port, 
                           shift_out(18) => positive_inputs_23_18_port, 
                           shift_out(17) => positive_inputs_23_17_port, 
                           shift_out(16) => positive_inputs_23_16_port, 
                           shift_out(15) => positive_inputs_23_15_port, 
                           shift_out(14) => positive_inputs_23_14_port, 
                           shift_out(13) => positive_inputs_23_13_port, 
                           shift_out(12) => positive_inputs_23_12_port, 
                           shift_out(11) => positive_inputs_23_11_port, 
                           shift_out(10) => positive_inputs_23_10_port, 
                           shift_out(9) => positive_inputs_23_9_port, 
                           shift_out(8) => positive_inputs_23_8_port, 
                           shift_out(7) => positive_inputs_23_7_port, 
                           shift_out(6) => positive_inputs_23_6_port, 
                           shift_out(5) => positive_inputs_23_5_port, 
                           shift_out(4) => positive_inputs_23_4_port, 
                           shift_out(3) => positive_inputs_23_3_port, 
                           shift_out(2) => positive_inputs_23_2_port, 
                           shift_out(1) => positive_inputs_23_1_port, 
                           shift_out(0) => n_1023);
   shifted_pos_24 : leftshifter_NbitShifter64_40 port map( shift_in(63) => 
                           positive_inputs_23_63_port, shift_in(62) => 
                           positive_inputs_23_62_port, shift_in(61) => 
                           positive_inputs_23_61_port, shift_in(60) => 
                           positive_inputs_23_60_port, shift_in(59) => 
                           positive_inputs_23_59_port, shift_in(58) => 
                           positive_inputs_23_58_port, shift_in(57) => 
                           positive_inputs_23_57_port, shift_in(56) => 
                           positive_inputs_23_56_port, shift_in(55) => 
                           positive_inputs_23_55_port, shift_in(54) => 
                           positive_inputs_23_54_port, shift_in(53) => 
                           positive_inputs_23_53_port, shift_in(52) => 
                           positive_inputs_23_52_port, shift_in(51) => 
                           positive_inputs_23_51_port, shift_in(50) => 
                           positive_inputs_23_50_port, shift_in(49) => 
                           positive_inputs_23_49_port, shift_in(48) => 
                           positive_inputs_23_48_port, shift_in(47) => 
                           positive_inputs_23_47_port, shift_in(46) => 
                           positive_inputs_23_46_port, shift_in(45) => 
                           positive_inputs_23_45_port, shift_in(44) => 
                           positive_inputs_23_44_port, shift_in(43) => 
                           positive_inputs_23_43_port, shift_in(42) => 
                           positive_inputs_23_42_port, shift_in(41) => 
                           positive_inputs_23_41_port, shift_in(40) => 
                           positive_inputs_23_40_port, shift_in(39) => 
                           positive_inputs_23_39_port, shift_in(38) => 
                           positive_inputs_23_38_port, shift_in(37) => 
                           positive_inputs_23_37_port, shift_in(36) => 
                           positive_inputs_23_36_port, shift_in(35) => 
                           positive_inputs_23_35_port, shift_in(34) => 
                           positive_inputs_23_34_port, shift_in(33) => 
                           positive_inputs_23_33_port, shift_in(32) => 
                           positive_inputs_23_32_port, shift_in(31) => 
                           positive_inputs_23_31_port, shift_in(30) => 
                           positive_inputs_23_30_port, shift_in(29) => 
                           positive_inputs_23_29_port, shift_in(28) => 
                           positive_inputs_23_28_port, shift_in(27) => 
                           positive_inputs_23_27_port, shift_in(26) => 
                           positive_inputs_23_26_port, shift_in(25) => 
                           positive_inputs_23_25_port, shift_in(24) => 
                           positive_inputs_23_24_port, shift_in(23) => 
                           positive_inputs_23_23_port, shift_in(22) => 
                           positive_inputs_23_22_port, shift_in(21) => 
                           positive_inputs_23_21_port, shift_in(20) => 
                           positive_inputs_23_20_port, shift_in(19) => 
                           positive_inputs_23_19_port, shift_in(18) => 
                           positive_inputs_23_18_port, shift_in(17) => 
                           positive_inputs_23_17_port, shift_in(16) => 
                           positive_inputs_23_16_port, shift_in(15) => 
                           positive_inputs_23_15_port, shift_in(14) => 
                           positive_inputs_23_14_port, shift_in(13) => 
                           positive_inputs_23_13_port, shift_in(12) => 
                           positive_inputs_23_12_port, shift_in(11) => 
                           positive_inputs_23_11_port, shift_in(10) => 
                           positive_inputs_23_10_port, shift_in(9) => 
                           positive_inputs_23_9_port, shift_in(8) => 
                           positive_inputs_23_8_port, shift_in(7) => 
                           positive_inputs_23_7_port, shift_in(6) => 
                           positive_inputs_23_6_port, shift_in(5) => 
                           positive_inputs_23_5_port, shift_in(4) => 
                           positive_inputs_23_4_port, shift_in(3) => 
                           positive_inputs_23_3_port, shift_in(2) => 
                           positive_inputs_23_2_port, shift_in(1) => 
                           positive_inputs_23_1_port, shift_in(0) => n9, 
                           shift_out(63) => positive_inputs_24_63_port, 
                           shift_out(62) => positive_inputs_24_62_port, 
                           shift_out(61) => positive_inputs_24_61_port, 
                           shift_out(60) => positive_inputs_24_60_port, 
                           shift_out(59) => positive_inputs_24_59_port, 
                           shift_out(58) => positive_inputs_24_58_port, 
                           shift_out(57) => positive_inputs_24_57_port, 
                           shift_out(56) => positive_inputs_24_56_port, 
                           shift_out(55) => positive_inputs_24_55_port, 
                           shift_out(54) => positive_inputs_24_54_port, 
                           shift_out(53) => positive_inputs_24_53_port, 
                           shift_out(52) => positive_inputs_24_52_port, 
                           shift_out(51) => positive_inputs_24_51_port, 
                           shift_out(50) => positive_inputs_24_50_port, 
                           shift_out(49) => positive_inputs_24_49_port, 
                           shift_out(48) => positive_inputs_24_48_port, 
                           shift_out(47) => positive_inputs_24_47_port, 
                           shift_out(46) => positive_inputs_24_46_port, 
                           shift_out(45) => positive_inputs_24_45_port, 
                           shift_out(44) => positive_inputs_24_44_port, 
                           shift_out(43) => positive_inputs_24_43_port, 
                           shift_out(42) => positive_inputs_24_42_port, 
                           shift_out(41) => positive_inputs_24_41_port, 
                           shift_out(40) => positive_inputs_24_40_port, 
                           shift_out(39) => positive_inputs_24_39_port, 
                           shift_out(38) => positive_inputs_24_38_port, 
                           shift_out(37) => positive_inputs_24_37_port, 
                           shift_out(36) => positive_inputs_24_36_port, 
                           shift_out(35) => positive_inputs_24_35_port, 
                           shift_out(34) => positive_inputs_24_34_port, 
                           shift_out(33) => positive_inputs_24_33_port, 
                           shift_out(32) => positive_inputs_24_32_port, 
                           shift_out(31) => positive_inputs_24_31_port, 
                           shift_out(30) => positive_inputs_24_30_port, 
                           shift_out(29) => positive_inputs_24_29_port, 
                           shift_out(28) => positive_inputs_24_28_port, 
                           shift_out(27) => positive_inputs_24_27_port, 
                           shift_out(26) => positive_inputs_24_26_port, 
                           shift_out(25) => positive_inputs_24_25_port, 
                           shift_out(24) => positive_inputs_24_24_port, 
                           shift_out(23) => positive_inputs_24_23_port, 
                           shift_out(22) => positive_inputs_24_22_port, 
                           shift_out(21) => positive_inputs_24_21_port, 
                           shift_out(20) => positive_inputs_24_20_port, 
                           shift_out(19) => positive_inputs_24_19_port, 
                           shift_out(18) => positive_inputs_24_18_port, 
                           shift_out(17) => positive_inputs_24_17_port, 
                           shift_out(16) => positive_inputs_24_16_port, 
                           shift_out(15) => positive_inputs_24_15_port, 
                           shift_out(14) => positive_inputs_24_14_port, 
                           shift_out(13) => positive_inputs_24_13_port, 
                           shift_out(12) => positive_inputs_24_12_port, 
                           shift_out(11) => positive_inputs_24_11_port, 
                           shift_out(10) => positive_inputs_24_10_port, 
                           shift_out(9) => positive_inputs_24_9_port, 
                           shift_out(8) => positive_inputs_24_8_port, 
                           shift_out(7) => positive_inputs_24_7_port, 
                           shift_out(6) => positive_inputs_24_6_port, 
                           shift_out(5) => positive_inputs_24_5_port, 
                           shift_out(4) => positive_inputs_24_4_port, 
                           shift_out(3) => positive_inputs_24_3_port, 
                           shift_out(2) => positive_inputs_24_2_port, 
                           shift_out(1) => positive_inputs_24_1_port, 
                           shift_out(0) => n_1024);
   shifted_pos_25 : leftshifter_NbitShifter64_39 port map( shift_in(63) => 
                           positive_inputs_24_63_port, shift_in(62) => 
                           positive_inputs_24_62_port, shift_in(61) => 
                           positive_inputs_24_61_port, shift_in(60) => 
                           positive_inputs_24_60_port, shift_in(59) => 
                           positive_inputs_24_59_port, shift_in(58) => 
                           positive_inputs_24_58_port, shift_in(57) => 
                           positive_inputs_24_57_port, shift_in(56) => 
                           positive_inputs_24_56_port, shift_in(55) => 
                           positive_inputs_24_55_port, shift_in(54) => 
                           positive_inputs_24_54_port, shift_in(53) => 
                           positive_inputs_24_53_port, shift_in(52) => 
                           positive_inputs_24_52_port, shift_in(51) => 
                           positive_inputs_24_51_port, shift_in(50) => 
                           positive_inputs_24_50_port, shift_in(49) => 
                           positive_inputs_24_49_port, shift_in(48) => 
                           positive_inputs_24_48_port, shift_in(47) => 
                           positive_inputs_24_47_port, shift_in(46) => 
                           positive_inputs_24_46_port, shift_in(45) => 
                           positive_inputs_24_45_port, shift_in(44) => 
                           positive_inputs_24_44_port, shift_in(43) => 
                           positive_inputs_24_43_port, shift_in(42) => 
                           positive_inputs_24_42_port, shift_in(41) => 
                           positive_inputs_24_41_port, shift_in(40) => 
                           positive_inputs_24_40_port, shift_in(39) => 
                           positive_inputs_24_39_port, shift_in(38) => 
                           positive_inputs_24_38_port, shift_in(37) => 
                           positive_inputs_24_37_port, shift_in(36) => 
                           positive_inputs_24_36_port, shift_in(35) => 
                           positive_inputs_24_35_port, shift_in(34) => 
                           positive_inputs_24_34_port, shift_in(33) => 
                           positive_inputs_24_33_port, shift_in(32) => 
                           positive_inputs_24_32_port, shift_in(31) => 
                           positive_inputs_24_31_port, shift_in(30) => 
                           positive_inputs_24_30_port, shift_in(29) => 
                           positive_inputs_24_29_port, shift_in(28) => 
                           positive_inputs_24_28_port, shift_in(27) => 
                           positive_inputs_24_27_port, shift_in(26) => 
                           positive_inputs_24_26_port, shift_in(25) => 
                           positive_inputs_24_25_port, shift_in(24) => 
                           positive_inputs_24_24_port, shift_in(23) => 
                           positive_inputs_24_23_port, shift_in(22) => 
                           positive_inputs_24_22_port, shift_in(21) => 
                           positive_inputs_24_21_port, shift_in(20) => 
                           positive_inputs_24_20_port, shift_in(19) => 
                           positive_inputs_24_19_port, shift_in(18) => 
                           positive_inputs_24_18_port, shift_in(17) => 
                           positive_inputs_24_17_port, shift_in(16) => 
                           positive_inputs_24_16_port, shift_in(15) => 
                           positive_inputs_24_15_port, shift_in(14) => 
                           positive_inputs_24_14_port, shift_in(13) => 
                           positive_inputs_24_13_port, shift_in(12) => 
                           positive_inputs_24_12_port, shift_in(11) => 
                           positive_inputs_24_11_port, shift_in(10) => 
                           positive_inputs_24_10_port, shift_in(9) => 
                           positive_inputs_24_9_port, shift_in(8) => 
                           positive_inputs_24_8_port, shift_in(7) => 
                           positive_inputs_24_7_port, shift_in(6) => 
                           positive_inputs_24_6_port, shift_in(5) => 
                           positive_inputs_24_5_port, shift_in(4) => 
                           positive_inputs_24_4_port, shift_in(3) => 
                           positive_inputs_24_3_port, shift_in(2) => 
                           positive_inputs_24_2_port, shift_in(1) => 
                           positive_inputs_24_1_port, shift_in(0) => n9, 
                           shift_out(63) => positive_inputs_25_63_port, 
                           shift_out(62) => positive_inputs_25_62_port, 
                           shift_out(61) => positive_inputs_25_61_port, 
                           shift_out(60) => positive_inputs_25_60_port, 
                           shift_out(59) => positive_inputs_25_59_port, 
                           shift_out(58) => positive_inputs_25_58_port, 
                           shift_out(57) => positive_inputs_25_57_port, 
                           shift_out(56) => positive_inputs_25_56_port, 
                           shift_out(55) => positive_inputs_25_55_port, 
                           shift_out(54) => positive_inputs_25_54_port, 
                           shift_out(53) => positive_inputs_25_53_port, 
                           shift_out(52) => positive_inputs_25_52_port, 
                           shift_out(51) => positive_inputs_25_51_port, 
                           shift_out(50) => positive_inputs_25_50_port, 
                           shift_out(49) => positive_inputs_25_49_port, 
                           shift_out(48) => positive_inputs_25_48_port, 
                           shift_out(47) => positive_inputs_25_47_port, 
                           shift_out(46) => positive_inputs_25_46_port, 
                           shift_out(45) => positive_inputs_25_45_port, 
                           shift_out(44) => positive_inputs_25_44_port, 
                           shift_out(43) => positive_inputs_25_43_port, 
                           shift_out(42) => positive_inputs_25_42_port, 
                           shift_out(41) => positive_inputs_25_41_port, 
                           shift_out(40) => positive_inputs_25_40_port, 
                           shift_out(39) => positive_inputs_25_39_port, 
                           shift_out(38) => positive_inputs_25_38_port, 
                           shift_out(37) => positive_inputs_25_37_port, 
                           shift_out(36) => positive_inputs_25_36_port, 
                           shift_out(35) => positive_inputs_25_35_port, 
                           shift_out(34) => positive_inputs_25_34_port, 
                           shift_out(33) => positive_inputs_25_33_port, 
                           shift_out(32) => positive_inputs_25_32_port, 
                           shift_out(31) => positive_inputs_25_31_port, 
                           shift_out(30) => positive_inputs_25_30_port, 
                           shift_out(29) => positive_inputs_25_29_port, 
                           shift_out(28) => positive_inputs_25_28_port, 
                           shift_out(27) => positive_inputs_25_27_port, 
                           shift_out(26) => positive_inputs_25_26_port, 
                           shift_out(25) => positive_inputs_25_25_port, 
                           shift_out(24) => positive_inputs_25_24_port, 
                           shift_out(23) => positive_inputs_25_23_port, 
                           shift_out(22) => positive_inputs_25_22_port, 
                           shift_out(21) => positive_inputs_25_21_port, 
                           shift_out(20) => positive_inputs_25_20_port, 
                           shift_out(19) => positive_inputs_25_19_port, 
                           shift_out(18) => positive_inputs_25_18_port, 
                           shift_out(17) => positive_inputs_25_17_port, 
                           shift_out(16) => positive_inputs_25_16_port, 
                           shift_out(15) => positive_inputs_25_15_port, 
                           shift_out(14) => positive_inputs_25_14_port, 
                           shift_out(13) => positive_inputs_25_13_port, 
                           shift_out(12) => positive_inputs_25_12_port, 
                           shift_out(11) => positive_inputs_25_11_port, 
                           shift_out(10) => positive_inputs_25_10_port, 
                           shift_out(9) => positive_inputs_25_9_port, 
                           shift_out(8) => positive_inputs_25_8_port, 
                           shift_out(7) => positive_inputs_25_7_port, 
                           shift_out(6) => positive_inputs_25_6_port, 
                           shift_out(5) => positive_inputs_25_5_port, 
                           shift_out(4) => positive_inputs_25_4_port, 
                           shift_out(3) => positive_inputs_25_3_port, 
                           shift_out(2) => positive_inputs_25_2_port, 
                           shift_out(1) => positive_inputs_25_1_port, 
                           shift_out(0) => n_1025);
   shifted_pos_26 : leftshifter_NbitShifter64_38 port map( shift_in(63) => 
                           positive_inputs_25_63_port, shift_in(62) => 
                           positive_inputs_25_62_port, shift_in(61) => 
                           positive_inputs_25_61_port, shift_in(60) => 
                           positive_inputs_25_60_port, shift_in(59) => 
                           positive_inputs_25_59_port, shift_in(58) => 
                           positive_inputs_25_58_port, shift_in(57) => 
                           positive_inputs_25_57_port, shift_in(56) => 
                           positive_inputs_25_56_port, shift_in(55) => 
                           positive_inputs_25_55_port, shift_in(54) => 
                           positive_inputs_25_54_port, shift_in(53) => 
                           positive_inputs_25_53_port, shift_in(52) => 
                           positive_inputs_25_52_port, shift_in(51) => 
                           positive_inputs_25_51_port, shift_in(50) => 
                           positive_inputs_25_50_port, shift_in(49) => 
                           positive_inputs_25_49_port, shift_in(48) => 
                           positive_inputs_25_48_port, shift_in(47) => 
                           positive_inputs_25_47_port, shift_in(46) => 
                           positive_inputs_25_46_port, shift_in(45) => 
                           positive_inputs_25_45_port, shift_in(44) => 
                           positive_inputs_25_44_port, shift_in(43) => 
                           positive_inputs_25_43_port, shift_in(42) => 
                           positive_inputs_25_42_port, shift_in(41) => 
                           positive_inputs_25_41_port, shift_in(40) => 
                           positive_inputs_25_40_port, shift_in(39) => 
                           positive_inputs_25_39_port, shift_in(38) => 
                           positive_inputs_25_38_port, shift_in(37) => 
                           positive_inputs_25_37_port, shift_in(36) => 
                           positive_inputs_25_36_port, shift_in(35) => 
                           positive_inputs_25_35_port, shift_in(34) => 
                           positive_inputs_25_34_port, shift_in(33) => 
                           positive_inputs_25_33_port, shift_in(32) => 
                           positive_inputs_25_32_port, shift_in(31) => 
                           positive_inputs_25_31_port, shift_in(30) => 
                           positive_inputs_25_30_port, shift_in(29) => 
                           positive_inputs_25_29_port, shift_in(28) => 
                           positive_inputs_25_28_port, shift_in(27) => 
                           positive_inputs_25_27_port, shift_in(26) => 
                           positive_inputs_25_26_port, shift_in(25) => 
                           positive_inputs_25_25_port, shift_in(24) => 
                           positive_inputs_25_24_port, shift_in(23) => 
                           positive_inputs_25_23_port, shift_in(22) => 
                           positive_inputs_25_22_port, shift_in(21) => 
                           positive_inputs_25_21_port, shift_in(20) => 
                           positive_inputs_25_20_port, shift_in(19) => 
                           positive_inputs_25_19_port, shift_in(18) => 
                           positive_inputs_25_18_port, shift_in(17) => 
                           positive_inputs_25_17_port, shift_in(16) => 
                           positive_inputs_25_16_port, shift_in(15) => 
                           positive_inputs_25_15_port, shift_in(14) => 
                           positive_inputs_25_14_port, shift_in(13) => 
                           positive_inputs_25_13_port, shift_in(12) => 
                           positive_inputs_25_12_port, shift_in(11) => 
                           positive_inputs_25_11_port, shift_in(10) => 
                           positive_inputs_25_10_port, shift_in(9) => 
                           positive_inputs_25_9_port, shift_in(8) => 
                           positive_inputs_25_8_port, shift_in(7) => 
                           positive_inputs_25_7_port, shift_in(6) => 
                           positive_inputs_25_6_port, shift_in(5) => 
                           positive_inputs_25_5_port, shift_in(4) => 
                           positive_inputs_25_4_port, shift_in(3) => 
                           positive_inputs_25_3_port, shift_in(2) => 
                           positive_inputs_25_2_port, shift_in(1) => 
                           positive_inputs_25_1_port, shift_in(0) => n9, 
                           shift_out(63) => positive_inputs_26_63_port, 
                           shift_out(62) => positive_inputs_26_62_port, 
                           shift_out(61) => positive_inputs_26_61_port, 
                           shift_out(60) => positive_inputs_26_60_port, 
                           shift_out(59) => positive_inputs_26_59_port, 
                           shift_out(58) => positive_inputs_26_58_port, 
                           shift_out(57) => positive_inputs_26_57_port, 
                           shift_out(56) => positive_inputs_26_56_port, 
                           shift_out(55) => positive_inputs_26_55_port, 
                           shift_out(54) => positive_inputs_26_54_port, 
                           shift_out(53) => positive_inputs_26_53_port, 
                           shift_out(52) => positive_inputs_26_52_port, 
                           shift_out(51) => positive_inputs_26_51_port, 
                           shift_out(50) => positive_inputs_26_50_port, 
                           shift_out(49) => positive_inputs_26_49_port, 
                           shift_out(48) => positive_inputs_26_48_port, 
                           shift_out(47) => positive_inputs_26_47_port, 
                           shift_out(46) => positive_inputs_26_46_port, 
                           shift_out(45) => positive_inputs_26_45_port, 
                           shift_out(44) => positive_inputs_26_44_port, 
                           shift_out(43) => positive_inputs_26_43_port, 
                           shift_out(42) => positive_inputs_26_42_port, 
                           shift_out(41) => positive_inputs_26_41_port, 
                           shift_out(40) => positive_inputs_26_40_port, 
                           shift_out(39) => positive_inputs_26_39_port, 
                           shift_out(38) => positive_inputs_26_38_port, 
                           shift_out(37) => positive_inputs_26_37_port, 
                           shift_out(36) => positive_inputs_26_36_port, 
                           shift_out(35) => positive_inputs_26_35_port, 
                           shift_out(34) => positive_inputs_26_34_port, 
                           shift_out(33) => positive_inputs_26_33_port, 
                           shift_out(32) => positive_inputs_26_32_port, 
                           shift_out(31) => positive_inputs_26_31_port, 
                           shift_out(30) => positive_inputs_26_30_port, 
                           shift_out(29) => positive_inputs_26_29_port, 
                           shift_out(28) => positive_inputs_26_28_port, 
                           shift_out(27) => positive_inputs_26_27_port, 
                           shift_out(26) => positive_inputs_26_26_port, 
                           shift_out(25) => positive_inputs_26_25_port, 
                           shift_out(24) => positive_inputs_26_24_port, 
                           shift_out(23) => positive_inputs_26_23_port, 
                           shift_out(22) => positive_inputs_26_22_port, 
                           shift_out(21) => positive_inputs_26_21_port, 
                           shift_out(20) => positive_inputs_26_20_port, 
                           shift_out(19) => positive_inputs_26_19_port, 
                           shift_out(18) => positive_inputs_26_18_port, 
                           shift_out(17) => positive_inputs_26_17_port, 
                           shift_out(16) => positive_inputs_26_16_port, 
                           shift_out(15) => positive_inputs_26_15_port, 
                           shift_out(14) => positive_inputs_26_14_port, 
                           shift_out(13) => positive_inputs_26_13_port, 
                           shift_out(12) => positive_inputs_26_12_port, 
                           shift_out(11) => positive_inputs_26_11_port, 
                           shift_out(10) => positive_inputs_26_10_port, 
                           shift_out(9) => positive_inputs_26_9_port, 
                           shift_out(8) => positive_inputs_26_8_port, 
                           shift_out(7) => positive_inputs_26_7_port, 
                           shift_out(6) => positive_inputs_26_6_port, 
                           shift_out(5) => positive_inputs_26_5_port, 
                           shift_out(4) => positive_inputs_26_4_port, 
                           shift_out(3) => positive_inputs_26_3_port, 
                           shift_out(2) => positive_inputs_26_2_port, 
                           shift_out(1) => positive_inputs_26_1_port, 
                           shift_out(0) => n_1026);
   shifted_pos_27 : leftshifter_NbitShifter64_37 port map( shift_in(63) => 
                           positive_inputs_26_63_port, shift_in(62) => 
                           positive_inputs_26_62_port, shift_in(61) => 
                           positive_inputs_26_61_port, shift_in(60) => 
                           positive_inputs_26_60_port, shift_in(59) => 
                           positive_inputs_26_59_port, shift_in(58) => 
                           positive_inputs_26_58_port, shift_in(57) => 
                           positive_inputs_26_57_port, shift_in(56) => 
                           positive_inputs_26_56_port, shift_in(55) => 
                           positive_inputs_26_55_port, shift_in(54) => 
                           positive_inputs_26_54_port, shift_in(53) => 
                           positive_inputs_26_53_port, shift_in(52) => 
                           positive_inputs_26_52_port, shift_in(51) => 
                           positive_inputs_26_51_port, shift_in(50) => 
                           positive_inputs_26_50_port, shift_in(49) => 
                           positive_inputs_26_49_port, shift_in(48) => 
                           positive_inputs_26_48_port, shift_in(47) => 
                           positive_inputs_26_47_port, shift_in(46) => 
                           positive_inputs_26_46_port, shift_in(45) => 
                           positive_inputs_26_45_port, shift_in(44) => 
                           positive_inputs_26_44_port, shift_in(43) => 
                           positive_inputs_26_43_port, shift_in(42) => 
                           positive_inputs_26_42_port, shift_in(41) => 
                           positive_inputs_26_41_port, shift_in(40) => 
                           positive_inputs_26_40_port, shift_in(39) => 
                           positive_inputs_26_39_port, shift_in(38) => 
                           positive_inputs_26_38_port, shift_in(37) => 
                           positive_inputs_26_37_port, shift_in(36) => 
                           positive_inputs_26_36_port, shift_in(35) => 
                           positive_inputs_26_35_port, shift_in(34) => 
                           positive_inputs_26_34_port, shift_in(33) => 
                           positive_inputs_26_33_port, shift_in(32) => 
                           positive_inputs_26_32_port, shift_in(31) => 
                           positive_inputs_26_31_port, shift_in(30) => 
                           positive_inputs_26_30_port, shift_in(29) => 
                           positive_inputs_26_29_port, shift_in(28) => 
                           positive_inputs_26_28_port, shift_in(27) => 
                           positive_inputs_26_27_port, shift_in(26) => 
                           positive_inputs_26_26_port, shift_in(25) => 
                           positive_inputs_26_25_port, shift_in(24) => 
                           positive_inputs_26_24_port, shift_in(23) => 
                           positive_inputs_26_23_port, shift_in(22) => 
                           positive_inputs_26_22_port, shift_in(21) => 
                           positive_inputs_26_21_port, shift_in(20) => 
                           positive_inputs_26_20_port, shift_in(19) => 
                           positive_inputs_26_19_port, shift_in(18) => 
                           positive_inputs_26_18_port, shift_in(17) => 
                           positive_inputs_26_17_port, shift_in(16) => 
                           positive_inputs_26_16_port, shift_in(15) => 
                           positive_inputs_26_15_port, shift_in(14) => 
                           positive_inputs_26_14_port, shift_in(13) => 
                           positive_inputs_26_13_port, shift_in(12) => 
                           positive_inputs_26_12_port, shift_in(11) => 
                           positive_inputs_26_11_port, shift_in(10) => 
                           positive_inputs_26_10_port, shift_in(9) => 
                           positive_inputs_26_9_port, shift_in(8) => 
                           positive_inputs_26_8_port, shift_in(7) => 
                           positive_inputs_26_7_port, shift_in(6) => 
                           positive_inputs_26_6_port, shift_in(5) => 
                           positive_inputs_26_5_port, shift_in(4) => 
                           positive_inputs_26_4_port, shift_in(3) => 
                           positive_inputs_26_3_port, shift_in(2) => 
                           positive_inputs_26_2_port, shift_in(1) => 
                           positive_inputs_26_1_port, shift_in(0) => n9, 
                           shift_out(63) => positive_inputs_27_63_port, 
                           shift_out(62) => positive_inputs_27_62_port, 
                           shift_out(61) => positive_inputs_27_61_port, 
                           shift_out(60) => positive_inputs_27_60_port, 
                           shift_out(59) => positive_inputs_27_59_port, 
                           shift_out(58) => positive_inputs_27_58_port, 
                           shift_out(57) => positive_inputs_27_57_port, 
                           shift_out(56) => positive_inputs_27_56_port, 
                           shift_out(55) => positive_inputs_27_55_port, 
                           shift_out(54) => positive_inputs_27_54_port, 
                           shift_out(53) => positive_inputs_27_53_port, 
                           shift_out(52) => positive_inputs_27_52_port, 
                           shift_out(51) => positive_inputs_27_51_port, 
                           shift_out(50) => positive_inputs_27_50_port, 
                           shift_out(49) => positive_inputs_27_49_port, 
                           shift_out(48) => positive_inputs_27_48_port, 
                           shift_out(47) => positive_inputs_27_47_port, 
                           shift_out(46) => positive_inputs_27_46_port, 
                           shift_out(45) => positive_inputs_27_45_port, 
                           shift_out(44) => positive_inputs_27_44_port, 
                           shift_out(43) => positive_inputs_27_43_port, 
                           shift_out(42) => positive_inputs_27_42_port, 
                           shift_out(41) => positive_inputs_27_41_port, 
                           shift_out(40) => positive_inputs_27_40_port, 
                           shift_out(39) => positive_inputs_27_39_port, 
                           shift_out(38) => positive_inputs_27_38_port, 
                           shift_out(37) => positive_inputs_27_37_port, 
                           shift_out(36) => positive_inputs_27_36_port, 
                           shift_out(35) => positive_inputs_27_35_port, 
                           shift_out(34) => positive_inputs_27_34_port, 
                           shift_out(33) => positive_inputs_27_33_port, 
                           shift_out(32) => positive_inputs_27_32_port, 
                           shift_out(31) => positive_inputs_27_31_port, 
                           shift_out(30) => positive_inputs_27_30_port, 
                           shift_out(29) => positive_inputs_27_29_port, 
                           shift_out(28) => positive_inputs_27_28_port, 
                           shift_out(27) => positive_inputs_27_27_port, 
                           shift_out(26) => positive_inputs_27_26_port, 
                           shift_out(25) => positive_inputs_27_25_port, 
                           shift_out(24) => positive_inputs_27_24_port, 
                           shift_out(23) => positive_inputs_27_23_port, 
                           shift_out(22) => positive_inputs_27_22_port, 
                           shift_out(21) => positive_inputs_27_21_port, 
                           shift_out(20) => positive_inputs_27_20_port, 
                           shift_out(19) => positive_inputs_27_19_port, 
                           shift_out(18) => positive_inputs_27_18_port, 
                           shift_out(17) => positive_inputs_27_17_port, 
                           shift_out(16) => positive_inputs_27_16_port, 
                           shift_out(15) => positive_inputs_27_15_port, 
                           shift_out(14) => positive_inputs_27_14_port, 
                           shift_out(13) => positive_inputs_27_13_port, 
                           shift_out(12) => positive_inputs_27_12_port, 
                           shift_out(11) => positive_inputs_27_11_port, 
                           shift_out(10) => positive_inputs_27_10_port, 
                           shift_out(9) => positive_inputs_27_9_port, 
                           shift_out(8) => positive_inputs_27_8_port, 
                           shift_out(7) => positive_inputs_27_7_port, 
                           shift_out(6) => positive_inputs_27_6_port, 
                           shift_out(5) => positive_inputs_27_5_port, 
                           shift_out(4) => positive_inputs_27_4_port, 
                           shift_out(3) => positive_inputs_27_3_port, 
                           shift_out(2) => positive_inputs_27_2_port, 
                           shift_out(1) => positive_inputs_27_1_port, 
                           shift_out(0) => n_1027);
   shifted_pos_28 : leftshifter_NbitShifter64_36 port map( shift_in(63) => 
                           positive_inputs_27_63_port, shift_in(62) => 
                           positive_inputs_27_62_port, shift_in(61) => 
                           positive_inputs_27_61_port, shift_in(60) => 
                           positive_inputs_27_60_port, shift_in(59) => 
                           positive_inputs_27_59_port, shift_in(58) => 
                           positive_inputs_27_58_port, shift_in(57) => 
                           positive_inputs_27_57_port, shift_in(56) => 
                           positive_inputs_27_56_port, shift_in(55) => 
                           positive_inputs_27_55_port, shift_in(54) => 
                           positive_inputs_27_54_port, shift_in(53) => 
                           positive_inputs_27_53_port, shift_in(52) => 
                           positive_inputs_27_52_port, shift_in(51) => 
                           positive_inputs_27_51_port, shift_in(50) => 
                           positive_inputs_27_50_port, shift_in(49) => 
                           positive_inputs_27_49_port, shift_in(48) => 
                           positive_inputs_27_48_port, shift_in(47) => 
                           positive_inputs_27_47_port, shift_in(46) => 
                           positive_inputs_27_46_port, shift_in(45) => 
                           positive_inputs_27_45_port, shift_in(44) => 
                           positive_inputs_27_44_port, shift_in(43) => 
                           positive_inputs_27_43_port, shift_in(42) => 
                           positive_inputs_27_42_port, shift_in(41) => 
                           positive_inputs_27_41_port, shift_in(40) => 
                           positive_inputs_27_40_port, shift_in(39) => 
                           positive_inputs_27_39_port, shift_in(38) => 
                           positive_inputs_27_38_port, shift_in(37) => 
                           positive_inputs_27_37_port, shift_in(36) => 
                           positive_inputs_27_36_port, shift_in(35) => 
                           positive_inputs_27_35_port, shift_in(34) => 
                           positive_inputs_27_34_port, shift_in(33) => 
                           positive_inputs_27_33_port, shift_in(32) => 
                           positive_inputs_27_32_port, shift_in(31) => 
                           positive_inputs_27_31_port, shift_in(30) => 
                           positive_inputs_27_30_port, shift_in(29) => 
                           positive_inputs_27_29_port, shift_in(28) => 
                           positive_inputs_27_28_port, shift_in(27) => 
                           positive_inputs_27_27_port, shift_in(26) => 
                           positive_inputs_27_26_port, shift_in(25) => 
                           positive_inputs_27_25_port, shift_in(24) => 
                           positive_inputs_27_24_port, shift_in(23) => 
                           positive_inputs_27_23_port, shift_in(22) => 
                           positive_inputs_27_22_port, shift_in(21) => 
                           positive_inputs_27_21_port, shift_in(20) => 
                           positive_inputs_27_20_port, shift_in(19) => 
                           positive_inputs_27_19_port, shift_in(18) => 
                           positive_inputs_27_18_port, shift_in(17) => 
                           positive_inputs_27_17_port, shift_in(16) => 
                           positive_inputs_27_16_port, shift_in(15) => 
                           positive_inputs_27_15_port, shift_in(14) => 
                           positive_inputs_27_14_port, shift_in(13) => 
                           positive_inputs_27_13_port, shift_in(12) => 
                           positive_inputs_27_12_port, shift_in(11) => 
                           positive_inputs_27_11_port, shift_in(10) => 
                           positive_inputs_27_10_port, shift_in(9) => 
                           positive_inputs_27_9_port, shift_in(8) => 
                           positive_inputs_27_8_port, shift_in(7) => 
                           positive_inputs_27_7_port, shift_in(6) => 
                           positive_inputs_27_6_port, shift_in(5) => 
                           positive_inputs_27_5_port, shift_in(4) => 
                           positive_inputs_27_4_port, shift_in(3) => 
                           positive_inputs_27_3_port, shift_in(2) => 
                           positive_inputs_27_2_port, shift_in(1) => 
                           positive_inputs_27_1_port, shift_in(0) => n9, 
                           shift_out(63) => positive_inputs_28_63_port, 
                           shift_out(62) => positive_inputs_28_62_port, 
                           shift_out(61) => positive_inputs_28_61_port, 
                           shift_out(60) => positive_inputs_28_60_port, 
                           shift_out(59) => positive_inputs_28_59_port, 
                           shift_out(58) => positive_inputs_28_58_port, 
                           shift_out(57) => positive_inputs_28_57_port, 
                           shift_out(56) => positive_inputs_28_56_port, 
                           shift_out(55) => positive_inputs_28_55_port, 
                           shift_out(54) => positive_inputs_28_54_port, 
                           shift_out(53) => positive_inputs_28_53_port, 
                           shift_out(52) => positive_inputs_28_52_port, 
                           shift_out(51) => positive_inputs_28_51_port, 
                           shift_out(50) => positive_inputs_28_50_port, 
                           shift_out(49) => positive_inputs_28_49_port, 
                           shift_out(48) => positive_inputs_28_48_port, 
                           shift_out(47) => positive_inputs_28_47_port, 
                           shift_out(46) => positive_inputs_28_46_port, 
                           shift_out(45) => positive_inputs_28_45_port, 
                           shift_out(44) => positive_inputs_28_44_port, 
                           shift_out(43) => positive_inputs_28_43_port, 
                           shift_out(42) => positive_inputs_28_42_port, 
                           shift_out(41) => positive_inputs_28_41_port, 
                           shift_out(40) => positive_inputs_28_40_port, 
                           shift_out(39) => positive_inputs_28_39_port, 
                           shift_out(38) => positive_inputs_28_38_port, 
                           shift_out(37) => positive_inputs_28_37_port, 
                           shift_out(36) => positive_inputs_28_36_port, 
                           shift_out(35) => positive_inputs_28_35_port, 
                           shift_out(34) => positive_inputs_28_34_port, 
                           shift_out(33) => positive_inputs_28_33_port, 
                           shift_out(32) => positive_inputs_28_32_port, 
                           shift_out(31) => positive_inputs_28_31_port, 
                           shift_out(30) => positive_inputs_28_30_port, 
                           shift_out(29) => positive_inputs_28_29_port, 
                           shift_out(28) => positive_inputs_28_28_port, 
                           shift_out(27) => positive_inputs_28_27_port, 
                           shift_out(26) => positive_inputs_28_26_port, 
                           shift_out(25) => positive_inputs_28_25_port, 
                           shift_out(24) => positive_inputs_28_24_port, 
                           shift_out(23) => positive_inputs_28_23_port, 
                           shift_out(22) => positive_inputs_28_22_port, 
                           shift_out(21) => positive_inputs_28_21_port, 
                           shift_out(20) => positive_inputs_28_20_port, 
                           shift_out(19) => positive_inputs_28_19_port, 
                           shift_out(18) => positive_inputs_28_18_port, 
                           shift_out(17) => positive_inputs_28_17_port, 
                           shift_out(16) => positive_inputs_28_16_port, 
                           shift_out(15) => positive_inputs_28_15_port, 
                           shift_out(14) => positive_inputs_28_14_port, 
                           shift_out(13) => positive_inputs_28_13_port, 
                           shift_out(12) => positive_inputs_28_12_port, 
                           shift_out(11) => positive_inputs_28_11_port, 
                           shift_out(10) => positive_inputs_28_10_port, 
                           shift_out(9) => positive_inputs_28_9_port, 
                           shift_out(8) => positive_inputs_28_8_port, 
                           shift_out(7) => positive_inputs_28_7_port, 
                           shift_out(6) => positive_inputs_28_6_port, 
                           shift_out(5) => positive_inputs_28_5_port, 
                           shift_out(4) => positive_inputs_28_4_port, 
                           shift_out(3) => positive_inputs_28_3_port, 
                           shift_out(2) => positive_inputs_28_2_port, 
                           shift_out(1) => positive_inputs_28_1_port, 
                           shift_out(0) => n_1028);
   shifted_pos_29 : leftshifter_NbitShifter64_35 port map( shift_in(63) => 
                           positive_inputs_28_63_port, shift_in(62) => 
                           positive_inputs_28_62_port, shift_in(61) => 
                           positive_inputs_28_61_port, shift_in(60) => 
                           positive_inputs_28_60_port, shift_in(59) => 
                           positive_inputs_28_59_port, shift_in(58) => 
                           positive_inputs_28_58_port, shift_in(57) => 
                           positive_inputs_28_57_port, shift_in(56) => 
                           positive_inputs_28_56_port, shift_in(55) => 
                           positive_inputs_28_55_port, shift_in(54) => 
                           positive_inputs_28_54_port, shift_in(53) => 
                           positive_inputs_28_53_port, shift_in(52) => 
                           positive_inputs_28_52_port, shift_in(51) => 
                           positive_inputs_28_51_port, shift_in(50) => 
                           positive_inputs_28_50_port, shift_in(49) => 
                           positive_inputs_28_49_port, shift_in(48) => 
                           positive_inputs_28_48_port, shift_in(47) => 
                           positive_inputs_28_47_port, shift_in(46) => 
                           positive_inputs_28_46_port, shift_in(45) => 
                           positive_inputs_28_45_port, shift_in(44) => 
                           positive_inputs_28_44_port, shift_in(43) => 
                           positive_inputs_28_43_port, shift_in(42) => 
                           positive_inputs_28_42_port, shift_in(41) => 
                           positive_inputs_28_41_port, shift_in(40) => 
                           positive_inputs_28_40_port, shift_in(39) => 
                           positive_inputs_28_39_port, shift_in(38) => 
                           positive_inputs_28_38_port, shift_in(37) => 
                           positive_inputs_28_37_port, shift_in(36) => 
                           positive_inputs_28_36_port, shift_in(35) => 
                           positive_inputs_28_35_port, shift_in(34) => 
                           positive_inputs_28_34_port, shift_in(33) => 
                           positive_inputs_28_33_port, shift_in(32) => 
                           positive_inputs_28_32_port, shift_in(31) => 
                           positive_inputs_28_31_port, shift_in(30) => 
                           positive_inputs_28_30_port, shift_in(29) => 
                           positive_inputs_28_29_port, shift_in(28) => 
                           positive_inputs_28_28_port, shift_in(27) => 
                           positive_inputs_28_27_port, shift_in(26) => 
                           positive_inputs_28_26_port, shift_in(25) => 
                           positive_inputs_28_25_port, shift_in(24) => 
                           positive_inputs_28_24_port, shift_in(23) => 
                           positive_inputs_28_23_port, shift_in(22) => 
                           positive_inputs_28_22_port, shift_in(21) => 
                           positive_inputs_28_21_port, shift_in(20) => 
                           positive_inputs_28_20_port, shift_in(19) => 
                           positive_inputs_28_19_port, shift_in(18) => 
                           positive_inputs_28_18_port, shift_in(17) => 
                           positive_inputs_28_17_port, shift_in(16) => 
                           positive_inputs_28_16_port, shift_in(15) => 
                           positive_inputs_28_15_port, shift_in(14) => 
                           positive_inputs_28_14_port, shift_in(13) => 
                           positive_inputs_28_13_port, shift_in(12) => 
                           positive_inputs_28_12_port, shift_in(11) => 
                           positive_inputs_28_11_port, shift_in(10) => 
                           positive_inputs_28_10_port, shift_in(9) => 
                           positive_inputs_28_9_port, shift_in(8) => 
                           positive_inputs_28_8_port, shift_in(7) => 
                           positive_inputs_28_7_port, shift_in(6) => 
                           positive_inputs_28_6_port, shift_in(5) => 
                           positive_inputs_28_5_port, shift_in(4) => 
                           positive_inputs_28_4_port, shift_in(3) => 
                           positive_inputs_28_3_port, shift_in(2) => 
                           positive_inputs_28_2_port, shift_in(1) => 
                           positive_inputs_28_1_port, shift_in(0) => n9, 
                           shift_out(63) => positive_inputs_29_63_port, 
                           shift_out(62) => positive_inputs_29_62_port, 
                           shift_out(61) => positive_inputs_29_61_port, 
                           shift_out(60) => positive_inputs_29_60_port, 
                           shift_out(59) => positive_inputs_29_59_port, 
                           shift_out(58) => positive_inputs_29_58_port, 
                           shift_out(57) => positive_inputs_29_57_port, 
                           shift_out(56) => positive_inputs_29_56_port, 
                           shift_out(55) => positive_inputs_29_55_port, 
                           shift_out(54) => positive_inputs_29_54_port, 
                           shift_out(53) => positive_inputs_29_53_port, 
                           shift_out(52) => positive_inputs_29_52_port, 
                           shift_out(51) => positive_inputs_29_51_port, 
                           shift_out(50) => positive_inputs_29_50_port, 
                           shift_out(49) => positive_inputs_29_49_port, 
                           shift_out(48) => positive_inputs_29_48_port, 
                           shift_out(47) => positive_inputs_29_47_port, 
                           shift_out(46) => positive_inputs_29_46_port, 
                           shift_out(45) => positive_inputs_29_45_port, 
                           shift_out(44) => positive_inputs_29_44_port, 
                           shift_out(43) => positive_inputs_29_43_port, 
                           shift_out(42) => positive_inputs_29_42_port, 
                           shift_out(41) => positive_inputs_29_41_port, 
                           shift_out(40) => positive_inputs_29_40_port, 
                           shift_out(39) => positive_inputs_29_39_port, 
                           shift_out(38) => positive_inputs_29_38_port, 
                           shift_out(37) => positive_inputs_29_37_port, 
                           shift_out(36) => positive_inputs_29_36_port, 
                           shift_out(35) => positive_inputs_29_35_port, 
                           shift_out(34) => positive_inputs_29_34_port, 
                           shift_out(33) => positive_inputs_29_33_port, 
                           shift_out(32) => positive_inputs_29_32_port, 
                           shift_out(31) => positive_inputs_29_31_port, 
                           shift_out(30) => positive_inputs_29_30_port, 
                           shift_out(29) => positive_inputs_29_29_port, 
                           shift_out(28) => positive_inputs_29_28_port, 
                           shift_out(27) => positive_inputs_29_27_port, 
                           shift_out(26) => positive_inputs_29_26_port, 
                           shift_out(25) => positive_inputs_29_25_port, 
                           shift_out(24) => positive_inputs_29_24_port, 
                           shift_out(23) => positive_inputs_29_23_port, 
                           shift_out(22) => positive_inputs_29_22_port, 
                           shift_out(21) => positive_inputs_29_21_port, 
                           shift_out(20) => positive_inputs_29_20_port, 
                           shift_out(19) => positive_inputs_29_19_port, 
                           shift_out(18) => positive_inputs_29_18_port, 
                           shift_out(17) => positive_inputs_29_17_port, 
                           shift_out(16) => positive_inputs_29_16_port, 
                           shift_out(15) => positive_inputs_29_15_port, 
                           shift_out(14) => positive_inputs_29_14_port, 
                           shift_out(13) => positive_inputs_29_13_port, 
                           shift_out(12) => positive_inputs_29_12_port, 
                           shift_out(11) => positive_inputs_29_11_port, 
                           shift_out(10) => positive_inputs_29_10_port, 
                           shift_out(9) => positive_inputs_29_9_port, 
                           shift_out(8) => positive_inputs_29_8_port, 
                           shift_out(7) => positive_inputs_29_7_port, 
                           shift_out(6) => positive_inputs_29_6_port, 
                           shift_out(5) => positive_inputs_29_5_port, 
                           shift_out(4) => positive_inputs_29_4_port, 
                           shift_out(3) => positive_inputs_29_3_port, 
                           shift_out(2) => positive_inputs_29_2_port, 
                           shift_out(1) => positive_inputs_29_1_port, 
                           shift_out(0) => n_1029);
   shifted_pos_30 : leftshifter_NbitShifter64_34 port map( shift_in(63) => 
                           positive_inputs_29_63_port, shift_in(62) => 
                           positive_inputs_29_62_port, shift_in(61) => 
                           positive_inputs_29_61_port, shift_in(60) => 
                           positive_inputs_29_60_port, shift_in(59) => 
                           positive_inputs_29_59_port, shift_in(58) => 
                           positive_inputs_29_58_port, shift_in(57) => 
                           positive_inputs_29_57_port, shift_in(56) => 
                           positive_inputs_29_56_port, shift_in(55) => 
                           positive_inputs_29_55_port, shift_in(54) => 
                           positive_inputs_29_54_port, shift_in(53) => 
                           positive_inputs_29_53_port, shift_in(52) => 
                           positive_inputs_29_52_port, shift_in(51) => 
                           positive_inputs_29_51_port, shift_in(50) => 
                           positive_inputs_29_50_port, shift_in(49) => 
                           positive_inputs_29_49_port, shift_in(48) => 
                           positive_inputs_29_48_port, shift_in(47) => 
                           positive_inputs_29_47_port, shift_in(46) => 
                           positive_inputs_29_46_port, shift_in(45) => 
                           positive_inputs_29_45_port, shift_in(44) => 
                           positive_inputs_29_44_port, shift_in(43) => 
                           positive_inputs_29_43_port, shift_in(42) => 
                           positive_inputs_29_42_port, shift_in(41) => 
                           positive_inputs_29_41_port, shift_in(40) => 
                           positive_inputs_29_40_port, shift_in(39) => 
                           positive_inputs_29_39_port, shift_in(38) => 
                           positive_inputs_29_38_port, shift_in(37) => 
                           positive_inputs_29_37_port, shift_in(36) => 
                           positive_inputs_29_36_port, shift_in(35) => 
                           positive_inputs_29_35_port, shift_in(34) => 
                           positive_inputs_29_34_port, shift_in(33) => 
                           positive_inputs_29_33_port, shift_in(32) => 
                           positive_inputs_29_32_port, shift_in(31) => 
                           positive_inputs_29_31_port, shift_in(30) => 
                           positive_inputs_29_30_port, shift_in(29) => 
                           positive_inputs_29_29_port, shift_in(28) => 
                           positive_inputs_29_28_port, shift_in(27) => 
                           positive_inputs_29_27_port, shift_in(26) => 
                           positive_inputs_29_26_port, shift_in(25) => 
                           positive_inputs_29_25_port, shift_in(24) => 
                           positive_inputs_29_24_port, shift_in(23) => 
                           positive_inputs_29_23_port, shift_in(22) => 
                           positive_inputs_29_22_port, shift_in(21) => 
                           positive_inputs_29_21_port, shift_in(20) => 
                           positive_inputs_29_20_port, shift_in(19) => 
                           positive_inputs_29_19_port, shift_in(18) => 
                           positive_inputs_29_18_port, shift_in(17) => 
                           positive_inputs_29_17_port, shift_in(16) => 
                           positive_inputs_29_16_port, shift_in(15) => 
                           positive_inputs_29_15_port, shift_in(14) => 
                           positive_inputs_29_14_port, shift_in(13) => 
                           positive_inputs_29_13_port, shift_in(12) => 
                           positive_inputs_29_12_port, shift_in(11) => 
                           positive_inputs_29_11_port, shift_in(10) => 
                           positive_inputs_29_10_port, shift_in(9) => 
                           positive_inputs_29_9_port, shift_in(8) => 
                           positive_inputs_29_8_port, shift_in(7) => 
                           positive_inputs_29_7_port, shift_in(6) => 
                           positive_inputs_29_6_port, shift_in(5) => 
                           positive_inputs_29_5_port, shift_in(4) => 
                           positive_inputs_29_4_port, shift_in(3) => 
                           positive_inputs_29_3_port, shift_in(2) => 
                           positive_inputs_29_2_port, shift_in(1) => 
                           positive_inputs_29_1_port, shift_in(0) => n9, 
                           shift_out(63) => positive_inputs_30_63_port, 
                           shift_out(62) => positive_inputs_30_62_port, 
                           shift_out(61) => positive_inputs_30_61_port, 
                           shift_out(60) => positive_inputs_30_60_port, 
                           shift_out(59) => positive_inputs_30_59_port, 
                           shift_out(58) => positive_inputs_30_58_port, 
                           shift_out(57) => positive_inputs_30_57_port, 
                           shift_out(56) => positive_inputs_30_56_port, 
                           shift_out(55) => positive_inputs_30_55_port, 
                           shift_out(54) => positive_inputs_30_54_port, 
                           shift_out(53) => positive_inputs_30_53_port, 
                           shift_out(52) => positive_inputs_30_52_port, 
                           shift_out(51) => positive_inputs_30_51_port, 
                           shift_out(50) => positive_inputs_30_50_port, 
                           shift_out(49) => positive_inputs_30_49_port, 
                           shift_out(48) => positive_inputs_30_48_port, 
                           shift_out(47) => positive_inputs_30_47_port, 
                           shift_out(46) => positive_inputs_30_46_port, 
                           shift_out(45) => positive_inputs_30_45_port, 
                           shift_out(44) => positive_inputs_30_44_port, 
                           shift_out(43) => positive_inputs_30_43_port, 
                           shift_out(42) => positive_inputs_30_42_port, 
                           shift_out(41) => positive_inputs_30_41_port, 
                           shift_out(40) => positive_inputs_30_40_port, 
                           shift_out(39) => positive_inputs_30_39_port, 
                           shift_out(38) => positive_inputs_30_38_port, 
                           shift_out(37) => positive_inputs_30_37_port, 
                           shift_out(36) => positive_inputs_30_36_port, 
                           shift_out(35) => positive_inputs_30_35_port, 
                           shift_out(34) => positive_inputs_30_34_port, 
                           shift_out(33) => positive_inputs_30_33_port, 
                           shift_out(32) => positive_inputs_30_32_port, 
                           shift_out(31) => positive_inputs_30_31_port, 
                           shift_out(30) => positive_inputs_30_30_port, 
                           shift_out(29) => positive_inputs_30_29_port, 
                           shift_out(28) => positive_inputs_30_28_port, 
                           shift_out(27) => positive_inputs_30_27_port, 
                           shift_out(26) => positive_inputs_30_26_port, 
                           shift_out(25) => positive_inputs_30_25_port, 
                           shift_out(24) => positive_inputs_30_24_port, 
                           shift_out(23) => positive_inputs_30_23_port, 
                           shift_out(22) => positive_inputs_30_22_port, 
                           shift_out(21) => positive_inputs_30_21_port, 
                           shift_out(20) => positive_inputs_30_20_port, 
                           shift_out(19) => positive_inputs_30_19_port, 
                           shift_out(18) => positive_inputs_30_18_port, 
                           shift_out(17) => positive_inputs_30_17_port, 
                           shift_out(16) => positive_inputs_30_16_port, 
                           shift_out(15) => positive_inputs_30_15_port, 
                           shift_out(14) => positive_inputs_30_14_port, 
                           shift_out(13) => positive_inputs_30_13_port, 
                           shift_out(12) => positive_inputs_30_12_port, 
                           shift_out(11) => positive_inputs_30_11_port, 
                           shift_out(10) => positive_inputs_30_10_port, 
                           shift_out(9) => positive_inputs_30_9_port, 
                           shift_out(8) => positive_inputs_30_8_port, 
                           shift_out(7) => positive_inputs_30_7_port, 
                           shift_out(6) => positive_inputs_30_6_port, 
                           shift_out(5) => positive_inputs_30_5_port, 
                           shift_out(4) => positive_inputs_30_4_port, 
                           shift_out(3) => positive_inputs_30_3_port, 
                           shift_out(2) => positive_inputs_30_2_port, 
                           shift_out(1) => positive_inputs_30_1_port, 
                           shift_out(0) => n_1030);
   shifted_pos_31 : leftshifter_NbitShifter64_33 port map( shift_in(63) => 
                           positive_inputs_30_63_port, shift_in(62) => 
                           positive_inputs_30_62_port, shift_in(61) => 
                           positive_inputs_30_61_port, shift_in(60) => 
                           positive_inputs_30_60_port, shift_in(59) => 
                           positive_inputs_30_59_port, shift_in(58) => 
                           positive_inputs_30_58_port, shift_in(57) => 
                           positive_inputs_30_57_port, shift_in(56) => 
                           positive_inputs_30_56_port, shift_in(55) => 
                           positive_inputs_30_55_port, shift_in(54) => 
                           positive_inputs_30_54_port, shift_in(53) => 
                           positive_inputs_30_53_port, shift_in(52) => 
                           positive_inputs_30_52_port, shift_in(51) => 
                           positive_inputs_30_51_port, shift_in(50) => 
                           positive_inputs_30_50_port, shift_in(49) => 
                           positive_inputs_30_49_port, shift_in(48) => 
                           positive_inputs_30_48_port, shift_in(47) => 
                           positive_inputs_30_47_port, shift_in(46) => 
                           positive_inputs_30_46_port, shift_in(45) => 
                           positive_inputs_30_45_port, shift_in(44) => 
                           positive_inputs_30_44_port, shift_in(43) => 
                           positive_inputs_30_43_port, shift_in(42) => 
                           positive_inputs_30_42_port, shift_in(41) => 
                           positive_inputs_30_41_port, shift_in(40) => 
                           positive_inputs_30_40_port, shift_in(39) => 
                           positive_inputs_30_39_port, shift_in(38) => 
                           positive_inputs_30_38_port, shift_in(37) => 
                           positive_inputs_30_37_port, shift_in(36) => 
                           positive_inputs_30_36_port, shift_in(35) => 
                           positive_inputs_30_35_port, shift_in(34) => 
                           positive_inputs_30_34_port, shift_in(33) => 
                           positive_inputs_30_33_port, shift_in(32) => 
                           positive_inputs_30_32_port, shift_in(31) => 
                           positive_inputs_30_31_port, shift_in(30) => 
                           positive_inputs_30_30_port, shift_in(29) => 
                           positive_inputs_30_29_port, shift_in(28) => 
                           positive_inputs_30_28_port, shift_in(27) => 
                           positive_inputs_30_27_port, shift_in(26) => 
                           positive_inputs_30_26_port, shift_in(25) => 
                           positive_inputs_30_25_port, shift_in(24) => 
                           positive_inputs_30_24_port, shift_in(23) => 
                           positive_inputs_30_23_port, shift_in(22) => 
                           positive_inputs_30_22_port, shift_in(21) => 
                           positive_inputs_30_21_port, shift_in(20) => 
                           positive_inputs_30_20_port, shift_in(19) => 
                           positive_inputs_30_19_port, shift_in(18) => 
                           positive_inputs_30_18_port, shift_in(17) => 
                           positive_inputs_30_17_port, shift_in(16) => 
                           positive_inputs_30_16_port, shift_in(15) => 
                           positive_inputs_30_15_port, shift_in(14) => 
                           positive_inputs_30_14_port, shift_in(13) => 
                           positive_inputs_30_13_port, shift_in(12) => 
                           positive_inputs_30_12_port, shift_in(11) => 
                           positive_inputs_30_11_port, shift_in(10) => 
                           positive_inputs_30_10_port, shift_in(9) => 
                           positive_inputs_30_9_port, shift_in(8) => 
                           positive_inputs_30_8_port, shift_in(7) => 
                           positive_inputs_30_7_port, shift_in(6) => 
                           positive_inputs_30_6_port, shift_in(5) => 
                           positive_inputs_30_5_port, shift_in(4) => 
                           positive_inputs_30_4_port, shift_in(3) => 
                           positive_inputs_30_3_port, shift_in(2) => 
                           positive_inputs_30_2_port, shift_in(1) => 
                           positive_inputs_30_1_port, shift_in(0) => n9, 
                           shift_out(63) => positive_inputs_31_63_port, 
                           shift_out(62) => positive_inputs_31_62_port, 
                           shift_out(61) => positive_inputs_31_61_port, 
                           shift_out(60) => positive_inputs_31_60_port, 
                           shift_out(59) => positive_inputs_31_59_port, 
                           shift_out(58) => positive_inputs_31_58_port, 
                           shift_out(57) => positive_inputs_31_57_port, 
                           shift_out(56) => positive_inputs_31_56_port, 
                           shift_out(55) => positive_inputs_31_55_port, 
                           shift_out(54) => positive_inputs_31_54_port, 
                           shift_out(53) => positive_inputs_31_53_port, 
                           shift_out(52) => positive_inputs_31_52_port, 
                           shift_out(51) => positive_inputs_31_51_port, 
                           shift_out(50) => positive_inputs_31_50_port, 
                           shift_out(49) => positive_inputs_31_49_port, 
                           shift_out(48) => positive_inputs_31_48_port, 
                           shift_out(47) => positive_inputs_31_47_port, 
                           shift_out(46) => positive_inputs_31_46_port, 
                           shift_out(45) => positive_inputs_31_45_port, 
                           shift_out(44) => positive_inputs_31_44_port, 
                           shift_out(43) => positive_inputs_31_43_port, 
                           shift_out(42) => positive_inputs_31_42_port, 
                           shift_out(41) => positive_inputs_31_41_port, 
                           shift_out(40) => positive_inputs_31_40_port, 
                           shift_out(39) => positive_inputs_31_39_port, 
                           shift_out(38) => positive_inputs_31_38_port, 
                           shift_out(37) => positive_inputs_31_37_port, 
                           shift_out(36) => positive_inputs_31_36_port, 
                           shift_out(35) => positive_inputs_31_35_port, 
                           shift_out(34) => positive_inputs_31_34_port, 
                           shift_out(33) => positive_inputs_31_33_port, 
                           shift_out(32) => positive_inputs_31_32_port, 
                           shift_out(31) => positive_inputs_31_31_port, 
                           shift_out(30) => positive_inputs_31_30_port, 
                           shift_out(29) => positive_inputs_31_29_port, 
                           shift_out(28) => positive_inputs_31_28_port, 
                           shift_out(27) => positive_inputs_31_27_port, 
                           shift_out(26) => positive_inputs_31_26_port, 
                           shift_out(25) => positive_inputs_31_25_port, 
                           shift_out(24) => positive_inputs_31_24_port, 
                           shift_out(23) => positive_inputs_31_23_port, 
                           shift_out(22) => positive_inputs_31_22_port, 
                           shift_out(21) => positive_inputs_31_21_port, 
                           shift_out(20) => positive_inputs_31_20_port, 
                           shift_out(19) => positive_inputs_31_19_port, 
                           shift_out(18) => positive_inputs_31_18_port, 
                           shift_out(17) => positive_inputs_31_17_port, 
                           shift_out(16) => positive_inputs_31_16_port, 
                           shift_out(15) => positive_inputs_31_15_port, 
                           shift_out(14) => positive_inputs_31_14_port, 
                           shift_out(13) => positive_inputs_31_13_port, 
                           shift_out(12) => positive_inputs_31_12_port, 
                           shift_out(11) => positive_inputs_31_11_port, 
                           shift_out(10) => positive_inputs_31_10_port, 
                           shift_out(9) => positive_inputs_31_9_port, 
                           shift_out(8) => positive_inputs_31_8_port, 
                           shift_out(7) => positive_inputs_31_7_port, 
                           shift_out(6) => positive_inputs_31_6_port, 
                           shift_out(5) => positive_inputs_31_5_port, 
                           shift_out(4) => positive_inputs_31_4_port, 
                           shift_out(3) => positive_inputs_31_3_port, 
                           shift_out(2) => positive_inputs_31_2_port, 
                           shift_out(1) => positive_inputs_31_1_port, 
                           shift_out(0) => n_1031);
   shifted_pos_32 : leftshifter_NbitShifter64_32 port map( shift_in(63) => 
                           positive_inputs_31_63_port, shift_in(62) => 
                           positive_inputs_31_62_port, shift_in(61) => 
                           positive_inputs_31_61_port, shift_in(60) => 
                           positive_inputs_31_60_port, shift_in(59) => 
                           positive_inputs_31_59_port, shift_in(58) => 
                           positive_inputs_31_58_port, shift_in(57) => 
                           positive_inputs_31_57_port, shift_in(56) => 
                           positive_inputs_31_56_port, shift_in(55) => 
                           positive_inputs_31_55_port, shift_in(54) => 
                           positive_inputs_31_54_port, shift_in(53) => 
                           positive_inputs_31_53_port, shift_in(52) => 
                           positive_inputs_31_52_port, shift_in(51) => 
                           positive_inputs_31_51_port, shift_in(50) => 
                           positive_inputs_31_50_port, shift_in(49) => 
                           positive_inputs_31_49_port, shift_in(48) => 
                           positive_inputs_31_48_port, shift_in(47) => 
                           positive_inputs_31_47_port, shift_in(46) => 
                           positive_inputs_31_46_port, shift_in(45) => 
                           positive_inputs_31_45_port, shift_in(44) => 
                           positive_inputs_31_44_port, shift_in(43) => 
                           positive_inputs_31_43_port, shift_in(42) => 
                           positive_inputs_31_42_port, shift_in(41) => 
                           positive_inputs_31_41_port, shift_in(40) => 
                           positive_inputs_31_40_port, shift_in(39) => 
                           positive_inputs_31_39_port, shift_in(38) => 
                           positive_inputs_31_38_port, shift_in(37) => 
                           positive_inputs_31_37_port, shift_in(36) => 
                           positive_inputs_31_36_port, shift_in(35) => 
                           positive_inputs_31_35_port, shift_in(34) => 
                           positive_inputs_31_34_port, shift_in(33) => 
                           positive_inputs_31_33_port, shift_in(32) => 
                           positive_inputs_31_32_port, shift_in(31) => 
                           positive_inputs_31_31_port, shift_in(30) => 
                           positive_inputs_31_30_port, shift_in(29) => 
                           positive_inputs_31_29_port, shift_in(28) => 
                           positive_inputs_31_28_port, shift_in(27) => 
                           positive_inputs_31_27_port, shift_in(26) => 
                           positive_inputs_31_26_port, shift_in(25) => 
                           positive_inputs_31_25_port, shift_in(24) => 
                           positive_inputs_31_24_port, shift_in(23) => 
                           positive_inputs_31_23_port, shift_in(22) => 
                           positive_inputs_31_22_port, shift_in(21) => 
                           positive_inputs_31_21_port, shift_in(20) => 
                           positive_inputs_31_20_port, shift_in(19) => 
                           positive_inputs_31_19_port, shift_in(18) => 
                           positive_inputs_31_18_port, shift_in(17) => 
                           positive_inputs_31_17_port, shift_in(16) => 
                           positive_inputs_31_16_port, shift_in(15) => 
                           positive_inputs_31_15_port, shift_in(14) => 
                           positive_inputs_31_14_port, shift_in(13) => 
                           positive_inputs_31_13_port, shift_in(12) => 
                           positive_inputs_31_12_port, shift_in(11) => 
                           positive_inputs_31_11_port, shift_in(10) => 
                           positive_inputs_31_10_port, shift_in(9) => 
                           positive_inputs_31_9_port, shift_in(8) => 
                           positive_inputs_31_8_port, shift_in(7) => 
                           positive_inputs_31_7_port, shift_in(6) => 
                           positive_inputs_31_6_port, shift_in(5) => 
                           positive_inputs_31_5_port, shift_in(4) => 
                           positive_inputs_31_4_port, shift_in(3) => 
                           positive_inputs_31_3_port, shift_in(2) => 
                           positive_inputs_31_2_port, shift_in(1) => 
                           positive_inputs_31_1_port, shift_in(0) => n9, 
                           shift_out(63) => n_1032, shift_out(62) => n_1033, 
                           shift_out(61) => n_1034, shift_out(60) => n_1035, 
                           shift_out(59) => n_1036, shift_out(58) => n_1037, 
                           shift_out(57) => n_1038, shift_out(56) => n_1039, 
                           shift_out(55) => n_1040, shift_out(54) => n_1041, 
                           shift_out(53) => n_1042, shift_out(52) => n_1043, 
                           shift_out(51) => n_1044, shift_out(50) => n_1045, 
                           shift_out(49) => n_1046, shift_out(48) => n_1047, 
                           shift_out(47) => n_1048, shift_out(46) => n_1049, 
                           shift_out(45) => n_1050, shift_out(44) => n_1051, 
                           shift_out(43) => n_1052, shift_out(42) => n_1053, 
                           shift_out(41) => n_1054, shift_out(40) => n_1055, 
                           shift_out(39) => n_1056, shift_out(38) => n_1057, 
                           shift_out(37) => n_1058, shift_out(36) => n_1059, 
                           shift_out(35) => n_1060, shift_out(34) => n_1061, 
                           shift_out(33) => n_1062, shift_out(32) => n_1063, 
                           shift_out(31) => n_1064, shift_out(30) => n_1065, 
                           shift_out(29) => n_1066, shift_out(28) => n_1067, 
                           shift_out(27) => n_1068, shift_out(26) => n_1069, 
                           shift_out(25) => n_1070, shift_out(24) => n_1071, 
                           shift_out(23) => n_1072, shift_out(22) => n_1073, 
                           shift_out(21) => n_1074, shift_out(20) => n_1075, 
                           shift_out(19) => n_1076, shift_out(18) => n_1077, 
                           shift_out(17) => n_1078, shift_out(16) => n_1079, 
                           shift_out(15) => n_1080, shift_out(14) => n_1081, 
                           shift_out(13) => n_1082, shift_out(12) => n_1083, 
                           shift_out(11) => n_1084, shift_out(10) => n_1085, 
                           shift_out(9) => n_1086, shift_out(8) => n_1087, 
                           shift_out(7) => n_1088, shift_out(6) => n_1089, 
                           shift_out(5) => n_1090, shift_out(4) => n_1091, 
                           shift_out(3) => n_1092, shift_out(2) => n_1093, 
                           shift_out(1) => n_1094, shift_out(0) => n_1095);
   shifted_neg_1 : leftshifter_NbitShifter64_31 port map( shift_in(63) => 
                           negative_inputs_0_63_port, shift_in(62) => 
                           negative_inputs_0_62_port, shift_in(61) => 
                           negative_inputs_0_61_port, shift_in(60) => 
                           negative_inputs_0_60_port, shift_in(59) => 
                           negative_inputs_0_59_port, shift_in(58) => 
                           negative_inputs_0_58_port, shift_in(57) => 
                           negative_inputs_0_57_port, shift_in(56) => 
                           negative_inputs_0_56_port, shift_in(55) => 
                           negative_inputs_0_55_port, shift_in(54) => 
                           negative_inputs_0_54_port, shift_in(53) => 
                           negative_inputs_0_53_port, shift_in(52) => 
                           negative_inputs_0_52_port, shift_in(51) => 
                           negative_inputs_0_51_port, shift_in(50) => 
                           negative_inputs_0_50_port, shift_in(49) => 
                           negative_inputs_0_49_port, shift_in(48) => 
                           negative_inputs_0_48_port, shift_in(47) => n14, 
                           shift_in(46) => n27, shift_in(45) => n31, 
                           shift_in(44) => negative_inputs_0_44_port, 
                           shift_in(43) => negative_inputs_0_43_port, 
                           shift_in(42) => negative_inputs_0_42_port, 
                           shift_in(41) => negative_inputs_0_41_port, 
                           shift_in(40) => negative_inputs_0_40_port, 
                           shift_in(39) => n151, shift_in(38) => 
                           negative_inputs_0_38_port, shift_in(37) => 
                           negative_inputs_0_37_port, shift_in(36) => 
                           negative_inputs_0_36_port, shift_in(35) => 
                           negative_inputs_0_35_port, shift_in(34) => 
                           negative_inputs_0_34_port, shift_in(33) => 
                           negative_inputs_0_33_port, shift_in(32) => n15, 
                           shift_in(31) => n23, shift_in(30) => n22, 
                           shift_in(29) => n24, shift_in(28) => n28, 
                           shift_in(27) => n25, shift_in(26) => 
                           negative_inputs_0_26_port, shift_in(25) => n36, 
                           shift_in(24) => n10, shift_in(23) => n39, 
                           shift_in(22) => n33, shift_in(21) => 
                           negative_inputs_0_21_port, shift_in(20) => n32, 
                           shift_in(19) => n29, shift_in(18) => 
                           negative_inputs_0_18_port, shift_in(17) => n16, 
                           shift_in(16) => n19, shift_in(15) => n40, 
                           shift_in(14) => n47, shift_in(13) => n38, 
                           shift_in(12) => negative_inputs_0_12_port, 
                           shift_in(11) => n43, shift_in(10) => n46, 
                           shift_in(9) => n45, shift_in(8) => n44, shift_in(7) 
                           => negative_inputs_0_7_port, shift_in(6) => 
                           negative_inputs_0_6_port, shift_in(5) => n48, 
                           shift_in(4) => n37, shift_in(3) => n71, shift_in(2) 
                           => negative_inputs_0_2_port, shift_in(1) => 
                           negative_inputs_0_1_port, shift_in(0) => 
                           negative_inputs_0_0_port, shift_out(63) => 
                           negative_inputs_1_63_port, shift_out(62) => 
                           negative_inputs_1_62_port, shift_out(61) => 
                           negative_inputs_1_61_port, shift_out(60) => 
                           negative_inputs_1_60_port, shift_out(59) => 
                           negative_inputs_1_59_port, shift_out(58) => 
                           negative_inputs_1_58_port, shift_out(57) => 
                           negative_inputs_1_57_port, shift_out(56) => 
                           negative_inputs_1_56_port, shift_out(55) => 
                           negative_inputs_1_55_port, shift_out(54) => 
                           negative_inputs_1_54_port, shift_out(53) => 
                           negative_inputs_1_53_port, shift_out(52) => 
                           negative_inputs_1_52_port, shift_out(51) => 
                           negative_inputs_1_51_port, shift_out(50) => 
                           negative_inputs_1_50_port, shift_out(49) => 
                           negative_inputs_1_49_port, shift_out(48) => 
                           negative_inputs_1_48_port, shift_out(47) => 
                           negative_inputs_1_47_port, shift_out(46) => 
                           negative_inputs_1_46_port, shift_out(45) => 
                           negative_inputs_1_45_port, shift_out(44) => 
                           negative_inputs_1_44_port, shift_out(43) => 
                           negative_inputs_1_43_port, shift_out(42) => 
                           negative_inputs_1_42_port, shift_out(41) => 
                           negative_inputs_1_41_port, shift_out(40) => 
                           negative_inputs_1_40_port, shift_out(39) => 
                           negative_inputs_1_39_port, shift_out(38) => 
                           negative_inputs_1_38_port, shift_out(37) => 
                           negative_inputs_1_37_port, shift_out(36) => 
                           negative_inputs_1_36_port, shift_out(35) => 
                           negative_inputs_1_35_port, shift_out(34) => 
                           negative_inputs_1_34_port, shift_out(33) => 
                           negative_inputs_1_33_port, shift_out(32) => 
                           negative_inputs_1_32_port, shift_out(31) => 
                           negative_inputs_1_31_port, shift_out(30) => 
                           negative_inputs_1_30_port, shift_out(29) => 
                           negative_inputs_1_29_port, shift_out(28) => 
                           negative_inputs_1_28_port, shift_out(27) => 
                           negative_inputs_1_27_port, shift_out(26) => 
                           negative_inputs_1_26_port, shift_out(25) => 
                           negative_inputs_1_25_port, shift_out(24) => 
                           negative_inputs_1_24_port, shift_out(23) => 
                           negative_inputs_1_23_port, shift_out(22) => 
                           negative_inputs_1_22_port, shift_out(21) => 
                           negative_inputs_1_21_port, shift_out(20) => 
                           negative_inputs_1_20_port, shift_out(19) => 
                           negative_inputs_1_19_port, shift_out(18) => 
                           negative_inputs_1_18_port, shift_out(17) => 
                           negative_inputs_1_17_port, shift_out(16) => 
                           negative_inputs_1_16_port, shift_out(15) => 
                           negative_inputs_1_15_port, shift_out(14) => 
                           negative_inputs_1_14_port, shift_out(13) => 
                           negative_inputs_1_13_port, shift_out(12) => 
                           negative_inputs_1_12_port, shift_out(11) => 
                           negative_inputs_1_11_port, shift_out(10) => 
                           negative_inputs_1_10_port, shift_out(9) => 
                           negative_inputs_1_9_port, shift_out(8) => 
                           negative_inputs_1_8_port, shift_out(7) => 
                           negative_inputs_1_7_port, shift_out(6) => 
                           negative_inputs_1_6_port, shift_out(5) => 
                           negative_inputs_1_5_port, shift_out(4) => 
                           negative_inputs_1_4_port, shift_out(3) => 
                           negative_inputs_1_3_port, shift_out(2) => 
                           negative_inputs_1_2_port, shift_out(1) => 
                           negative_inputs_1_1_port, shift_out(0) => n_1096);
   shifted_neg_2 : leftshifter_NbitShifter64_30 port map( shift_in(63) => 
                           negative_inputs_1_63_port, shift_in(62) => 
                           negative_inputs_1_62_port, shift_in(61) => 
                           negative_inputs_1_61_port, shift_in(60) => 
                           negative_inputs_1_60_port, shift_in(59) => 
                           negative_inputs_1_59_port, shift_in(58) => 
                           negative_inputs_1_58_port, shift_in(57) => 
                           negative_inputs_1_57_port, shift_in(56) => 
                           negative_inputs_1_56_port, shift_in(55) => 
                           negative_inputs_1_55_port, shift_in(54) => 
                           negative_inputs_1_54_port, shift_in(53) => 
                           negative_inputs_1_53_port, shift_in(52) => 
                           negative_inputs_1_52_port, shift_in(51) => 
                           negative_inputs_1_51_port, shift_in(50) => 
                           negative_inputs_1_50_port, shift_in(49) => 
                           negative_inputs_1_49_port, shift_in(48) => 
                           negative_inputs_1_48_port, shift_in(47) => 
                           negative_inputs_1_47_port, shift_in(46) => 
                           negative_inputs_1_46_port, shift_in(45) => 
                           negative_inputs_1_45_port, shift_in(44) => 
                           negative_inputs_1_44_port, shift_in(43) => n42, 
                           shift_in(42) => negative_inputs_1_42_port, 
                           shift_in(41) => negative_inputs_1_41_port, 
                           shift_in(40) => negative_inputs_1_40_port, 
                           shift_in(39) => n149, shift_in(38) => 
                           negative_inputs_1_38_port, shift_in(37) => 
                           negative_inputs_1_37_port, shift_in(36) => 
                           negative_inputs_1_36_port, shift_in(35) => 
                           negative_inputs_1_35_port, shift_in(34) => 
                           negative_inputs_1_34_port, shift_in(33) => 
                           negative_inputs_1_33_port, shift_in(32) => 
                           negative_inputs_1_32_port, shift_in(31) => 
                           negative_inputs_1_31_port, shift_in(30) => 
                           negative_inputs_1_30_port, shift_in(29) => 
                           negative_inputs_1_29_port, shift_in(28) => 
                           negative_inputs_1_28_port, shift_in(27) => 
                           negative_inputs_1_27_port, shift_in(26) => 
                           negative_inputs_1_26_port, shift_in(25) => 
                           negative_inputs_1_25_port, shift_in(24) => 
                           negative_inputs_1_24_port, shift_in(23) => 
                           negative_inputs_1_23_port, shift_in(22) => 
                           negative_inputs_1_22_port, shift_in(21) => 
                           negative_inputs_1_21_port, shift_in(20) => 
                           negative_inputs_1_20_port, shift_in(19) => 
                           negative_inputs_1_19_port, shift_in(18) => 
                           negative_inputs_1_18_port, shift_in(17) => 
                           negative_inputs_1_17_port, shift_in(16) => 
                           negative_inputs_1_16_port, shift_in(15) => 
                           negative_inputs_1_15_port, shift_in(14) => 
                           negative_inputs_1_14_port, shift_in(13) => n13, 
                           shift_in(12) => negative_inputs_1_12_port, 
                           shift_in(11) => n17, shift_in(10) => n18, 
                           shift_in(9) => negative_inputs_1_9_port, shift_in(8)
                           => n20, shift_in(7) => n35, shift_in(6) => n34, 
                           shift_in(5) => n21, shift_in(4) => 
                           negative_inputs_1_4_port, shift_in(3) => n12, 
                           shift_in(2) => negative_inputs_1_2_port, shift_in(1)
                           => negative_inputs_1_1_port, shift_in(0) => n9, 
                           shift_out(63) => negative_inputs_2_63_port, 
                           shift_out(62) => negative_inputs_2_62_port, 
                           shift_out(61) => negative_inputs_2_61_port, 
                           shift_out(60) => negative_inputs_2_60_port, 
                           shift_out(59) => negative_inputs_2_59_port, 
                           shift_out(58) => negative_inputs_2_58_port, 
                           shift_out(57) => negative_inputs_2_57_port, 
                           shift_out(56) => negative_inputs_2_56_port, 
                           shift_out(55) => negative_inputs_2_55_port, 
                           shift_out(54) => negative_inputs_2_54_port, 
                           shift_out(53) => negative_inputs_2_53_port, 
                           shift_out(52) => negative_inputs_2_52_port, 
                           shift_out(51) => negative_inputs_2_51_port, 
                           shift_out(50) => negative_inputs_2_50_port, 
                           shift_out(49) => negative_inputs_2_49_port, 
                           shift_out(48) => negative_inputs_2_48_port, 
                           shift_out(47) => negative_inputs_2_47_port, 
                           shift_out(46) => negative_inputs_2_46_port, 
                           shift_out(45) => negative_inputs_2_45_port, 
                           shift_out(44) => negative_inputs_2_44_port, 
                           shift_out(43) => negative_inputs_2_43_port, 
                           shift_out(42) => negative_inputs_2_42_port, 
                           shift_out(41) => negative_inputs_2_41_port, 
                           shift_out(40) => negative_inputs_2_40_port, 
                           shift_out(39) => negative_inputs_2_39_port, 
                           shift_out(38) => negative_inputs_2_38_port, 
                           shift_out(37) => negative_inputs_2_37_port, 
                           shift_out(36) => negative_inputs_2_36_port, 
                           shift_out(35) => negative_inputs_2_35_port, 
                           shift_out(34) => negative_inputs_2_34_port, 
                           shift_out(33) => negative_inputs_2_33_port, 
                           shift_out(32) => negative_inputs_2_32_port, 
                           shift_out(31) => negative_inputs_2_31_port, 
                           shift_out(30) => negative_inputs_2_30_port, 
                           shift_out(29) => negative_inputs_2_29_port, 
                           shift_out(28) => negative_inputs_2_28_port, 
                           shift_out(27) => negative_inputs_2_27_port, 
                           shift_out(26) => negative_inputs_2_26_port, 
                           shift_out(25) => negative_inputs_2_25_port, 
                           shift_out(24) => negative_inputs_2_24_port, 
                           shift_out(23) => negative_inputs_2_23_port, 
                           shift_out(22) => negative_inputs_2_22_port, 
                           shift_out(21) => negative_inputs_2_21_port, 
                           shift_out(20) => negative_inputs_2_20_port, 
                           shift_out(19) => negative_inputs_2_19_port, 
                           shift_out(18) => negative_inputs_2_18_port, 
                           shift_out(17) => negative_inputs_2_17_port, 
                           shift_out(16) => negative_inputs_2_16_port, 
                           shift_out(15) => negative_inputs_2_15_port, 
                           shift_out(14) => negative_inputs_2_14_port, 
                           shift_out(13) => negative_inputs_2_13_port, 
                           shift_out(12) => negative_inputs_2_12_port, 
                           shift_out(11) => negative_inputs_2_11_port, 
                           shift_out(10) => negative_inputs_2_10_port, 
                           shift_out(9) => negative_inputs_2_9_port, 
                           shift_out(8) => negative_inputs_2_8_port, 
                           shift_out(7) => negative_inputs_2_7_port, 
                           shift_out(6) => negative_inputs_2_6_port, 
                           shift_out(5) => negative_inputs_2_5_port, 
                           shift_out(4) => negative_inputs_2_4_port, 
                           shift_out(3) => negative_inputs_2_3_port, 
                           shift_out(2) => negative_inputs_2_2_port, 
                           shift_out(1) => negative_inputs_2_1_port, 
                           shift_out(0) => n_1097);
   shifted_neg_3 : leftshifter_NbitShifter64_29 port map( shift_in(63) => 
                           negative_inputs_2_63_port, shift_in(62) => 
                           negative_inputs_2_62_port, shift_in(61) => 
                           negative_inputs_2_61_port, shift_in(60) => 
                           negative_inputs_2_60_port, shift_in(59) => 
                           negative_inputs_2_59_port, shift_in(58) => 
                           negative_inputs_2_58_port, shift_in(57) => 
                           negative_inputs_2_57_port, shift_in(56) => 
                           negative_inputs_2_56_port, shift_in(55) => 
                           negative_inputs_2_55_port, shift_in(54) => 
                           negative_inputs_2_54_port, shift_in(53) => 
                           negative_inputs_2_53_port, shift_in(52) => 
                           negative_inputs_2_52_port, shift_in(51) => 
                           negative_inputs_2_51_port, shift_in(50) => 
                           negative_inputs_2_50_port, shift_in(49) => 
                           negative_inputs_2_49_port, shift_in(48) => 
                           negative_inputs_2_48_port, shift_in(47) => 
                           negative_inputs_2_47_port, shift_in(46) => 
                           negative_inputs_2_46_port, shift_in(45) => 
                           negative_inputs_2_45_port, shift_in(44) => 
                           negative_inputs_2_44_port, shift_in(43) => 
                           negative_inputs_2_43_port, shift_in(42) => 
                           negative_inputs_2_42_port, shift_in(41) => 
                           negative_inputs_2_41_port, shift_in(40) => 
                           negative_inputs_2_40_port, shift_in(39) => n147, 
                           shift_in(38) => negative_inputs_2_38_port, 
                           shift_in(37) => negative_inputs_2_37_port, 
                           shift_in(36) => negative_inputs_2_36_port, 
                           shift_in(35) => negative_inputs_2_35_port, 
                           shift_in(34) => negative_inputs_2_34_port, 
                           shift_in(33) => negative_inputs_2_33_port, 
                           shift_in(32) => negative_inputs_2_32_port, 
                           shift_in(31) => negative_inputs_2_31_port, 
                           shift_in(30) => negative_inputs_2_30_port, 
                           shift_in(29) => negative_inputs_2_29_port, 
                           shift_in(28) => negative_inputs_2_28_port, 
                           shift_in(27) => negative_inputs_2_27_port, 
                           shift_in(26) => negative_inputs_2_26_port, 
                           shift_in(25) => negative_inputs_2_25_port, 
                           shift_in(24) => negative_inputs_2_24_port, 
                           shift_in(23) => negative_inputs_2_23_port, 
                           shift_in(22) => negative_inputs_2_22_port, 
                           shift_in(21) => negative_inputs_2_21_port, 
                           shift_in(20) => negative_inputs_2_20_port, 
                           shift_in(19) => negative_inputs_2_19_port, 
                           shift_in(18) => negative_inputs_2_18_port, 
                           shift_in(17) => negative_inputs_2_17_port, 
                           shift_in(16) => negative_inputs_2_16_port, 
                           shift_in(15) => negative_inputs_2_15_port, 
                           shift_in(14) => negative_inputs_2_14_port, 
                           shift_in(13) => negative_inputs_2_13_port, 
                           shift_in(12) => negative_inputs_2_12_port, 
                           shift_in(11) => negative_inputs_2_11_port, 
                           shift_in(10) => negative_inputs_2_10_port, 
                           shift_in(9) => negative_inputs_2_9_port, shift_in(8)
                           => negative_inputs_2_8_port, shift_in(7) => 
                           negative_inputs_2_7_port, shift_in(6) => 
                           negative_inputs_2_6_port, shift_in(5) => 
                           negative_inputs_2_5_port, shift_in(4) => 
                           negative_inputs_2_4_port, shift_in(3) => 
                           negative_inputs_2_3_port, shift_in(2) => 
                           negative_inputs_2_2_port, shift_in(1) => 
                           negative_inputs_2_1_port, shift_in(0) => n9, 
                           shift_out(63) => negative_inputs_3_63_port, 
                           shift_out(62) => negative_inputs_3_62_port, 
                           shift_out(61) => negative_inputs_3_61_port, 
                           shift_out(60) => negative_inputs_3_60_port, 
                           shift_out(59) => negative_inputs_3_59_port, 
                           shift_out(58) => negative_inputs_3_58_port, 
                           shift_out(57) => negative_inputs_3_57_port, 
                           shift_out(56) => negative_inputs_3_56_port, 
                           shift_out(55) => negative_inputs_3_55_port, 
                           shift_out(54) => negative_inputs_3_54_port, 
                           shift_out(53) => negative_inputs_3_53_port, 
                           shift_out(52) => negative_inputs_3_52_port, 
                           shift_out(51) => negative_inputs_3_51_port, 
                           shift_out(50) => negative_inputs_3_50_port, 
                           shift_out(49) => negative_inputs_3_49_port, 
                           shift_out(48) => negative_inputs_3_48_port, 
                           shift_out(47) => negative_inputs_3_47_port, 
                           shift_out(46) => negative_inputs_3_46_port, 
                           shift_out(45) => negative_inputs_3_45_port, 
                           shift_out(44) => negative_inputs_3_44_port, 
                           shift_out(43) => negative_inputs_3_43_port, 
                           shift_out(42) => negative_inputs_3_42_port, 
                           shift_out(41) => negative_inputs_3_41_port, 
                           shift_out(40) => negative_inputs_3_40_port, 
                           shift_out(39) => negative_inputs_3_39_port, 
                           shift_out(38) => negative_inputs_3_38_port, 
                           shift_out(37) => negative_inputs_3_37_port, 
                           shift_out(36) => negative_inputs_3_36_port, 
                           shift_out(35) => negative_inputs_3_35_port, 
                           shift_out(34) => negative_inputs_3_34_port, 
                           shift_out(33) => negative_inputs_3_33_port, 
                           shift_out(32) => negative_inputs_3_32_port, 
                           shift_out(31) => negative_inputs_3_31_port, 
                           shift_out(30) => negative_inputs_3_30_port, 
                           shift_out(29) => negative_inputs_3_29_port, 
                           shift_out(28) => negative_inputs_3_28_port, 
                           shift_out(27) => negative_inputs_3_27_port, 
                           shift_out(26) => negative_inputs_3_26_port, 
                           shift_out(25) => negative_inputs_3_25_port, 
                           shift_out(24) => negative_inputs_3_24_port, 
                           shift_out(23) => negative_inputs_3_23_port, 
                           shift_out(22) => negative_inputs_3_22_port, 
                           shift_out(21) => negative_inputs_3_21_port, 
                           shift_out(20) => negative_inputs_3_20_port, 
                           shift_out(19) => negative_inputs_3_19_port, 
                           shift_out(18) => negative_inputs_3_18_port, 
                           shift_out(17) => negative_inputs_3_17_port, 
                           shift_out(16) => negative_inputs_3_16_port, 
                           shift_out(15) => negative_inputs_3_15_port, 
                           shift_out(14) => negative_inputs_3_14_port, 
                           shift_out(13) => negative_inputs_3_13_port, 
                           shift_out(12) => negative_inputs_3_12_port, 
                           shift_out(11) => negative_inputs_3_11_port, 
                           shift_out(10) => negative_inputs_3_10_port, 
                           shift_out(9) => negative_inputs_3_9_port, 
                           shift_out(8) => negative_inputs_3_8_port, 
                           shift_out(7) => negative_inputs_3_7_port, 
                           shift_out(6) => negative_inputs_3_6_port, 
                           shift_out(5) => negative_inputs_3_5_port, 
                           shift_out(4) => negative_inputs_3_4_port, 
                           shift_out(3) => negative_inputs_3_3_port, 
                           shift_out(2) => negative_inputs_3_2_port, 
                           shift_out(1) => negative_inputs_3_1_port, 
                           shift_out(0) => n_1098);
   shifted_neg_4 : leftshifter_NbitShifter64_28 port map( shift_in(63) => 
                           negative_inputs_3_63_port, shift_in(62) => 
                           negative_inputs_3_62_port, shift_in(61) => 
                           negative_inputs_3_61_port, shift_in(60) => 
                           negative_inputs_3_60_port, shift_in(59) => 
                           negative_inputs_3_59_port, shift_in(58) => 
                           negative_inputs_3_58_port, shift_in(57) => 
                           negative_inputs_3_57_port, shift_in(56) => 
                           negative_inputs_3_56_port, shift_in(55) => 
                           negative_inputs_3_55_port, shift_in(54) => 
                           negative_inputs_3_54_port, shift_in(53) => 
                           negative_inputs_3_53_port, shift_in(52) => 
                           negative_inputs_3_52_port, shift_in(51) => 
                           negative_inputs_3_51_port, shift_in(50) => 
                           negative_inputs_3_50_port, shift_in(49) => 
                           negative_inputs_3_49_port, shift_in(48) => 
                           negative_inputs_3_48_port, shift_in(47) => 
                           negative_inputs_3_47_port, shift_in(46) => 
                           negative_inputs_3_46_port, shift_in(45) => 
                           negative_inputs_3_45_port, shift_in(44) => 
                           negative_inputs_3_44_port, shift_in(43) => 
                           negative_inputs_3_43_port, shift_in(42) => 
                           negative_inputs_3_42_port, shift_in(41) => 
                           negative_inputs_3_41_port, shift_in(40) => 
                           negative_inputs_3_40_port, shift_in(39) => n145, 
                           shift_in(38) => negative_inputs_3_38_port, 
                           shift_in(37) => negative_inputs_3_37_port, 
                           shift_in(36) => negative_inputs_3_36_port, 
                           shift_in(35) => negative_inputs_3_35_port, 
                           shift_in(34) => negative_inputs_3_34_port, 
                           shift_in(33) => negative_inputs_3_33_port, 
                           shift_in(32) => negative_inputs_3_32_port, 
                           shift_in(31) => negative_inputs_3_31_port, 
                           shift_in(30) => negative_inputs_3_30_port, 
                           shift_in(29) => negative_inputs_3_29_port, 
                           shift_in(28) => negative_inputs_3_28_port, 
                           shift_in(27) => negative_inputs_3_27_port, 
                           shift_in(26) => negative_inputs_3_26_port, 
                           shift_in(25) => negative_inputs_3_25_port, 
                           shift_in(24) => negative_inputs_3_24_port, 
                           shift_in(23) => negative_inputs_3_23_port, 
                           shift_in(22) => negative_inputs_3_22_port, 
                           shift_in(21) => negative_inputs_3_21_port, 
                           shift_in(20) => negative_inputs_3_20_port, 
                           shift_in(19) => negative_inputs_3_19_port, 
                           shift_in(18) => negative_inputs_3_18_port, 
                           shift_in(17) => negative_inputs_3_17_port, 
                           shift_in(16) => negative_inputs_3_16_port, 
                           shift_in(15) => negative_inputs_3_15_port, 
                           shift_in(14) => negative_inputs_3_14_port, 
                           shift_in(13) => negative_inputs_3_13_port, 
                           shift_in(12) => negative_inputs_3_12_port, 
                           shift_in(11) => negative_inputs_3_11_port, 
                           shift_in(10) => negative_inputs_3_10_port, 
                           shift_in(9) => negative_inputs_3_9_port, shift_in(8)
                           => negative_inputs_3_8_port, shift_in(7) => 
                           negative_inputs_3_7_port, shift_in(6) => 
                           negative_inputs_3_6_port, shift_in(5) => 
                           negative_inputs_3_5_port, shift_in(4) => 
                           negative_inputs_3_4_port, shift_in(3) => 
                           negative_inputs_3_3_port, shift_in(2) => 
                           negative_inputs_3_2_port, shift_in(1) => 
                           negative_inputs_3_1_port, shift_in(0) => n9, 
                           shift_out(63) => negative_inputs_4_63_port, 
                           shift_out(62) => negative_inputs_4_62_port, 
                           shift_out(61) => negative_inputs_4_61_port, 
                           shift_out(60) => negative_inputs_4_60_port, 
                           shift_out(59) => negative_inputs_4_59_port, 
                           shift_out(58) => negative_inputs_4_58_port, 
                           shift_out(57) => negative_inputs_4_57_port, 
                           shift_out(56) => negative_inputs_4_56_port, 
                           shift_out(55) => negative_inputs_4_55_port, 
                           shift_out(54) => negative_inputs_4_54_port, 
                           shift_out(53) => negative_inputs_4_53_port, 
                           shift_out(52) => negative_inputs_4_52_port, 
                           shift_out(51) => negative_inputs_4_51_port, 
                           shift_out(50) => negative_inputs_4_50_port, 
                           shift_out(49) => negative_inputs_4_49_port, 
                           shift_out(48) => negative_inputs_4_48_port, 
                           shift_out(47) => negative_inputs_4_47_port, 
                           shift_out(46) => negative_inputs_4_46_port, 
                           shift_out(45) => negative_inputs_4_45_port, 
                           shift_out(44) => negative_inputs_4_44_port, 
                           shift_out(43) => negative_inputs_4_43_port, 
                           shift_out(42) => negative_inputs_4_42_port, 
                           shift_out(41) => negative_inputs_4_41_port, 
                           shift_out(40) => negative_inputs_4_40_port, 
                           shift_out(39) => negative_inputs_4_39_port, 
                           shift_out(38) => negative_inputs_4_38_port, 
                           shift_out(37) => negative_inputs_4_37_port, 
                           shift_out(36) => negative_inputs_4_36_port, 
                           shift_out(35) => negative_inputs_4_35_port, 
                           shift_out(34) => negative_inputs_4_34_port, 
                           shift_out(33) => negative_inputs_4_33_port, 
                           shift_out(32) => negative_inputs_4_32_port, 
                           shift_out(31) => negative_inputs_4_31_port, 
                           shift_out(30) => negative_inputs_4_30_port, 
                           shift_out(29) => negative_inputs_4_29_port, 
                           shift_out(28) => negative_inputs_4_28_port, 
                           shift_out(27) => negative_inputs_4_27_port, 
                           shift_out(26) => negative_inputs_4_26_port, 
                           shift_out(25) => negative_inputs_4_25_port, 
                           shift_out(24) => negative_inputs_4_24_port, 
                           shift_out(23) => negative_inputs_4_23_port, 
                           shift_out(22) => negative_inputs_4_22_port, 
                           shift_out(21) => negative_inputs_4_21_port, 
                           shift_out(20) => negative_inputs_4_20_port, 
                           shift_out(19) => negative_inputs_4_19_port, 
                           shift_out(18) => negative_inputs_4_18_port, 
                           shift_out(17) => negative_inputs_4_17_port, 
                           shift_out(16) => negative_inputs_4_16_port, 
                           shift_out(15) => negative_inputs_4_15_port, 
                           shift_out(14) => negative_inputs_4_14_port, 
                           shift_out(13) => negative_inputs_4_13_port, 
                           shift_out(12) => negative_inputs_4_12_port, 
                           shift_out(11) => negative_inputs_4_11_port, 
                           shift_out(10) => negative_inputs_4_10_port, 
                           shift_out(9) => negative_inputs_4_9_port, 
                           shift_out(8) => negative_inputs_4_8_port, 
                           shift_out(7) => negative_inputs_4_7_port, 
                           shift_out(6) => negative_inputs_4_6_port, 
                           shift_out(5) => negative_inputs_4_5_port, 
                           shift_out(4) => negative_inputs_4_4_port, 
                           shift_out(3) => negative_inputs_4_3_port, 
                           shift_out(2) => negative_inputs_4_2_port, 
                           shift_out(1) => negative_inputs_4_1_port, 
                           shift_out(0) => n_1099);
   shifted_neg_5 : leftshifter_NbitShifter64_27 port map( shift_in(63) => 
                           negative_inputs_4_63_port, shift_in(62) => 
                           negative_inputs_4_62_port, shift_in(61) => 
                           negative_inputs_4_61_port, shift_in(60) => 
                           negative_inputs_4_60_port, shift_in(59) => 
                           negative_inputs_4_59_port, shift_in(58) => 
                           negative_inputs_4_58_port, shift_in(57) => 
                           negative_inputs_4_57_port, shift_in(56) => 
                           negative_inputs_4_56_port, shift_in(55) => 
                           negative_inputs_4_55_port, shift_in(54) => 
                           negative_inputs_4_54_port, shift_in(53) => 
                           negative_inputs_4_53_port, shift_in(52) => 
                           negative_inputs_4_52_port, shift_in(51) => 
                           negative_inputs_4_51_port, shift_in(50) => 
                           negative_inputs_4_50_port, shift_in(49) => 
                           negative_inputs_4_49_port, shift_in(48) => 
                           negative_inputs_4_48_port, shift_in(47) => 
                           negative_inputs_4_47_port, shift_in(46) => 
                           negative_inputs_4_46_port, shift_in(45) => 
                           negative_inputs_4_45_port, shift_in(44) => 
                           negative_inputs_4_44_port, shift_in(43) => 
                           negative_inputs_4_43_port, shift_in(42) => 
                           negative_inputs_4_42_port, shift_in(41) => 
                           negative_inputs_4_41_port, shift_in(40) => 
                           negative_inputs_4_40_port, shift_in(39) => n143, 
                           shift_in(38) => negative_inputs_4_38_port, 
                           shift_in(37) => negative_inputs_4_37_port, 
                           shift_in(36) => negative_inputs_4_36_port, 
                           shift_in(35) => negative_inputs_4_35_port, 
                           shift_in(34) => negative_inputs_4_34_port, 
                           shift_in(33) => negative_inputs_4_33_port, 
                           shift_in(32) => negative_inputs_4_32_port, 
                           shift_in(31) => negative_inputs_4_31_port, 
                           shift_in(30) => negative_inputs_4_30_port, 
                           shift_in(29) => negative_inputs_4_29_port, 
                           shift_in(28) => negative_inputs_4_28_port, 
                           shift_in(27) => negative_inputs_4_27_port, 
                           shift_in(26) => negative_inputs_4_26_port, 
                           shift_in(25) => negative_inputs_4_25_port, 
                           shift_in(24) => negative_inputs_4_24_port, 
                           shift_in(23) => negative_inputs_4_23_port, 
                           shift_in(22) => negative_inputs_4_22_port, 
                           shift_in(21) => negative_inputs_4_21_port, 
                           shift_in(20) => negative_inputs_4_20_port, 
                           shift_in(19) => negative_inputs_4_19_port, 
                           shift_in(18) => negative_inputs_4_18_port, 
                           shift_in(17) => negative_inputs_4_17_port, 
                           shift_in(16) => negative_inputs_4_16_port, 
                           shift_in(15) => negative_inputs_4_15_port, 
                           shift_in(14) => negative_inputs_4_14_port, 
                           shift_in(13) => negative_inputs_4_13_port, 
                           shift_in(12) => negative_inputs_4_12_port, 
                           shift_in(11) => negative_inputs_4_11_port, 
                           shift_in(10) => negative_inputs_4_10_port, 
                           shift_in(9) => negative_inputs_4_9_port, shift_in(8)
                           => negative_inputs_4_8_port, shift_in(7) => 
                           negative_inputs_4_7_port, shift_in(6) => 
                           negative_inputs_4_6_port, shift_in(5) => 
                           negative_inputs_4_5_port, shift_in(4) => 
                           negative_inputs_4_4_port, shift_in(3) => 
                           negative_inputs_4_3_port, shift_in(2) => 
                           negative_inputs_4_2_port, shift_in(1) => 
                           negative_inputs_4_1_port, shift_in(0) => n9, 
                           shift_out(63) => negative_inputs_5_63_port, 
                           shift_out(62) => negative_inputs_5_62_port, 
                           shift_out(61) => negative_inputs_5_61_port, 
                           shift_out(60) => negative_inputs_5_60_port, 
                           shift_out(59) => negative_inputs_5_59_port, 
                           shift_out(58) => negative_inputs_5_58_port, 
                           shift_out(57) => negative_inputs_5_57_port, 
                           shift_out(56) => negative_inputs_5_56_port, 
                           shift_out(55) => negative_inputs_5_55_port, 
                           shift_out(54) => negative_inputs_5_54_port, 
                           shift_out(53) => negative_inputs_5_53_port, 
                           shift_out(52) => negative_inputs_5_52_port, 
                           shift_out(51) => negative_inputs_5_51_port, 
                           shift_out(50) => negative_inputs_5_50_port, 
                           shift_out(49) => negative_inputs_5_49_port, 
                           shift_out(48) => negative_inputs_5_48_port, 
                           shift_out(47) => negative_inputs_5_47_port, 
                           shift_out(46) => negative_inputs_5_46_port, 
                           shift_out(45) => negative_inputs_5_45_port, 
                           shift_out(44) => negative_inputs_5_44_port, 
                           shift_out(43) => negative_inputs_5_43_port, 
                           shift_out(42) => negative_inputs_5_42_port, 
                           shift_out(41) => negative_inputs_5_41_port, 
                           shift_out(40) => negative_inputs_5_40_port, 
                           shift_out(39) => negative_inputs_5_39_port, 
                           shift_out(38) => negative_inputs_5_38_port, 
                           shift_out(37) => negative_inputs_5_37_port, 
                           shift_out(36) => negative_inputs_5_36_port, 
                           shift_out(35) => negative_inputs_5_35_port, 
                           shift_out(34) => negative_inputs_5_34_port, 
                           shift_out(33) => negative_inputs_5_33_port, 
                           shift_out(32) => negative_inputs_5_32_port, 
                           shift_out(31) => negative_inputs_5_31_port, 
                           shift_out(30) => negative_inputs_5_30_port, 
                           shift_out(29) => negative_inputs_5_29_port, 
                           shift_out(28) => negative_inputs_5_28_port, 
                           shift_out(27) => negative_inputs_5_27_port, 
                           shift_out(26) => negative_inputs_5_26_port, 
                           shift_out(25) => negative_inputs_5_25_port, 
                           shift_out(24) => negative_inputs_5_24_port, 
                           shift_out(23) => negative_inputs_5_23_port, 
                           shift_out(22) => negative_inputs_5_22_port, 
                           shift_out(21) => negative_inputs_5_21_port, 
                           shift_out(20) => negative_inputs_5_20_port, 
                           shift_out(19) => negative_inputs_5_19_port, 
                           shift_out(18) => negative_inputs_5_18_port, 
                           shift_out(17) => negative_inputs_5_17_port, 
                           shift_out(16) => negative_inputs_5_16_port, 
                           shift_out(15) => negative_inputs_5_15_port, 
                           shift_out(14) => negative_inputs_5_14_port, 
                           shift_out(13) => negative_inputs_5_13_port, 
                           shift_out(12) => negative_inputs_5_12_port, 
                           shift_out(11) => negative_inputs_5_11_port, 
                           shift_out(10) => negative_inputs_5_10_port, 
                           shift_out(9) => negative_inputs_5_9_port, 
                           shift_out(8) => negative_inputs_5_8_port, 
                           shift_out(7) => negative_inputs_5_7_port, 
                           shift_out(6) => negative_inputs_5_6_port, 
                           shift_out(5) => negative_inputs_5_5_port, 
                           shift_out(4) => negative_inputs_5_4_port, 
                           shift_out(3) => negative_inputs_5_3_port, 
                           shift_out(2) => negative_inputs_5_2_port, 
                           shift_out(1) => negative_inputs_5_1_port, 
                           shift_out(0) => n_1100);
   shifted_neg_6 : leftshifter_NbitShifter64_26 port map( shift_in(63) => 
                           negative_inputs_5_63_port, shift_in(62) => 
                           negative_inputs_5_62_port, shift_in(61) => 
                           negative_inputs_5_61_port, shift_in(60) => 
                           negative_inputs_5_60_port, shift_in(59) => 
                           negative_inputs_5_59_port, shift_in(58) => 
                           negative_inputs_5_58_port, shift_in(57) => 
                           negative_inputs_5_57_port, shift_in(56) => 
                           negative_inputs_5_56_port, shift_in(55) => 
                           negative_inputs_5_55_port, shift_in(54) => 
                           negative_inputs_5_54_port, shift_in(53) => 
                           negative_inputs_5_53_port, shift_in(52) => 
                           negative_inputs_5_52_port, shift_in(51) => 
                           negative_inputs_5_51_port, shift_in(50) => 
                           negative_inputs_5_50_port, shift_in(49) => 
                           negative_inputs_5_49_port, shift_in(48) => 
                           negative_inputs_5_48_port, shift_in(47) => 
                           negative_inputs_5_47_port, shift_in(46) => 
                           negative_inputs_5_46_port, shift_in(45) => 
                           negative_inputs_5_45_port, shift_in(44) => 
                           negative_inputs_5_44_port, shift_in(43) => 
                           negative_inputs_5_43_port, shift_in(42) => 
                           negative_inputs_5_42_port, shift_in(41) => 
                           negative_inputs_5_41_port, shift_in(40) => 
                           negative_inputs_5_40_port, shift_in(39) => n141, 
                           shift_in(38) => negative_inputs_5_38_port, 
                           shift_in(37) => negative_inputs_5_37_port, 
                           shift_in(36) => negative_inputs_5_36_port, 
                           shift_in(35) => negative_inputs_5_35_port, 
                           shift_in(34) => negative_inputs_5_34_port, 
                           shift_in(33) => negative_inputs_5_33_port, 
                           shift_in(32) => negative_inputs_5_32_port, 
                           shift_in(31) => negative_inputs_5_31_port, 
                           shift_in(30) => negative_inputs_5_30_port, 
                           shift_in(29) => negative_inputs_5_29_port, 
                           shift_in(28) => negative_inputs_5_28_port, 
                           shift_in(27) => negative_inputs_5_27_port, 
                           shift_in(26) => negative_inputs_5_26_port, 
                           shift_in(25) => negative_inputs_5_25_port, 
                           shift_in(24) => negative_inputs_5_24_port, 
                           shift_in(23) => negative_inputs_5_23_port, 
                           shift_in(22) => negative_inputs_5_22_port, 
                           shift_in(21) => negative_inputs_5_21_port, 
                           shift_in(20) => negative_inputs_5_20_port, 
                           shift_in(19) => negative_inputs_5_19_port, 
                           shift_in(18) => negative_inputs_5_18_port, 
                           shift_in(17) => negative_inputs_5_17_port, 
                           shift_in(16) => negative_inputs_5_16_port, 
                           shift_in(15) => negative_inputs_5_15_port, 
                           shift_in(14) => negative_inputs_5_14_port, 
                           shift_in(13) => negative_inputs_5_13_port, 
                           shift_in(12) => negative_inputs_5_12_port, 
                           shift_in(11) => negative_inputs_5_11_port, 
                           shift_in(10) => negative_inputs_5_10_port, 
                           shift_in(9) => negative_inputs_5_9_port, shift_in(8)
                           => negative_inputs_5_8_port, shift_in(7) => 
                           negative_inputs_5_7_port, shift_in(6) => 
                           negative_inputs_5_6_port, shift_in(5) => 
                           negative_inputs_5_5_port, shift_in(4) => 
                           negative_inputs_5_4_port, shift_in(3) => 
                           negative_inputs_5_3_port, shift_in(2) => 
                           negative_inputs_5_2_port, shift_in(1) => 
                           negative_inputs_5_1_port, shift_in(0) => n9, 
                           shift_out(63) => negative_inputs_6_63_port, 
                           shift_out(62) => negative_inputs_6_62_port, 
                           shift_out(61) => negative_inputs_6_61_port, 
                           shift_out(60) => negative_inputs_6_60_port, 
                           shift_out(59) => negative_inputs_6_59_port, 
                           shift_out(58) => negative_inputs_6_58_port, 
                           shift_out(57) => negative_inputs_6_57_port, 
                           shift_out(56) => negative_inputs_6_56_port, 
                           shift_out(55) => negative_inputs_6_55_port, 
                           shift_out(54) => negative_inputs_6_54_port, 
                           shift_out(53) => negative_inputs_6_53_port, 
                           shift_out(52) => negative_inputs_6_52_port, 
                           shift_out(51) => negative_inputs_6_51_port, 
                           shift_out(50) => negative_inputs_6_50_port, 
                           shift_out(49) => negative_inputs_6_49_port, 
                           shift_out(48) => negative_inputs_6_48_port, 
                           shift_out(47) => negative_inputs_6_47_port, 
                           shift_out(46) => negative_inputs_6_46_port, 
                           shift_out(45) => negative_inputs_6_45_port, 
                           shift_out(44) => negative_inputs_6_44_port, 
                           shift_out(43) => negative_inputs_6_43_port, 
                           shift_out(42) => negative_inputs_6_42_port, 
                           shift_out(41) => negative_inputs_6_41_port, 
                           shift_out(40) => negative_inputs_6_40_port, 
                           shift_out(39) => negative_inputs_6_39_port, 
                           shift_out(38) => negative_inputs_6_38_port, 
                           shift_out(37) => negative_inputs_6_37_port, 
                           shift_out(36) => negative_inputs_6_36_port, 
                           shift_out(35) => negative_inputs_6_35_port, 
                           shift_out(34) => negative_inputs_6_34_port, 
                           shift_out(33) => negative_inputs_6_33_port, 
                           shift_out(32) => negative_inputs_6_32_port, 
                           shift_out(31) => negative_inputs_6_31_port, 
                           shift_out(30) => negative_inputs_6_30_port, 
                           shift_out(29) => negative_inputs_6_29_port, 
                           shift_out(28) => negative_inputs_6_28_port, 
                           shift_out(27) => negative_inputs_6_27_port, 
                           shift_out(26) => negative_inputs_6_26_port, 
                           shift_out(25) => negative_inputs_6_25_port, 
                           shift_out(24) => negative_inputs_6_24_port, 
                           shift_out(23) => negative_inputs_6_23_port, 
                           shift_out(22) => negative_inputs_6_22_port, 
                           shift_out(21) => negative_inputs_6_21_port, 
                           shift_out(20) => negative_inputs_6_20_port, 
                           shift_out(19) => negative_inputs_6_19_port, 
                           shift_out(18) => negative_inputs_6_18_port, 
                           shift_out(17) => negative_inputs_6_17_port, 
                           shift_out(16) => negative_inputs_6_16_port, 
                           shift_out(15) => negative_inputs_6_15_port, 
                           shift_out(14) => negative_inputs_6_14_port, 
                           shift_out(13) => negative_inputs_6_13_port, 
                           shift_out(12) => negative_inputs_6_12_port, 
                           shift_out(11) => negative_inputs_6_11_port, 
                           shift_out(10) => negative_inputs_6_10_port, 
                           shift_out(9) => negative_inputs_6_9_port, 
                           shift_out(8) => negative_inputs_6_8_port, 
                           shift_out(7) => negative_inputs_6_7_port, 
                           shift_out(6) => negative_inputs_6_6_port, 
                           shift_out(5) => negative_inputs_6_5_port, 
                           shift_out(4) => negative_inputs_6_4_port, 
                           shift_out(3) => negative_inputs_6_3_port, 
                           shift_out(2) => negative_inputs_6_2_port, 
                           shift_out(1) => negative_inputs_6_1_port, 
                           shift_out(0) => n_1101);
   shifted_neg_7 : leftshifter_NbitShifter64_25 port map( shift_in(63) => 
                           negative_inputs_6_63_port, shift_in(62) => 
                           negative_inputs_6_62_port, shift_in(61) => 
                           negative_inputs_6_61_port, shift_in(60) => 
                           negative_inputs_6_60_port, shift_in(59) => 
                           negative_inputs_6_59_port, shift_in(58) => 
                           negative_inputs_6_58_port, shift_in(57) => 
                           negative_inputs_6_57_port, shift_in(56) => 
                           negative_inputs_6_56_port, shift_in(55) => 
                           negative_inputs_6_55_port, shift_in(54) => 
                           negative_inputs_6_54_port, shift_in(53) => 
                           negative_inputs_6_53_port, shift_in(52) => 
                           negative_inputs_6_52_port, shift_in(51) => 
                           negative_inputs_6_51_port, shift_in(50) => 
                           negative_inputs_6_50_port, shift_in(49) => 
                           negative_inputs_6_49_port, shift_in(48) => 
                           negative_inputs_6_48_port, shift_in(47) => 
                           negative_inputs_6_47_port, shift_in(46) => 
                           negative_inputs_6_46_port, shift_in(45) => 
                           negative_inputs_6_45_port, shift_in(44) => 
                           negative_inputs_6_44_port, shift_in(43) => 
                           negative_inputs_6_43_port, shift_in(42) => 
                           negative_inputs_6_42_port, shift_in(41) => 
                           negative_inputs_6_41_port, shift_in(40) => 
                           negative_inputs_6_40_port, shift_in(39) => n139, 
                           shift_in(38) => negative_inputs_6_38_port, 
                           shift_in(37) => negative_inputs_6_37_port, 
                           shift_in(36) => negative_inputs_6_36_port, 
                           shift_in(35) => negative_inputs_6_35_port, 
                           shift_in(34) => negative_inputs_6_34_port, 
                           shift_in(33) => negative_inputs_6_33_port, 
                           shift_in(32) => negative_inputs_6_32_port, 
                           shift_in(31) => negative_inputs_6_31_port, 
                           shift_in(30) => negative_inputs_6_30_port, 
                           shift_in(29) => negative_inputs_6_29_port, 
                           shift_in(28) => negative_inputs_6_28_port, 
                           shift_in(27) => negative_inputs_6_27_port, 
                           shift_in(26) => negative_inputs_6_26_port, 
                           shift_in(25) => negative_inputs_6_25_port, 
                           shift_in(24) => negative_inputs_6_24_port, 
                           shift_in(23) => negative_inputs_6_23_port, 
                           shift_in(22) => negative_inputs_6_22_port, 
                           shift_in(21) => negative_inputs_6_21_port, 
                           shift_in(20) => negative_inputs_6_20_port, 
                           shift_in(19) => negative_inputs_6_19_port, 
                           shift_in(18) => negative_inputs_6_18_port, 
                           shift_in(17) => negative_inputs_6_17_port, 
                           shift_in(16) => negative_inputs_6_16_port, 
                           shift_in(15) => negative_inputs_6_15_port, 
                           shift_in(14) => negative_inputs_6_14_port, 
                           shift_in(13) => negative_inputs_6_13_port, 
                           shift_in(12) => negative_inputs_6_12_port, 
                           shift_in(11) => negative_inputs_6_11_port, 
                           shift_in(10) => negative_inputs_6_10_port, 
                           shift_in(9) => negative_inputs_6_9_port, shift_in(8)
                           => negative_inputs_6_8_port, shift_in(7) => 
                           negative_inputs_6_7_port, shift_in(6) => 
                           negative_inputs_6_6_port, shift_in(5) => 
                           negative_inputs_6_5_port, shift_in(4) => 
                           negative_inputs_6_4_port, shift_in(3) => 
                           negative_inputs_6_3_port, shift_in(2) => 
                           negative_inputs_6_2_port, shift_in(1) => 
                           negative_inputs_6_1_port, shift_in(0) => n9, 
                           shift_out(63) => negative_inputs_7_63_port, 
                           shift_out(62) => negative_inputs_7_62_port, 
                           shift_out(61) => negative_inputs_7_61_port, 
                           shift_out(60) => negative_inputs_7_60_port, 
                           shift_out(59) => negative_inputs_7_59_port, 
                           shift_out(58) => negative_inputs_7_58_port, 
                           shift_out(57) => negative_inputs_7_57_port, 
                           shift_out(56) => negative_inputs_7_56_port, 
                           shift_out(55) => negative_inputs_7_55_port, 
                           shift_out(54) => negative_inputs_7_54_port, 
                           shift_out(53) => negative_inputs_7_53_port, 
                           shift_out(52) => negative_inputs_7_52_port, 
                           shift_out(51) => negative_inputs_7_51_port, 
                           shift_out(50) => negative_inputs_7_50_port, 
                           shift_out(49) => negative_inputs_7_49_port, 
                           shift_out(48) => negative_inputs_7_48_port, 
                           shift_out(47) => negative_inputs_7_47_port, 
                           shift_out(46) => negative_inputs_7_46_port, 
                           shift_out(45) => negative_inputs_7_45_port, 
                           shift_out(44) => negative_inputs_7_44_port, 
                           shift_out(43) => negative_inputs_7_43_port, 
                           shift_out(42) => negative_inputs_7_42_port, 
                           shift_out(41) => negative_inputs_7_41_port, 
                           shift_out(40) => negative_inputs_7_40_port, 
                           shift_out(39) => negative_inputs_7_39_port, 
                           shift_out(38) => negative_inputs_7_38_port, 
                           shift_out(37) => negative_inputs_7_37_port, 
                           shift_out(36) => negative_inputs_7_36_port, 
                           shift_out(35) => negative_inputs_7_35_port, 
                           shift_out(34) => negative_inputs_7_34_port, 
                           shift_out(33) => negative_inputs_7_33_port, 
                           shift_out(32) => negative_inputs_7_32_port, 
                           shift_out(31) => negative_inputs_7_31_port, 
                           shift_out(30) => negative_inputs_7_30_port, 
                           shift_out(29) => negative_inputs_7_29_port, 
                           shift_out(28) => negative_inputs_7_28_port, 
                           shift_out(27) => negative_inputs_7_27_port, 
                           shift_out(26) => negative_inputs_7_26_port, 
                           shift_out(25) => negative_inputs_7_25_port, 
                           shift_out(24) => negative_inputs_7_24_port, 
                           shift_out(23) => negative_inputs_7_23_port, 
                           shift_out(22) => negative_inputs_7_22_port, 
                           shift_out(21) => negative_inputs_7_21_port, 
                           shift_out(20) => negative_inputs_7_20_port, 
                           shift_out(19) => negative_inputs_7_19_port, 
                           shift_out(18) => negative_inputs_7_18_port, 
                           shift_out(17) => negative_inputs_7_17_port, 
                           shift_out(16) => negative_inputs_7_16_port, 
                           shift_out(15) => negative_inputs_7_15_port, 
                           shift_out(14) => negative_inputs_7_14_port, 
                           shift_out(13) => negative_inputs_7_13_port, 
                           shift_out(12) => negative_inputs_7_12_port, 
                           shift_out(11) => negative_inputs_7_11_port, 
                           shift_out(10) => negative_inputs_7_10_port, 
                           shift_out(9) => negative_inputs_7_9_port, 
                           shift_out(8) => negative_inputs_7_8_port, 
                           shift_out(7) => negative_inputs_7_7_port, 
                           shift_out(6) => negative_inputs_7_6_port, 
                           shift_out(5) => negative_inputs_7_5_port, 
                           shift_out(4) => negative_inputs_7_4_port, 
                           shift_out(3) => negative_inputs_7_3_port, 
                           shift_out(2) => negative_inputs_7_2_port, 
                           shift_out(1) => negative_inputs_7_1_port, 
                           shift_out(0) => n_1102);
   shifted_neg_8 : leftshifter_NbitShifter64_24 port map( shift_in(63) => 
                           negative_inputs_7_63_port, shift_in(62) => 
                           negative_inputs_7_62_port, shift_in(61) => 
                           negative_inputs_7_61_port, shift_in(60) => 
                           negative_inputs_7_60_port, shift_in(59) => 
                           negative_inputs_7_59_port, shift_in(58) => 
                           negative_inputs_7_58_port, shift_in(57) => 
                           negative_inputs_7_57_port, shift_in(56) => 
                           negative_inputs_7_56_port, shift_in(55) => 
                           negative_inputs_7_55_port, shift_in(54) => 
                           negative_inputs_7_54_port, shift_in(53) => 
                           negative_inputs_7_53_port, shift_in(52) => 
                           negative_inputs_7_52_port, shift_in(51) => 
                           negative_inputs_7_51_port, shift_in(50) => 
                           negative_inputs_7_50_port, shift_in(49) => 
                           negative_inputs_7_49_port, shift_in(48) => 
                           negative_inputs_7_48_port, shift_in(47) => 
                           negative_inputs_7_47_port, shift_in(46) => 
                           negative_inputs_7_46_port, shift_in(45) => 
                           negative_inputs_7_45_port, shift_in(44) => 
                           negative_inputs_7_44_port, shift_in(43) => 
                           negative_inputs_7_43_port, shift_in(42) => 
                           negative_inputs_7_42_port, shift_in(41) => 
                           negative_inputs_7_41_port, shift_in(40) => 
                           negative_inputs_7_40_port, shift_in(39) => n137, 
                           shift_in(38) => n135, shift_in(37) => n133, 
                           shift_in(36) => n131, shift_in(35) => n129, 
                           shift_in(34) => n127, shift_in(33) => n125, 
                           shift_in(32) => n123, shift_in(31) => n121, 
                           shift_in(30) => n119, shift_in(29) => n117, 
                           shift_in(28) => n115, shift_in(27) => n113, 
                           shift_in(26) => n111, shift_in(25) => n109, 
                           shift_in(24) => n107, shift_in(23) => n105, 
                           shift_in(22) => n103, shift_in(21) => n101, 
                           shift_in(20) => n99, shift_in(19) => n97, 
                           shift_in(18) => n95, shift_in(17) => n93, 
                           shift_in(16) => n91, shift_in(15) => n89, 
                           shift_in(14) => n87, shift_in(13) => n85, 
                           shift_in(12) => n83, shift_in(11) => n81, 
                           shift_in(10) => n79, shift_in(9) => n77, shift_in(8)
                           => n75, shift_in(7) => n73, shift_in(6) => 
                           negative_inputs_7_6_port, shift_in(5) => 
                           negative_inputs_7_5_port, shift_in(4) => 
                           negative_inputs_7_4_port, shift_in(3) => 
                           negative_inputs_7_3_port, shift_in(2) => 
                           negative_inputs_7_2_port, shift_in(1) => 
                           negative_inputs_7_1_port, shift_in(0) => n9, 
                           shift_out(63) => negative_inputs_8_63_port, 
                           shift_out(62) => negative_inputs_8_62_port, 
                           shift_out(61) => negative_inputs_8_61_port, 
                           shift_out(60) => negative_inputs_8_60_port, 
                           shift_out(59) => negative_inputs_8_59_port, 
                           shift_out(58) => negative_inputs_8_58_port, 
                           shift_out(57) => negative_inputs_8_57_port, 
                           shift_out(56) => negative_inputs_8_56_port, 
                           shift_out(55) => negative_inputs_8_55_port, 
                           shift_out(54) => negative_inputs_8_54_port, 
                           shift_out(53) => negative_inputs_8_53_port, 
                           shift_out(52) => negative_inputs_8_52_port, 
                           shift_out(51) => negative_inputs_8_51_port, 
                           shift_out(50) => negative_inputs_8_50_port, 
                           shift_out(49) => negative_inputs_8_49_port, 
                           shift_out(48) => negative_inputs_8_48_port, 
                           shift_out(47) => negative_inputs_8_47_port, 
                           shift_out(46) => negative_inputs_8_46_port, 
                           shift_out(45) => negative_inputs_8_45_port, 
                           shift_out(44) => negative_inputs_8_44_port, 
                           shift_out(43) => negative_inputs_8_43_port, 
                           shift_out(42) => negative_inputs_8_42_port, 
                           shift_out(41) => negative_inputs_8_41_port, 
                           shift_out(40) => negative_inputs_8_40_port, 
                           shift_out(39) => negative_inputs_8_39_port, 
                           shift_out(38) => negative_inputs_8_38_port, 
                           shift_out(37) => negative_inputs_8_37_port, 
                           shift_out(36) => negative_inputs_8_36_port, 
                           shift_out(35) => negative_inputs_8_35_port, 
                           shift_out(34) => negative_inputs_8_34_port, 
                           shift_out(33) => negative_inputs_8_33_port, 
                           shift_out(32) => negative_inputs_8_32_port, 
                           shift_out(31) => negative_inputs_8_31_port, 
                           shift_out(30) => negative_inputs_8_30_port, 
                           shift_out(29) => negative_inputs_8_29_port, 
                           shift_out(28) => negative_inputs_8_28_port, 
                           shift_out(27) => negative_inputs_8_27_port, 
                           shift_out(26) => negative_inputs_8_26_port, 
                           shift_out(25) => negative_inputs_8_25_port, 
                           shift_out(24) => negative_inputs_8_24_port, 
                           shift_out(23) => negative_inputs_8_23_port, 
                           shift_out(22) => negative_inputs_8_22_port, 
                           shift_out(21) => negative_inputs_8_21_port, 
                           shift_out(20) => negative_inputs_8_20_port, 
                           shift_out(19) => negative_inputs_8_19_port, 
                           shift_out(18) => negative_inputs_8_18_port, 
                           shift_out(17) => negative_inputs_8_17_port, 
                           shift_out(16) => negative_inputs_8_16_port, 
                           shift_out(15) => negative_inputs_8_15_port, 
                           shift_out(14) => negative_inputs_8_14_port, 
                           shift_out(13) => negative_inputs_8_13_port, 
                           shift_out(12) => negative_inputs_8_12_port, 
                           shift_out(11) => negative_inputs_8_11_port, 
                           shift_out(10) => negative_inputs_8_10_port, 
                           shift_out(9) => negative_inputs_8_9_port, 
                           shift_out(8) => negative_inputs_8_8_port, 
                           shift_out(7) => negative_inputs_8_7_port, 
                           shift_out(6) => negative_inputs_8_6_port, 
                           shift_out(5) => negative_inputs_8_5_port, 
                           shift_out(4) => negative_inputs_8_4_port, 
                           shift_out(3) => negative_inputs_8_3_port, 
                           shift_out(2) => negative_inputs_8_2_port, 
                           shift_out(1) => negative_inputs_8_1_port, 
                           shift_out(0) => n_1103);
   shifted_neg_9 : leftshifter_NbitShifter64_23 port map( shift_in(63) => 
                           negative_inputs_8_63_port, shift_in(62) => 
                           negative_inputs_8_62_port, shift_in(61) => 
                           negative_inputs_8_61_port, shift_in(60) => 
                           negative_inputs_8_60_port, shift_in(59) => 
                           negative_inputs_8_59_port, shift_in(58) => 
                           negative_inputs_8_58_port, shift_in(57) => 
                           negative_inputs_8_57_port, shift_in(56) => 
                           negative_inputs_8_56_port, shift_in(55) => 
                           negative_inputs_8_55_port, shift_in(54) => 
                           negative_inputs_8_54_port, shift_in(53) => 
                           negative_inputs_8_53_port, shift_in(52) => 
                           negative_inputs_8_52_port, shift_in(51) => 
                           negative_inputs_8_51_port, shift_in(50) => 
                           negative_inputs_8_50_port, shift_in(49) => 
                           negative_inputs_8_49_port, shift_in(48) => n153, 
                           shift_in(47) => negative_inputs_8_47_port, 
                           shift_in(46) => negative_inputs_8_46_port, 
                           shift_in(45) => negative_inputs_8_45_port, 
                           shift_in(44) => negative_inputs_8_44_port, 
                           shift_in(43) => negative_inputs_8_43_port, 
                           shift_in(42) => negative_inputs_8_42_port, 
                           shift_in(41) => negative_inputs_8_41_port, 
                           shift_in(40) => negative_inputs_8_40_port, 
                           shift_in(39) => negative_inputs_8_39_port, 
                           shift_in(38) => negative_inputs_8_38_port, 
                           shift_in(37) => negative_inputs_8_37_port, 
                           shift_in(36) => negative_inputs_8_36_port, 
                           shift_in(35) => negative_inputs_8_35_port, 
                           shift_in(34) => negative_inputs_8_34_port, 
                           shift_in(33) => negative_inputs_8_33_port, 
                           shift_in(32) => negative_inputs_8_32_port, 
                           shift_in(31) => negative_inputs_8_31_port, 
                           shift_in(30) => negative_inputs_8_30_port, 
                           shift_in(29) => negative_inputs_8_29_port, 
                           shift_in(28) => negative_inputs_8_28_port, 
                           shift_in(27) => negative_inputs_8_27_port, 
                           shift_in(26) => negative_inputs_8_26_port, 
                           shift_in(25) => negative_inputs_8_25_port, 
                           shift_in(24) => negative_inputs_8_24_port, 
                           shift_in(23) => negative_inputs_8_23_port, 
                           shift_in(22) => negative_inputs_8_22_port, 
                           shift_in(21) => negative_inputs_8_21_port, 
                           shift_in(20) => negative_inputs_8_20_port, 
                           shift_in(19) => negative_inputs_8_19_port, 
                           shift_in(18) => negative_inputs_8_18_port, 
                           shift_in(17) => negative_inputs_8_17_port, 
                           shift_in(16) => negative_inputs_8_16_port, 
                           shift_in(15) => negative_inputs_8_15_port, 
                           shift_in(14) => negative_inputs_8_14_port, 
                           shift_in(13) => negative_inputs_8_13_port, 
                           shift_in(12) => negative_inputs_8_12_port, 
                           shift_in(11) => negative_inputs_8_11_port, 
                           shift_in(10) => negative_inputs_8_10_port, 
                           shift_in(9) => negative_inputs_8_9_port, shift_in(8)
                           => negative_inputs_8_8_port, shift_in(7) => 
                           negative_inputs_8_7_port, shift_in(6) => 
                           negative_inputs_8_6_port, shift_in(5) => 
                           negative_inputs_8_5_port, shift_in(4) => 
                           negative_inputs_8_4_port, shift_in(3) => 
                           negative_inputs_8_3_port, shift_in(2) => 
                           negative_inputs_8_2_port, shift_in(1) => 
                           negative_inputs_8_1_port, shift_in(0) => n9, 
                           shift_out(63) => negative_inputs_9_63_port, 
                           shift_out(62) => negative_inputs_9_62_port, 
                           shift_out(61) => negative_inputs_9_61_port, 
                           shift_out(60) => negative_inputs_9_60_port, 
                           shift_out(59) => negative_inputs_9_59_port, 
                           shift_out(58) => negative_inputs_9_58_port, 
                           shift_out(57) => negative_inputs_9_57_port, 
                           shift_out(56) => negative_inputs_9_56_port, 
                           shift_out(55) => negative_inputs_9_55_port, 
                           shift_out(54) => negative_inputs_9_54_port, 
                           shift_out(53) => negative_inputs_9_53_port, 
                           shift_out(52) => negative_inputs_9_52_port, 
                           shift_out(51) => negative_inputs_9_51_port, 
                           shift_out(50) => negative_inputs_9_50_port, 
                           shift_out(49) => negative_inputs_9_49_port, 
                           shift_out(48) => negative_inputs_9_48_port, 
                           shift_out(47) => negative_inputs_9_47_port, 
                           shift_out(46) => negative_inputs_9_46_port, 
                           shift_out(45) => negative_inputs_9_45_port, 
                           shift_out(44) => negative_inputs_9_44_port, 
                           shift_out(43) => negative_inputs_9_43_port, 
                           shift_out(42) => negative_inputs_9_42_port, 
                           shift_out(41) => negative_inputs_9_41_port, 
                           shift_out(40) => negative_inputs_9_40_port, 
                           shift_out(39) => negative_inputs_9_39_port, 
                           shift_out(38) => negative_inputs_9_38_port, 
                           shift_out(37) => negative_inputs_9_37_port, 
                           shift_out(36) => negative_inputs_9_36_port, 
                           shift_out(35) => negative_inputs_9_35_port, 
                           shift_out(34) => negative_inputs_9_34_port, 
                           shift_out(33) => negative_inputs_9_33_port, 
                           shift_out(32) => negative_inputs_9_32_port, 
                           shift_out(31) => negative_inputs_9_31_port, 
                           shift_out(30) => negative_inputs_9_30_port, 
                           shift_out(29) => negative_inputs_9_29_port, 
                           shift_out(28) => negative_inputs_9_28_port, 
                           shift_out(27) => negative_inputs_9_27_port, 
                           shift_out(26) => negative_inputs_9_26_port, 
                           shift_out(25) => negative_inputs_9_25_port, 
                           shift_out(24) => negative_inputs_9_24_port, 
                           shift_out(23) => negative_inputs_9_23_port, 
                           shift_out(22) => negative_inputs_9_22_port, 
                           shift_out(21) => negative_inputs_9_21_port, 
                           shift_out(20) => negative_inputs_9_20_port, 
                           shift_out(19) => negative_inputs_9_19_port, 
                           shift_out(18) => negative_inputs_9_18_port, 
                           shift_out(17) => negative_inputs_9_17_port, 
                           shift_out(16) => negative_inputs_9_16_port, 
                           shift_out(15) => negative_inputs_9_15_port, 
                           shift_out(14) => negative_inputs_9_14_port, 
                           shift_out(13) => negative_inputs_9_13_port, 
                           shift_out(12) => negative_inputs_9_12_port, 
                           shift_out(11) => negative_inputs_9_11_port, 
                           shift_out(10) => negative_inputs_9_10_port, 
                           shift_out(9) => negative_inputs_9_9_port, 
                           shift_out(8) => negative_inputs_9_8_port, 
                           shift_out(7) => negative_inputs_9_7_port, 
                           shift_out(6) => negative_inputs_9_6_port, 
                           shift_out(5) => negative_inputs_9_5_port, 
                           shift_out(4) => negative_inputs_9_4_port, 
                           shift_out(3) => negative_inputs_9_3_port, 
                           shift_out(2) => negative_inputs_9_2_port, 
                           shift_out(1) => negative_inputs_9_1_port, 
                           shift_out(0) => n_1104);
   shifted_neg_10 : leftshifter_NbitShifter64_22 port map( shift_in(63) => 
                           negative_inputs_9_63_port, shift_in(62) => 
                           negative_inputs_9_62_port, shift_in(61) => 
                           negative_inputs_9_61_port, shift_in(60) => 
                           negative_inputs_9_60_port, shift_in(59) => 
                           negative_inputs_9_59_port, shift_in(58) => 
                           negative_inputs_9_58_port, shift_in(57) => 
                           negative_inputs_9_57_port, shift_in(56) => 
                           negative_inputs_9_56_port, shift_in(55) => 
                           negative_inputs_9_55_port, shift_in(54) => 
                           negative_inputs_9_54_port, shift_in(53) => 
                           negative_inputs_9_53_port, shift_in(52) => 
                           negative_inputs_9_52_port, shift_in(51) => 
                           negative_inputs_9_51_port, shift_in(50) => 
                           negative_inputs_9_50_port, shift_in(49) => 
                           negative_inputs_9_49_port, shift_in(48) => n152, 
                           shift_in(47) => negative_inputs_9_47_port, 
                           shift_in(46) => negative_inputs_9_46_port, 
                           shift_in(45) => negative_inputs_9_45_port, 
                           shift_in(44) => negative_inputs_9_44_port, 
                           shift_in(43) => negative_inputs_9_43_port, 
                           shift_in(42) => negative_inputs_9_42_port, 
                           shift_in(41) => negative_inputs_9_41_port, 
                           shift_in(40) => negative_inputs_9_40_port, 
                           shift_in(39) => negative_inputs_9_39_port, 
                           shift_in(38) => negative_inputs_9_38_port, 
                           shift_in(37) => negative_inputs_9_37_port, 
                           shift_in(36) => negative_inputs_9_36_port, 
                           shift_in(35) => negative_inputs_9_35_port, 
                           shift_in(34) => negative_inputs_9_34_port, 
                           shift_in(33) => negative_inputs_9_33_port, 
                           shift_in(32) => negative_inputs_9_32_port, 
                           shift_in(31) => negative_inputs_9_31_port, 
                           shift_in(30) => negative_inputs_9_30_port, 
                           shift_in(29) => negative_inputs_9_29_port, 
                           shift_in(28) => negative_inputs_9_28_port, 
                           shift_in(27) => negative_inputs_9_27_port, 
                           shift_in(26) => negative_inputs_9_26_port, 
                           shift_in(25) => negative_inputs_9_25_port, 
                           shift_in(24) => negative_inputs_9_24_port, 
                           shift_in(23) => negative_inputs_9_23_port, 
                           shift_in(22) => negative_inputs_9_22_port, 
                           shift_in(21) => negative_inputs_9_21_port, 
                           shift_in(20) => negative_inputs_9_20_port, 
                           shift_in(19) => negative_inputs_9_19_port, 
                           shift_in(18) => negative_inputs_9_18_port, 
                           shift_in(17) => negative_inputs_9_17_port, 
                           shift_in(16) => negative_inputs_9_16_port, 
                           shift_in(15) => negative_inputs_9_15_port, 
                           shift_in(14) => negative_inputs_9_14_port, 
                           shift_in(13) => negative_inputs_9_13_port, 
                           shift_in(12) => negative_inputs_9_12_port, 
                           shift_in(11) => negative_inputs_9_11_port, 
                           shift_in(10) => negative_inputs_9_10_port, 
                           shift_in(9) => negative_inputs_9_9_port, shift_in(8)
                           => negative_inputs_9_8_port, shift_in(7) => 
                           negative_inputs_9_7_port, shift_in(6) => 
                           negative_inputs_9_6_port, shift_in(5) => 
                           negative_inputs_9_5_port, shift_in(4) => 
                           negative_inputs_9_4_port, shift_in(3) => 
                           negative_inputs_9_3_port, shift_in(2) => 
                           negative_inputs_9_2_port, shift_in(1) => 
                           negative_inputs_9_1_port, shift_in(0) => n9, 
                           shift_out(63) => negative_inputs_10_63_port, 
                           shift_out(62) => negative_inputs_10_62_port, 
                           shift_out(61) => negative_inputs_10_61_port, 
                           shift_out(60) => negative_inputs_10_60_port, 
                           shift_out(59) => negative_inputs_10_59_port, 
                           shift_out(58) => negative_inputs_10_58_port, 
                           shift_out(57) => negative_inputs_10_57_port, 
                           shift_out(56) => negative_inputs_10_56_port, 
                           shift_out(55) => negative_inputs_10_55_port, 
                           shift_out(54) => negative_inputs_10_54_port, 
                           shift_out(53) => negative_inputs_10_53_port, 
                           shift_out(52) => negative_inputs_10_52_port, 
                           shift_out(51) => negative_inputs_10_51_port, 
                           shift_out(50) => negative_inputs_10_50_port, 
                           shift_out(49) => negative_inputs_10_49_port, 
                           shift_out(48) => negative_inputs_10_48_port, 
                           shift_out(47) => negative_inputs_10_47_port, 
                           shift_out(46) => negative_inputs_10_46_port, 
                           shift_out(45) => negative_inputs_10_45_port, 
                           shift_out(44) => negative_inputs_10_44_port, 
                           shift_out(43) => negative_inputs_10_43_port, 
                           shift_out(42) => negative_inputs_10_42_port, 
                           shift_out(41) => negative_inputs_10_41_port, 
                           shift_out(40) => negative_inputs_10_40_port, 
                           shift_out(39) => negative_inputs_10_39_port, 
                           shift_out(38) => negative_inputs_10_38_port, 
                           shift_out(37) => negative_inputs_10_37_port, 
                           shift_out(36) => negative_inputs_10_36_port, 
                           shift_out(35) => negative_inputs_10_35_port, 
                           shift_out(34) => negative_inputs_10_34_port, 
                           shift_out(33) => negative_inputs_10_33_port, 
                           shift_out(32) => negative_inputs_10_32_port, 
                           shift_out(31) => negative_inputs_10_31_port, 
                           shift_out(30) => negative_inputs_10_30_port, 
                           shift_out(29) => negative_inputs_10_29_port, 
                           shift_out(28) => negative_inputs_10_28_port, 
                           shift_out(27) => negative_inputs_10_27_port, 
                           shift_out(26) => negative_inputs_10_26_port, 
                           shift_out(25) => negative_inputs_10_25_port, 
                           shift_out(24) => negative_inputs_10_24_port, 
                           shift_out(23) => negative_inputs_10_23_port, 
                           shift_out(22) => negative_inputs_10_22_port, 
                           shift_out(21) => negative_inputs_10_21_port, 
                           shift_out(20) => negative_inputs_10_20_port, 
                           shift_out(19) => negative_inputs_10_19_port, 
                           shift_out(18) => negative_inputs_10_18_port, 
                           shift_out(17) => negative_inputs_10_17_port, 
                           shift_out(16) => negative_inputs_10_16_port, 
                           shift_out(15) => negative_inputs_10_15_port, 
                           shift_out(14) => negative_inputs_10_14_port, 
                           shift_out(13) => negative_inputs_10_13_port, 
                           shift_out(12) => negative_inputs_10_12_port, 
                           shift_out(11) => negative_inputs_10_11_port, 
                           shift_out(10) => negative_inputs_10_10_port, 
                           shift_out(9) => negative_inputs_10_9_port, 
                           shift_out(8) => negative_inputs_10_8_port, 
                           shift_out(7) => negative_inputs_10_7_port, 
                           shift_out(6) => negative_inputs_10_6_port, 
                           shift_out(5) => negative_inputs_10_5_port, 
                           shift_out(4) => negative_inputs_10_4_port, 
                           shift_out(3) => negative_inputs_10_3_port, 
                           shift_out(2) => negative_inputs_10_2_port, 
                           shift_out(1) => negative_inputs_10_1_port, 
                           shift_out(0) => n_1105);
   shifted_neg_11 : leftshifter_NbitShifter64_21 port map( shift_in(63) => 
                           negative_inputs_10_63_port, shift_in(62) => 
                           negative_inputs_10_62_port, shift_in(61) => 
                           negative_inputs_10_61_port, shift_in(60) => 
                           negative_inputs_10_60_port, shift_in(59) => 
                           negative_inputs_10_59_port, shift_in(58) => 
                           negative_inputs_10_58_port, shift_in(57) => 
                           negative_inputs_10_57_port, shift_in(56) => 
                           negative_inputs_10_56_port, shift_in(55) => 
                           negative_inputs_10_55_port, shift_in(54) => 
                           negative_inputs_10_54_port, shift_in(53) => 
                           negative_inputs_10_53_port, shift_in(52) => 
                           negative_inputs_10_52_port, shift_in(51) => 
                           negative_inputs_10_51_port, shift_in(50) => 
                           negative_inputs_10_50_port, shift_in(49) => 
                           negative_inputs_10_49_port, shift_in(48) => n150, 
                           shift_in(47) => negative_inputs_10_47_port, 
                           shift_in(46) => negative_inputs_10_46_port, 
                           shift_in(45) => negative_inputs_10_45_port, 
                           shift_in(44) => negative_inputs_10_44_port, 
                           shift_in(43) => negative_inputs_10_43_port, 
                           shift_in(42) => negative_inputs_10_42_port, 
                           shift_in(41) => negative_inputs_10_41_port, 
                           shift_in(40) => negative_inputs_10_40_port, 
                           shift_in(39) => negative_inputs_10_39_port, 
                           shift_in(38) => negative_inputs_10_38_port, 
                           shift_in(37) => negative_inputs_10_37_port, 
                           shift_in(36) => negative_inputs_10_36_port, 
                           shift_in(35) => negative_inputs_10_35_port, 
                           shift_in(34) => negative_inputs_10_34_port, 
                           shift_in(33) => negative_inputs_10_33_port, 
                           shift_in(32) => negative_inputs_10_32_port, 
                           shift_in(31) => negative_inputs_10_31_port, 
                           shift_in(30) => negative_inputs_10_30_port, 
                           shift_in(29) => negative_inputs_10_29_port, 
                           shift_in(28) => negative_inputs_10_28_port, 
                           shift_in(27) => negative_inputs_10_27_port, 
                           shift_in(26) => negative_inputs_10_26_port, 
                           shift_in(25) => negative_inputs_10_25_port, 
                           shift_in(24) => negative_inputs_10_24_port, 
                           shift_in(23) => negative_inputs_10_23_port, 
                           shift_in(22) => negative_inputs_10_22_port, 
                           shift_in(21) => negative_inputs_10_21_port, 
                           shift_in(20) => negative_inputs_10_20_port, 
                           shift_in(19) => negative_inputs_10_19_port, 
                           shift_in(18) => negative_inputs_10_18_port, 
                           shift_in(17) => negative_inputs_10_17_port, 
                           shift_in(16) => negative_inputs_10_16_port, 
                           shift_in(15) => negative_inputs_10_15_port, 
                           shift_in(14) => negative_inputs_10_14_port, 
                           shift_in(13) => negative_inputs_10_13_port, 
                           shift_in(12) => negative_inputs_10_12_port, 
                           shift_in(11) => negative_inputs_10_11_port, 
                           shift_in(10) => negative_inputs_10_10_port, 
                           shift_in(9) => negative_inputs_10_9_port, 
                           shift_in(8) => negative_inputs_10_8_port, 
                           shift_in(7) => negative_inputs_10_7_port, 
                           shift_in(6) => negative_inputs_10_6_port, 
                           shift_in(5) => negative_inputs_10_5_port, 
                           shift_in(4) => negative_inputs_10_4_port, 
                           shift_in(3) => negative_inputs_10_3_port, 
                           shift_in(2) => negative_inputs_10_2_port, 
                           shift_in(1) => negative_inputs_10_1_port, 
                           shift_in(0) => n9, shift_out(63) => 
                           negative_inputs_11_63_port, shift_out(62) => 
                           negative_inputs_11_62_port, shift_out(61) => 
                           negative_inputs_11_61_port, shift_out(60) => 
                           negative_inputs_11_60_port, shift_out(59) => 
                           negative_inputs_11_59_port, shift_out(58) => 
                           negative_inputs_11_58_port, shift_out(57) => 
                           negative_inputs_11_57_port, shift_out(56) => 
                           negative_inputs_11_56_port, shift_out(55) => 
                           negative_inputs_11_55_port, shift_out(54) => 
                           negative_inputs_11_54_port, shift_out(53) => 
                           negative_inputs_11_53_port, shift_out(52) => 
                           negative_inputs_11_52_port, shift_out(51) => 
                           negative_inputs_11_51_port, shift_out(50) => 
                           negative_inputs_11_50_port, shift_out(49) => 
                           negative_inputs_11_49_port, shift_out(48) => 
                           negative_inputs_11_48_port, shift_out(47) => 
                           negative_inputs_11_47_port, shift_out(46) => 
                           negative_inputs_11_46_port, shift_out(45) => 
                           negative_inputs_11_45_port, shift_out(44) => 
                           negative_inputs_11_44_port, shift_out(43) => 
                           negative_inputs_11_43_port, shift_out(42) => 
                           negative_inputs_11_42_port, shift_out(41) => 
                           negative_inputs_11_41_port, shift_out(40) => 
                           negative_inputs_11_40_port, shift_out(39) => 
                           negative_inputs_11_39_port, shift_out(38) => 
                           negative_inputs_11_38_port, shift_out(37) => 
                           negative_inputs_11_37_port, shift_out(36) => 
                           negative_inputs_11_36_port, shift_out(35) => 
                           negative_inputs_11_35_port, shift_out(34) => 
                           negative_inputs_11_34_port, shift_out(33) => 
                           negative_inputs_11_33_port, shift_out(32) => 
                           negative_inputs_11_32_port, shift_out(31) => 
                           negative_inputs_11_31_port, shift_out(30) => 
                           negative_inputs_11_30_port, shift_out(29) => 
                           negative_inputs_11_29_port, shift_out(28) => 
                           negative_inputs_11_28_port, shift_out(27) => 
                           negative_inputs_11_27_port, shift_out(26) => 
                           negative_inputs_11_26_port, shift_out(25) => 
                           negative_inputs_11_25_port, shift_out(24) => 
                           negative_inputs_11_24_port, shift_out(23) => 
                           negative_inputs_11_23_port, shift_out(22) => 
                           negative_inputs_11_22_port, shift_out(21) => 
                           negative_inputs_11_21_port, shift_out(20) => 
                           negative_inputs_11_20_port, shift_out(19) => 
                           negative_inputs_11_19_port, shift_out(18) => 
                           negative_inputs_11_18_port, shift_out(17) => 
                           negative_inputs_11_17_port, shift_out(16) => 
                           negative_inputs_11_16_port, shift_out(15) => 
                           negative_inputs_11_15_port, shift_out(14) => 
                           negative_inputs_11_14_port, shift_out(13) => 
                           negative_inputs_11_13_port, shift_out(12) => 
                           negative_inputs_11_12_port, shift_out(11) => 
                           negative_inputs_11_11_port, shift_out(10) => 
                           negative_inputs_11_10_port, shift_out(9) => 
                           negative_inputs_11_9_port, shift_out(8) => 
                           negative_inputs_11_8_port, shift_out(7) => 
                           negative_inputs_11_7_port, shift_out(6) => 
                           negative_inputs_11_6_port, shift_out(5) => 
                           negative_inputs_11_5_port, shift_out(4) => 
                           negative_inputs_11_4_port, shift_out(3) => 
                           negative_inputs_11_3_port, shift_out(2) => 
                           negative_inputs_11_2_port, shift_out(1) => 
                           negative_inputs_11_1_port, shift_out(0) => n_1106);
   shifted_neg_12 : leftshifter_NbitShifter64_20 port map( shift_in(63) => 
                           negative_inputs_11_63_port, shift_in(62) => 
                           negative_inputs_11_62_port, shift_in(61) => 
                           negative_inputs_11_61_port, shift_in(60) => 
                           negative_inputs_11_60_port, shift_in(59) => 
                           negative_inputs_11_59_port, shift_in(58) => 
                           negative_inputs_11_58_port, shift_in(57) => 
                           negative_inputs_11_57_port, shift_in(56) => 
                           negative_inputs_11_56_port, shift_in(55) => 
                           negative_inputs_11_55_port, shift_in(54) => 
                           negative_inputs_11_54_port, shift_in(53) => 
                           negative_inputs_11_53_port, shift_in(52) => 
                           negative_inputs_11_52_port, shift_in(51) => 
                           negative_inputs_11_51_port, shift_in(50) => 
                           negative_inputs_11_50_port, shift_in(49) => 
                           negative_inputs_11_49_port, shift_in(48) => n148, 
                           shift_in(47) => negative_inputs_11_47_port, 
                           shift_in(46) => negative_inputs_11_46_port, 
                           shift_in(45) => negative_inputs_11_45_port, 
                           shift_in(44) => negative_inputs_11_44_port, 
                           shift_in(43) => negative_inputs_11_43_port, 
                           shift_in(42) => negative_inputs_11_42_port, 
                           shift_in(41) => negative_inputs_11_41_port, 
                           shift_in(40) => negative_inputs_11_40_port, 
                           shift_in(39) => negative_inputs_11_39_port, 
                           shift_in(38) => negative_inputs_11_38_port, 
                           shift_in(37) => negative_inputs_11_37_port, 
                           shift_in(36) => negative_inputs_11_36_port, 
                           shift_in(35) => negative_inputs_11_35_port, 
                           shift_in(34) => negative_inputs_11_34_port, 
                           shift_in(33) => negative_inputs_11_33_port, 
                           shift_in(32) => negative_inputs_11_32_port, 
                           shift_in(31) => negative_inputs_11_31_port, 
                           shift_in(30) => negative_inputs_11_30_port, 
                           shift_in(29) => negative_inputs_11_29_port, 
                           shift_in(28) => negative_inputs_11_28_port, 
                           shift_in(27) => negative_inputs_11_27_port, 
                           shift_in(26) => negative_inputs_11_26_port, 
                           shift_in(25) => negative_inputs_11_25_port, 
                           shift_in(24) => negative_inputs_11_24_port, 
                           shift_in(23) => negative_inputs_11_23_port, 
                           shift_in(22) => negative_inputs_11_22_port, 
                           shift_in(21) => negative_inputs_11_21_port, 
                           shift_in(20) => negative_inputs_11_20_port, 
                           shift_in(19) => negative_inputs_11_19_port, 
                           shift_in(18) => negative_inputs_11_18_port, 
                           shift_in(17) => negative_inputs_11_17_port, 
                           shift_in(16) => negative_inputs_11_16_port, 
                           shift_in(15) => negative_inputs_11_15_port, 
                           shift_in(14) => negative_inputs_11_14_port, 
                           shift_in(13) => negative_inputs_11_13_port, 
                           shift_in(12) => negative_inputs_11_12_port, 
                           shift_in(11) => negative_inputs_11_11_port, 
                           shift_in(10) => negative_inputs_11_10_port, 
                           shift_in(9) => negative_inputs_11_9_port, 
                           shift_in(8) => negative_inputs_11_8_port, 
                           shift_in(7) => negative_inputs_11_7_port, 
                           shift_in(6) => negative_inputs_11_6_port, 
                           shift_in(5) => negative_inputs_11_5_port, 
                           shift_in(4) => negative_inputs_11_4_port, 
                           shift_in(3) => negative_inputs_11_3_port, 
                           shift_in(2) => negative_inputs_11_2_port, 
                           shift_in(1) => negative_inputs_11_1_port, 
                           shift_in(0) => n9, shift_out(63) => 
                           negative_inputs_12_63_port, shift_out(62) => 
                           negative_inputs_12_62_port, shift_out(61) => 
                           negative_inputs_12_61_port, shift_out(60) => 
                           negative_inputs_12_60_port, shift_out(59) => 
                           negative_inputs_12_59_port, shift_out(58) => 
                           negative_inputs_12_58_port, shift_out(57) => 
                           negative_inputs_12_57_port, shift_out(56) => 
                           negative_inputs_12_56_port, shift_out(55) => 
                           negative_inputs_12_55_port, shift_out(54) => 
                           negative_inputs_12_54_port, shift_out(53) => 
                           negative_inputs_12_53_port, shift_out(52) => 
                           negative_inputs_12_52_port, shift_out(51) => 
                           negative_inputs_12_51_port, shift_out(50) => 
                           negative_inputs_12_50_port, shift_out(49) => 
                           negative_inputs_12_49_port, shift_out(48) => 
                           negative_inputs_12_48_port, shift_out(47) => 
                           negative_inputs_12_47_port, shift_out(46) => 
                           negative_inputs_12_46_port, shift_out(45) => 
                           negative_inputs_12_45_port, shift_out(44) => 
                           negative_inputs_12_44_port, shift_out(43) => 
                           negative_inputs_12_43_port, shift_out(42) => 
                           negative_inputs_12_42_port, shift_out(41) => 
                           negative_inputs_12_41_port, shift_out(40) => 
                           negative_inputs_12_40_port, shift_out(39) => 
                           negative_inputs_12_39_port, shift_out(38) => 
                           negative_inputs_12_38_port, shift_out(37) => 
                           negative_inputs_12_37_port, shift_out(36) => 
                           negative_inputs_12_36_port, shift_out(35) => 
                           negative_inputs_12_35_port, shift_out(34) => 
                           negative_inputs_12_34_port, shift_out(33) => 
                           negative_inputs_12_33_port, shift_out(32) => 
                           negative_inputs_12_32_port, shift_out(31) => 
                           negative_inputs_12_31_port, shift_out(30) => 
                           negative_inputs_12_30_port, shift_out(29) => 
                           negative_inputs_12_29_port, shift_out(28) => 
                           negative_inputs_12_28_port, shift_out(27) => 
                           negative_inputs_12_27_port, shift_out(26) => 
                           negative_inputs_12_26_port, shift_out(25) => 
                           negative_inputs_12_25_port, shift_out(24) => 
                           negative_inputs_12_24_port, shift_out(23) => 
                           negative_inputs_12_23_port, shift_out(22) => 
                           negative_inputs_12_22_port, shift_out(21) => 
                           negative_inputs_12_21_port, shift_out(20) => 
                           negative_inputs_12_20_port, shift_out(19) => 
                           negative_inputs_12_19_port, shift_out(18) => 
                           negative_inputs_12_18_port, shift_out(17) => 
                           negative_inputs_12_17_port, shift_out(16) => 
                           negative_inputs_12_16_port, shift_out(15) => 
                           negative_inputs_12_15_port, shift_out(14) => 
                           negative_inputs_12_14_port, shift_out(13) => 
                           negative_inputs_12_13_port, shift_out(12) => 
                           negative_inputs_12_12_port, shift_out(11) => 
                           negative_inputs_12_11_port, shift_out(10) => 
                           negative_inputs_12_10_port, shift_out(9) => 
                           negative_inputs_12_9_port, shift_out(8) => 
                           negative_inputs_12_8_port, shift_out(7) => 
                           negative_inputs_12_7_port, shift_out(6) => 
                           negative_inputs_12_6_port, shift_out(5) => 
                           negative_inputs_12_5_port, shift_out(4) => 
                           negative_inputs_12_4_port, shift_out(3) => 
                           negative_inputs_12_3_port, shift_out(2) => 
                           negative_inputs_12_2_port, shift_out(1) => 
                           negative_inputs_12_1_port, shift_out(0) => n_1107);
   shifted_neg_13 : leftshifter_NbitShifter64_19 port map( shift_in(63) => 
                           negative_inputs_12_63_port, shift_in(62) => 
                           negative_inputs_12_62_port, shift_in(61) => 
                           negative_inputs_12_61_port, shift_in(60) => 
                           negative_inputs_12_60_port, shift_in(59) => 
                           negative_inputs_12_59_port, shift_in(58) => 
                           negative_inputs_12_58_port, shift_in(57) => 
                           negative_inputs_12_57_port, shift_in(56) => 
                           negative_inputs_12_56_port, shift_in(55) => 
                           negative_inputs_12_55_port, shift_in(54) => 
                           negative_inputs_12_54_port, shift_in(53) => 
                           negative_inputs_12_53_port, shift_in(52) => 
                           negative_inputs_12_52_port, shift_in(51) => 
                           negative_inputs_12_51_port, shift_in(50) => 
                           negative_inputs_12_50_port, shift_in(49) => 
                           negative_inputs_12_49_port, shift_in(48) => n146, 
                           shift_in(47) => negative_inputs_12_47_port, 
                           shift_in(46) => negative_inputs_12_46_port, 
                           shift_in(45) => negative_inputs_12_45_port, 
                           shift_in(44) => negative_inputs_12_44_port, 
                           shift_in(43) => negative_inputs_12_43_port, 
                           shift_in(42) => negative_inputs_12_42_port, 
                           shift_in(41) => negative_inputs_12_41_port, 
                           shift_in(40) => negative_inputs_12_40_port, 
                           shift_in(39) => negative_inputs_12_39_port, 
                           shift_in(38) => negative_inputs_12_38_port, 
                           shift_in(37) => negative_inputs_12_37_port, 
                           shift_in(36) => negative_inputs_12_36_port, 
                           shift_in(35) => negative_inputs_12_35_port, 
                           shift_in(34) => negative_inputs_12_34_port, 
                           shift_in(33) => negative_inputs_12_33_port, 
                           shift_in(32) => negative_inputs_12_32_port, 
                           shift_in(31) => negative_inputs_12_31_port, 
                           shift_in(30) => negative_inputs_12_30_port, 
                           shift_in(29) => negative_inputs_12_29_port, 
                           shift_in(28) => negative_inputs_12_28_port, 
                           shift_in(27) => negative_inputs_12_27_port, 
                           shift_in(26) => negative_inputs_12_26_port, 
                           shift_in(25) => negative_inputs_12_25_port, 
                           shift_in(24) => negative_inputs_12_24_port, 
                           shift_in(23) => negative_inputs_12_23_port, 
                           shift_in(22) => negative_inputs_12_22_port, 
                           shift_in(21) => negative_inputs_12_21_port, 
                           shift_in(20) => negative_inputs_12_20_port, 
                           shift_in(19) => negative_inputs_12_19_port, 
                           shift_in(18) => negative_inputs_12_18_port, 
                           shift_in(17) => negative_inputs_12_17_port, 
                           shift_in(16) => negative_inputs_12_16_port, 
                           shift_in(15) => negative_inputs_12_15_port, 
                           shift_in(14) => negative_inputs_12_14_port, 
                           shift_in(13) => negative_inputs_12_13_port, 
                           shift_in(12) => negative_inputs_12_12_port, 
                           shift_in(11) => negative_inputs_12_11_port, 
                           shift_in(10) => negative_inputs_12_10_port, 
                           shift_in(9) => negative_inputs_12_9_port, 
                           shift_in(8) => negative_inputs_12_8_port, 
                           shift_in(7) => negative_inputs_12_7_port, 
                           shift_in(6) => negative_inputs_12_6_port, 
                           shift_in(5) => negative_inputs_12_5_port, 
                           shift_in(4) => negative_inputs_12_4_port, 
                           shift_in(3) => negative_inputs_12_3_port, 
                           shift_in(2) => negative_inputs_12_2_port, 
                           shift_in(1) => negative_inputs_12_1_port, 
                           shift_in(0) => n9, shift_out(63) => 
                           negative_inputs_13_63_port, shift_out(62) => 
                           negative_inputs_13_62_port, shift_out(61) => 
                           negative_inputs_13_61_port, shift_out(60) => 
                           negative_inputs_13_60_port, shift_out(59) => 
                           negative_inputs_13_59_port, shift_out(58) => 
                           negative_inputs_13_58_port, shift_out(57) => 
                           negative_inputs_13_57_port, shift_out(56) => 
                           negative_inputs_13_56_port, shift_out(55) => 
                           negative_inputs_13_55_port, shift_out(54) => 
                           negative_inputs_13_54_port, shift_out(53) => 
                           negative_inputs_13_53_port, shift_out(52) => 
                           negative_inputs_13_52_port, shift_out(51) => 
                           negative_inputs_13_51_port, shift_out(50) => 
                           negative_inputs_13_50_port, shift_out(49) => 
                           negative_inputs_13_49_port, shift_out(48) => 
                           negative_inputs_13_48_port, shift_out(47) => 
                           negative_inputs_13_47_port, shift_out(46) => 
                           negative_inputs_13_46_port, shift_out(45) => 
                           negative_inputs_13_45_port, shift_out(44) => 
                           negative_inputs_13_44_port, shift_out(43) => 
                           negative_inputs_13_43_port, shift_out(42) => 
                           negative_inputs_13_42_port, shift_out(41) => 
                           negative_inputs_13_41_port, shift_out(40) => 
                           negative_inputs_13_40_port, shift_out(39) => 
                           negative_inputs_13_39_port, shift_out(38) => 
                           negative_inputs_13_38_port, shift_out(37) => 
                           negative_inputs_13_37_port, shift_out(36) => 
                           negative_inputs_13_36_port, shift_out(35) => 
                           negative_inputs_13_35_port, shift_out(34) => 
                           negative_inputs_13_34_port, shift_out(33) => 
                           negative_inputs_13_33_port, shift_out(32) => 
                           negative_inputs_13_32_port, shift_out(31) => 
                           negative_inputs_13_31_port, shift_out(30) => 
                           negative_inputs_13_30_port, shift_out(29) => 
                           negative_inputs_13_29_port, shift_out(28) => 
                           negative_inputs_13_28_port, shift_out(27) => 
                           negative_inputs_13_27_port, shift_out(26) => 
                           negative_inputs_13_26_port, shift_out(25) => 
                           negative_inputs_13_25_port, shift_out(24) => 
                           negative_inputs_13_24_port, shift_out(23) => 
                           negative_inputs_13_23_port, shift_out(22) => 
                           negative_inputs_13_22_port, shift_out(21) => 
                           negative_inputs_13_21_port, shift_out(20) => 
                           negative_inputs_13_20_port, shift_out(19) => 
                           negative_inputs_13_19_port, shift_out(18) => 
                           negative_inputs_13_18_port, shift_out(17) => 
                           negative_inputs_13_17_port, shift_out(16) => 
                           negative_inputs_13_16_port, shift_out(15) => 
                           negative_inputs_13_15_port, shift_out(14) => 
                           negative_inputs_13_14_port, shift_out(13) => 
                           negative_inputs_13_13_port, shift_out(12) => 
                           negative_inputs_13_12_port, shift_out(11) => 
                           negative_inputs_13_11_port, shift_out(10) => 
                           negative_inputs_13_10_port, shift_out(9) => 
                           negative_inputs_13_9_port, shift_out(8) => 
                           negative_inputs_13_8_port, shift_out(7) => 
                           negative_inputs_13_7_port, shift_out(6) => 
                           negative_inputs_13_6_port, shift_out(5) => 
                           negative_inputs_13_5_port, shift_out(4) => 
                           negative_inputs_13_4_port, shift_out(3) => 
                           negative_inputs_13_3_port, shift_out(2) => 
                           negative_inputs_13_2_port, shift_out(1) => 
                           negative_inputs_13_1_port, shift_out(0) => n_1108);
   shifted_neg_14 : leftshifter_NbitShifter64_18 port map( shift_in(63) => 
                           negative_inputs_13_63_port, shift_in(62) => 
                           negative_inputs_13_62_port, shift_in(61) => 
                           negative_inputs_13_61_port, shift_in(60) => 
                           negative_inputs_13_60_port, shift_in(59) => 
                           negative_inputs_13_59_port, shift_in(58) => 
                           negative_inputs_13_58_port, shift_in(57) => 
                           negative_inputs_13_57_port, shift_in(56) => 
                           negative_inputs_13_56_port, shift_in(55) => 
                           negative_inputs_13_55_port, shift_in(54) => 
                           negative_inputs_13_54_port, shift_in(53) => 
                           negative_inputs_13_53_port, shift_in(52) => 
                           negative_inputs_13_52_port, shift_in(51) => 
                           negative_inputs_13_51_port, shift_in(50) => 
                           negative_inputs_13_50_port, shift_in(49) => 
                           negative_inputs_13_49_port, shift_in(48) => n144, 
                           shift_in(47) => negative_inputs_13_47_port, 
                           shift_in(46) => negative_inputs_13_46_port, 
                           shift_in(45) => negative_inputs_13_45_port, 
                           shift_in(44) => negative_inputs_13_44_port, 
                           shift_in(43) => negative_inputs_13_43_port, 
                           shift_in(42) => negative_inputs_13_42_port, 
                           shift_in(41) => negative_inputs_13_41_port, 
                           shift_in(40) => negative_inputs_13_40_port, 
                           shift_in(39) => negative_inputs_13_39_port, 
                           shift_in(38) => negative_inputs_13_38_port, 
                           shift_in(37) => negative_inputs_13_37_port, 
                           shift_in(36) => negative_inputs_13_36_port, 
                           shift_in(35) => negative_inputs_13_35_port, 
                           shift_in(34) => negative_inputs_13_34_port, 
                           shift_in(33) => negative_inputs_13_33_port, 
                           shift_in(32) => negative_inputs_13_32_port, 
                           shift_in(31) => negative_inputs_13_31_port, 
                           shift_in(30) => negative_inputs_13_30_port, 
                           shift_in(29) => negative_inputs_13_29_port, 
                           shift_in(28) => negative_inputs_13_28_port, 
                           shift_in(27) => negative_inputs_13_27_port, 
                           shift_in(26) => negative_inputs_13_26_port, 
                           shift_in(25) => negative_inputs_13_25_port, 
                           shift_in(24) => negative_inputs_13_24_port, 
                           shift_in(23) => negative_inputs_13_23_port, 
                           shift_in(22) => negative_inputs_13_22_port, 
                           shift_in(21) => negative_inputs_13_21_port, 
                           shift_in(20) => negative_inputs_13_20_port, 
                           shift_in(19) => negative_inputs_13_19_port, 
                           shift_in(18) => negative_inputs_13_18_port, 
                           shift_in(17) => negative_inputs_13_17_port, 
                           shift_in(16) => negative_inputs_13_16_port, 
                           shift_in(15) => negative_inputs_13_15_port, 
                           shift_in(14) => negative_inputs_13_14_port, 
                           shift_in(13) => negative_inputs_13_13_port, 
                           shift_in(12) => negative_inputs_13_12_port, 
                           shift_in(11) => negative_inputs_13_11_port, 
                           shift_in(10) => negative_inputs_13_10_port, 
                           shift_in(9) => negative_inputs_13_9_port, 
                           shift_in(8) => negative_inputs_13_8_port, 
                           shift_in(7) => negative_inputs_13_7_port, 
                           shift_in(6) => negative_inputs_13_6_port, 
                           shift_in(5) => negative_inputs_13_5_port, 
                           shift_in(4) => negative_inputs_13_4_port, 
                           shift_in(3) => negative_inputs_13_3_port, 
                           shift_in(2) => negative_inputs_13_2_port, 
                           shift_in(1) => negative_inputs_13_1_port, 
                           shift_in(0) => n9, shift_out(63) => 
                           negative_inputs_14_63_port, shift_out(62) => 
                           negative_inputs_14_62_port, shift_out(61) => 
                           negative_inputs_14_61_port, shift_out(60) => 
                           negative_inputs_14_60_port, shift_out(59) => 
                           negative_inputs_14_59_port, shift_out(58) => 
                           negative_inputs_14_58_port, shift_out(57) => 
                           negative_inputs_14_57_port, shift_out(56) => 
                           negative_inputs_14_56_port, shift_out(55) => 
                           negative_inputs_14_55_port, shift_out(54) => 
                           negative_inputs_14_54_port, shift_out(53) => 
                           negative_inputs_14_53_port, shift_out(52) => 
                           negative_inputs_14_52_port, shift_out(51) => 
                           negative_inputs_14_51_port, shift_out(50) => 
                           negative_inputs_14_50_port, shift_out(49) => 
                           negative_inputs_14_49_port, shift_out(48) => 
                           negative_inputs_14_48_port, shift_out(47) => 
                           negative_inputs_14_47_port, shift_out(46) => 
                           negative_inputs_14_46_port, shift_out(45) => 
                           negative_inputs_14_45_port, shift_out(44) => 
                           negative_inputs_14_44_port, shift_out(43) => 
                           negative_inputs_14_43_port, shift_out(42) => 
                           negative_inputs_14_42_port, shift_out(41) => 
                           negative_inputs_14_41_port, shift_out(40) => 
                           negative_inputs_14_40_port, shift_out(39) => 
                           negative_inputs_14_39_port, shift_out(38) => 
                           negative_inputs_14_38_port, shift_out(37) => 
                           negative_inputs_14_37_port, shift_out(36) => 
                           negative_inputs_14_36_port, shift_out(35) => 
                           negative_inputs_14_35_port, shift_out(34) => 
                           negative_inputs_14_34_port, shift_out(33) => 
                           negative_inputs_14_33_port, shift_out(32) => 
                           negative_inputs_14_32_port, shift_out(31) => 
                           negative_inputs_14_31_port, shift_out(30) => 
                           negative_inputs_14_30_port, shift_out(29) => 
                           negative_inputs_14_29_port, shift_out(28) => 
                           negative_inputs_14_28_port, shift_out(27) => 
                           negative_inputs_14_27_port, shift_out(26) => 
                           negative_inputs_14_26_port, shift_out(25) => 
                           negative_inputs_14_25_port, shift_out(24) => 
                           negative_inputs_14_24_port, shift_out(23) => 
                           negative_inputs_14_23_port, shift_out(22) => 
                           negative_inputs_14_22_port, shift_out(21) => 
                           negative_inputs_14_21_port, shift_out(20) => 
                           negative_inputs_14_20_port, shift_out(19) => 
                           negative_inputs_14_19_port, shift_out(18) => 
                           negative_inputs_14_18_port, shift_out(17) => 
                           negative_inputs_14_17_port, shift_out(16) => 
                           negative_inputs_14_16_port, shift_out(15) => 
                           negative_inputs_14_15_port, shift_out(14) => 
                           negative_inputs_14_14_port, shift_out(13) => 
                           negative_inputs_14_13_port, shift_out(12) => 
                           negative_inputs_14_12_port, shift_out(11) => 
                           negative_inputs_14_11_port, shift_out(10) => 
                           negative_inputs_14_10_port, shift_out(9) => 
                           negative_inputs_14_9_port, shift_out(8) => 
                           negative_inputs_14_8_port, shift_out(7) => 
                           negative_inputs_14_7_port, shift_out(6) => 
                           negative_inputs_14_6_port, shift_out(5) => 
                           negative_inputs_14_5_port, shift_out(4) => 
                           negative_inputs_14_4_port, shift_out(3) => 
                           negative_inputs_14_3_port, shift_out(2) => 
                           negative_inputs_14_2_port, shift_out(1) => 
                           negative_inputs_14_1_port, shift_out(0) => n_1109);
   shifted_neg_15 : leftshifter_NbitShifter64_17 port map( shift_in(63) => 
                           negative_inputs_14_63_port, shift_in(62) => 
                           negative_inputs_14_62_port, shift_in(61) => 
                           negative_inputs_14_61_port, shift_in(60) => 
                           negative_inputs_14_60_port, shift_in(59) => 
                           negative_inputs_14_59_port, shift_in(58) => 
                           negative_inputs_14_58_port, shift_in(57) => 
                           negative_inputs_14_57_port, shift_in(56) => 
                           negative_inputs_14_56_port, shift_in(55) => 
                           negative_inputs_14_55_port, shift_in(54) => 
                           negative_inputs_14_54_port, shift_in(53) => 
                           negative_inputs_14_53_port, shift_in(52) => 
                           negative_inputs_14_52_port, shift_in(51) => 
                           negative_inputs_14_51_port, shift_in(50) => 
                           negative_inputs_14_50_port, shift_in(49) => 
                           negative_inputs_14_49_port, shift_in(48) => n142, 
                           shift_in(47) => negative_inputs_14_47_port, 
                           shift_in(46) => negative_inputs_14_46_port, 
                           shift_in(45) => negative_inputs_14_45_port, 
                           shift_in(44) => negative_inputs_14_44_port, 
                           shift_in(43) => negative_inputs_14_43_port, 
                           shift_in(42) => negative_inputs_14_42_port, 
                           shift_in(41) => negative_inputs_14_41_port, 
                           shift_in(40) => negative_inputs_14_40_port, 
                           shift_in(39) => negative_inputs_14_39_port, 
                           shift_in(38) => negative_inputs_14_38_port, 
                           shift_in(37) => negative_inputs_14_37_port, 
                           shift_in(36) => negative_inputs_14_36_port, 
                           shift_in(35) => negative_inputs_14_35_port, 
                           shift_in(34) => negative_inputs_14_34_port, 
                           shift_in(33) => negative_inputs_14_33_port, 
                           shift_in(32) => negative_inputs_14_32_port, 
                           shift_in(31) => negative_inputs_14_31_port, 
                           shift_in(30) => negative_inputs_14_30_port, 
                           shift_in(29) => negative_inputs_14_29_port, 
                           shift_in(28) => negative_inputs_14_28_port, 
                           shift_in(27) => negative_inputs_14_27_port, 
                           shift_in(26) => negative_inputs_14_26_port, 
                           shift_in(25) => negative_inputs_14_25_port, 
                           shift_in(24) => negative_inputs_14_24_port, 
                           shift_in(23) => negative_inputs_14_23_port, 
                           shift_in(22) => negative_inputs_14_22_port, 
                           shift_in(21) => negative_inputs_14_21_port, 
                           shift_in(20) => negative_inputs_14_20_port, 
                           shift_in(19) => negative_inputs_14_19_port, 
                           shift_in(18) => negative_inputs_14_18_port, 
                           shift_in(17) => negative_inputs_14_17_port, 
                           shift_in(16) => negative_inputs_14_16_port, 
                           shift_in(15) => negative_inputs_14_15_port, 
                           shift_in(14) => negative_inputs_14_14_port, 
                           shift_in(13) => negative_inputs_14_13_port, 
                           shift_in(12) => negative_inputs_14_12_port, 
                           shift_in(11) => negative_inputs_14_11_port, 
                           shift_in(10) => negative_inputs_14_10_port, 
                           shift_in(9) => negative_inputs_14_9_port, 
                           shift_in(8) => negative_inputs_14_8_port, 
                           shift_in(7) => negative_inputs_14_7_port, 
                           shift_in(6) => negative_inputs_14_6_port, 
                           shift_in(5) => negative_inputs_14_5_port, 
                           shift_in(4) => negative_inputs_14_4_port, 
                           shift_in(3) => negative_inputs_14_3_port, 
                           shift_in(2) => negative_inputs_14_2_port, 
                           shift_in(1) => negative_inputs_14_1_port, 
                           shift_in(0) => n9, shift_out(63) => 
                           negative_inputs_15_63_port, shift_out(62) => 
                           negative_inputs_15_62_port, shift_out(61) => 
                           negative_inputs_15_61_port, shift_out(60) => 
                           negative_inputs_15_60_port, shift_out(59) => 
                           negative_inputs_15_59_port, shift_out(58) => 
                           negative_inputs_15_58_port, shift_out(57) => 
                           negative_inputs_15_57_port, shift_out(56) => 
                           negative_inputs_15_56_port, shift_out(55) => 
                           negative_inputs_15_55_port, shift_out(54) => 
                           negative_inputs_15_54_port, shift_out(53) => 
                           negative_inputs_15_53_port, shift_out(52) => 
                           negative_inputs_15_52_port, shift_out(51) => 
                           negative_inputs_15_51_port, shift_out(50) => 
                           negative_inputs_15_50_port, shift_out(49) => 
                           negative_inputs_15_49_port, shift_out(48) => 
                           negative_inputs_15_48_port, shift_out(47) => 
                           negative_inputs_15_47_port, shift_out(46) => 
                           negative_inputs_15_46_port, shift_out(45) => 
                           negative_inputs_15_45_port, shift_out(44) => 
                           negative_inputs_15_44_port, shift_out(43) => 
                           negative_inputs_15_43_port, shift_out(42) => 
                           negative_inputs_15_42_port, shift_out(41) => 
                           negative_inputs_15_41_port, shift_out(40) => 
                           negative_inputs_15_40_port, shift_out(39) => 
                           negative_inputs_15_39_port, shift_out(38) => 
                           negative_inputs_15_38_port, shift_out(37) => 
                           negative_inputs_15_37_port, shift_out(36) => 
                           negative_inputs_15_36_port, shift_out(35) => 
                           negative_inputs_15_35_port, shift_out(34) => 
                           negative_inputs_15_34_port, shift_out(33) => 
                           negative_inputs_15_33_port, shift_out(32) => 
                           negative_inputs_15_32_port, shift_out(31) => 
                           negative_inputs_15_31_port, shift_out(30) => 
                           negative_inputs_15_30_port, shift_out(29) => 
                           negative_inputs_15_29_port, shift_out(28) => 
                           negative_inputs_15_28_port, shift_out(27) => 
                           negative_inputs_15_27_port, shift_out(26) => 
                           negative_inputs_15_26_port, shift_out(25) => 
                           negative_inputs_15_25_port, shift_out(24) => 
                           negative_inputs_15_24_port, shift_out(23) => 
                           negative_inputs_15_23_port, shift_out(22) => 
                           negative_inputs_15_22_port, shift_out(21) => 
                           negative_inputs_15_21_port, shift_out(20) => 
                           negative_inputs_15_20_port, shift_out(19) => 
                           negative_inputs_15_19_port, shift_out(18) => 
                           negative_inputs_15_18_port, shift_out(17) => 
                           negative_inputs_15_17_port, shift_out(16) => 
                           negative_inputs_15_16_port, shift_out(15) => 
                           negative_inputs_15_15_port, shift_out(14) => 
                           negative_inputs_15_14_port, shift_out(13) => 
                           negative_inputs_15_13_port, shift_out(12) => 
                           negative_inputs_15_12_port, shift_out(11) => 
                           negative_inputs_15_11_port, shift_out(10) => 
                           negative_inputs_15_10_port, shift_out(9) => 
                           negative_inputs_15_9_port, shift_out(8) => 
                           negative_inputs_15_8_port, shift_out(7) => 
                           negative_inputs_15_7_port, shift_out(6) => 
                           negative_inputs_15_6_port, shift_out(5) => 
                           negative_inputs_15_5_port, shift_out(4) => 
                           negative_inputs_15_4_port, shift_out(3) => 
                           negative_inputs_15_3_port, shift_out(2) => 
                           negative_inputs_15_2_port, shift_out(1) => 
                           negative_inputs_15_1_port, shift_out(0) => n_1110);
   shifted_neg_16 : leftshifter_NbitShifter64_16 port map( shift_in(63) => 
                           negative_inputs_15_63_port, shift_in(62) => 
                           negative_inputs_15_62_port, shift_in(61) => 
                           negative_inputs_15_61_port, shift_in(60) => 
                           negative_inputs_15_60_port, shift_in(59) => 
                           negative_inputs_15_59_port, shift_in(58) => 
                           negative_inputs_15_58_port, shift_in(57) => 
                           negative_inputs_15_57_port, shift_in(56) => 
                           negative_inputs_15_56_port, shift_in(55) => 
                           negative_inputs_15_55_port, shift_in(54) => 
                           negative_inputs_15_54_port, shift_in(53) => 
                           negative_inputs_15_53_port, shift_in(52) => 
                           negative_inputs_15_52_port, shift_in(51) => 
                           negative_inputs_15_51_port, shift_in(50) => 
                           negative_inputs_15_50_port, shift_in(49) => 
                           negative_inputs_15_49_port, shift_in(48) => n140, 
                           shift_in(47) => negative_inputs_15_47_port, 
                           shift_in(46) => negative_inputs_15_46_port, 
                           shift_in(45) => negative_inputs_15_45_port, 
                           shift_in(44) => negative_inputs_15_44_port, 
                           shift_in(43) => negative_inputs_15_43_port, 
                           shift_in(42) => negative_inputs_15_42_port, 
                           shift_in(41) => negative_inputs_15_41_port, 
                           shift_in(40) => negative_inputs_15_40_port, 
                           shift_in(39) => negative_inputs_15_39_port, 
                           shift_in(38) => negative_inputs_15_38_port, 
                           shift_in(37) => negative_inputs_15_37_port, 
                           shift_in(36) => negative_inputs_15_36_port, 
                           shift_in(35) => negative_inputs_15_35_port, 
                           shift_in(34) => negative_inputs_15_34_port, 
                           shift_in(33) => negative_inputs_15_33_port, 
                           shift_in(32) => negative_inputs_15_32_port, 
                           shift_in(31) => negative_inputs_15_31_port, 
                           shift_in(30) => negative_inputs_15_30_port, 
                           shift_in(29) => negative_inputs_15_29_port, 
                           shift_in(28) => negative_inputs_15_28_port, 
                           shift_in(27) => negative_inputs_15_27_port, 
                           shift_in(26) => negative_inputs_15_26_port, 
                           shift_in(25) => negative_inputs_15_25_port, 
                           shift_in(24) => negative_inputs_15_24_port, 
                           shift_in(23) => negative_inputs_15_23_port, 
                           shift_in(22) => negative_inputs_15_22_port, 
                           shift_in(21) => negative_inputs_15_21_port, 
                           shift_in(20) => negative_inputs_15_20_port, 
                           shift_in(19) => negative_inputs_15_19_port, 
                           shift_in(18) => negative_inputs_15_18_port, 
                           shift_in(17) => negative_inputs_15_17_port, 
                           shift_in(16) => negative_inputs_15_16_port, 
                           shift_in(15) => negative_inputs_15_15_port, 
                           shift_in(14) => negative_inputs_15_14_port, 
                           shift_in(13) => negative_inputs_15_13_port, 
                           shift_in(12) => negative_inputs_15_12_port, 
                           shift_in(11) => negative_inputs_15_11_port, 
                           shift_in(10) => negative_inputs_15_10_port, 
                           shift_in(9) => negative_inputs_15_9_port, 
                           shift_in(8) => negative_inputs_15_8_port, 
                           shift_in(7) => negative_inputs_15_7_port, 
                           shift_in(6) => negative_inputs_15_6_port, 
                           shift_in(5) => negative_inputs_15_5_port, 
                           shift_in(4) => negative_inputs_15_4_port, 
                           shift_in(3) => negative_inputs_15_3_port, 
                           shift_in(2) => negative_inputs_15_2_port, 
                           shift_in(1) => negative_inputs_15_1_port, 
                           shift_in(0) => n9, shift_out(63) => 
                           negative_inputs_16_63_port, shift_out(62) => 
                           negative_inputs_16_62_port, shift_out(61) => 
                           negative_inputs_16_61_port, shift_out(60) => 
                           negative_inputs_16_60_port, shift_out(59) => 
                           negative_inputs_16_59_port, shift_out(58) => 
                           negative_inputs_16_58_port, shift_out(57) => 
                           negative_inputs_16_57_port, shift_out(56) => 
                           negative_inputs_16_56_port, shift_out(55) => 
                           negative_inputs_16_55_port, shift_out(54) => 
                           negative_inputs_16_54_port, shift_out(53) => 
                           negative_inputs_16_53_port, shift_out(52) => 
                           negative_inputs_16_52_port, shift_out(51) => 
                           negative_inputs_16_51_port, shift_out(50) => 
                           negative_inputs_16_50_port, shift_out(49) => 
                           negative_inputs_16_49_port, shift_out(48) => 
                           negative_inputs_16_48_port, shift_out(47) => 
                           negative_inputs_16_47_port, shift_out(46) => 
                           negative_inputs_16_46_port, shift_out(45) => 
                           negative_inputs_16_45_port, shift_out(44) => 
                           negative_inputs_16_44_port, shift_out(43) => 
                           negative_inputs_16_43_port, shift_out(42) => 
                           negative_inputs_16_42_port, shift_out(41) => 
                           negative_inputs_16_41_port, shift_out(40) => 
                           negative_inputs_16_40_port, shift_out(39) => 
                           negative_inputs_16_39_port, shift_out(38) => 
                           negative_inputs_16_38_port, shift_out(37) => 
                           negative_inputs_16_37_port, shift_out(36) => 
                           negative_inputs_16_36_port, shift_out(35) => 
                           negative_inputs_16_35_port, shift_out(34) => 
                           negative_inputs_16_34_port, shift_out(33) => 
                           negative_inputs_16_33_port, shift_out(32) => 
                           negative_inputs_16_32_port, shift_out(31) => 
                           negative_inputs_16_31_port, shift_out(30) => 
                           negative_inputs_16_30_port, shift_out(29) => 
                           negative_inputs_16_29_port, shift_out(28) => 
                           negative_inputs_16_28_port, shift_out(27) => 
                           negative_inputs_16_27_port, shift_out(26) => 
                           negative_inputs_16_26_port, shift_out(25) => 
                           negative_inputs_16_25_port, shift_out(24) => 
                           negative_inputs_16_24_port, shift_out(23) => 
                           negative_inputs_16_23_port, shift_out(22) => 
                           negative_inputs_16_22_port, shift_out(21) => 
                           negative_inputs_16_21_port, shift_out(20) => 
                           negative_inputs_16_20_port, shift_out(19) => 
                           negative_inputs_16_19_port, shift_out(18) => 
                           negative_inputs_16_18_port, shift_out(17) => 
                           negative_inputs_16_17_port, shift_out(16) => 
                           negative_inputs_16_16_port, shift_out(15) => 
                           negative_inputs_16_15_port, shift_out(14) => 
                           negative_inputs_16_14_port, shift_out(13) => 
                           negative_inputs_16_13_port, shift_out(12) => 
                           negative_inputs_16_12_port, shift_out(11) => 
                           negative_inputs_16_11_port, shift_out(10) => 
                           negative_inputs_16_10_port, shift_out(9) => 
                           negative_inputs_16_9_port, shift_out(8) => 
                           negative_inputs_16_8_port, shift_out(7) => 
                           negative_inputs_16_7_port, shift_out(6) => 
                           negative_inputs_16_6_port, shift_out(5) => 
                           negative_inputs_16_5_port, shift_out(4) => 
                           negative_inputs_16_4_port, shift_out(3) => 
                           negative_inputs_16_3_port, shift_out(2) => 
                           negative_inputs_16_2_port, shift_out(1) => 
                           negative_inputs_16_1_port, shift_out(0) => n_1111);
   shifted_neg_17 : leftshifter_NbitShifter64_15 port map( shift_in(63) => 
                           negative_inputs_16_63_port, shift_in(62) => 
                           negative_inputs_16_62_port, shift_in(61) => 
                           negative_inputs_16_61_port, shift_in(60) => 
                           negative_inputs_16_60_port, shift_in(59) => 
                           negative_inputs_16_59_port, shift_in(58) => 
                           negative_inputs_16_58_port, shift_in(57) => 
                           negative_inputs_16_57_port, shift_in(56) => 
                           negative_inputs_16_56_port, shift_in(55) => 
                           negative_inputs_16_55_port, shift_in(54) => 
                           negative_inputs_16_54_port, shift_in(53) => 
                           negative_inputs_16_53_port, shift_in(52) => 
                           negative_inputs_16_52_port, shift_in(51) => 
                           negative_inputs_16_51_port, shift_in(50) => 
                           negative_inputs_16_50_port, shift_in(49) => 
                           negative_inputs_16_49_port, shift_in(48) => n138, 
                           shift_in(47) => n136, shift_in(46) => n134, 
                           shift_in(45) => n132, shift_in(44) => n130, 
                           shift_in(43) => n128, shift_in(42) => n126, 
                           shift_in(41) => n124, shift_in(40) => n122, 
                           shift_in(39) => n120, shift_in(38) => n118, 
                           shift_in(37) => n116, shift_in(36) => n114, 
                           shift_in(35) => n112, shift_in(34) => n110, 
                           shift_in(33) => n108, shift_in(32) => n106, 
                           shift_in(31) => n104, shift_in(30) => n102, 
                           shift_in(29) => n100, shift_in(28) => n98, 
                           shift_in(27) => n96, shift_in(26) => n94, 
                           shift_in(25) => n92, shift_in(24) => n90, 
                           shift_in(23) => n88, shift_in(22) => n86, 
                           shift_in(21) => n84, shift_in(20) => n82, 
                           shift_in(19) => n80, shift_in(18) => n78, 
                           shift_in(17) => n76, shift_in(16) => n74, 
                           shift_in(15) => negative_inputs_16_15_port, 
                           shift_in(14) => negative_inputs_16_14_port, 
                           shift_in(13) => negative_inputs_16_13_port, 
                           shift_in(12) => negative_inputs_16_12_port, 
                           shift_in(11) => negative_inputs_16_11_port, 
                           shift_in(10) => negative_inputs_16_10_port, 
                           shift_in(9) => negative_inputs_16_9_port, 
                           shift_in(8) => negative_inputs_16_8_port, 
                           shift_in(7) => negative_inputs_16_7_port, 
                           shift_in(6) => negative_inputs_16_6_port, 
                           shift_in(5) => negative_inputs_16_5_port, 
                           shift_in(4) => negative_inputs_16_4_port, 
                           shift_in(3) => negative_inputs_16_3_port, 
                           shift_in(2) => negative_inputs_16_2_port, 
                           shift_in(1) => negative_inputs_16_1_port, 
                           shift_in(0) => n9, shift_out(63) => 
                           negative_inputs_17_63_port, shift_out(62) => 
                           negative_inputs_17_62_port, shift_out(61) => 
                           negative_inputs_17_61_port, shift_out(60) => 
                           negative_inputs_17_60_port, shift_out(59) => 
                           negative_inputs_17_59_port, shift_out(58) => 
                           negative_inputs_17_58_port, shift_out(57) => 
                           negative_inputs_17_57_port, shift_out(56) => 
                           negative_inputs_17_56_port, shift_out(55) => 
                           negative_inputs_17_55_port, shift_out(54) => 
                           negative_inputs_17_54_port, shift_out(53) => 
                           negative_inputs_17_53_port, shift_out(52) => 
                           negative_inputs_17_52_port, shift_out(51) => 
                           negative_inputs_17_51_port, shift_out(50) => 
                           negative_inputs_17_50_port, shift_out(49) => 
                           negative_inputs_17_49_port, shift_out(48) => 
                           negative_inputs_17_48_port, shift_out(47) => 
                           negative_inputs_17_47_port, shift_out(46) => 
                           negative_inputs_17_46_port, shift_out(45) => 
                           negative_inputs_17_45_port, shift_out(44) => 
                           negative_inputs_17_44_port, shift_out(43) => 
                           negative_inputs_17_43_port, shift_out(42) => 
                           negative_inputs_17_42_port, shift_out(41) => 
                           negative_inputs_17_41_port, shift_out(40) => 
                           negative_inputs_17_40_port, shift_out(39) => 
                           negative_inputs_17_39_port, shift_out(38) => 
                           negative_inputs_17_38_port, shift_out(37) => 
                           negative_inputs_17_37_port, shift_out(36) => 
                           negative_inputs_17_36_port, shift_out(35) => 
                           negative_inputs_17_35_port, shift_out(34) => 
                           negative_inputs_17_34_port, shift_out(33) => 
                           negative_inputs_17_33_port, shift_out(32) => 
                           negative_inputs_17_32_port, shift_out(31) => 
                           negative_inputs_17_31_port, shift_out(30) => 
                           negative_inputs_17_30_port, shift_out(29) => 
                           negative_inputs_17_29_port, shift_out(28) => 
                           negative_inputs_17_28_port, shift_out(27) => 
                           negative_inputs_17_27_port, shift_out(26) => 
                           negative_inputs_17_26_port, shift_out(25) => 
                           negative_inputs_17_25_port, shift_out(24) => 
                           negative_inputs_17_24_port, shift_out(23) => 
                           negative_inputs_17_23_port, shift_out(22) => 
                           negative_inputs_17_22_port, shift_out(21) => 
                           negative_inputs_17_21_port, shift_out(20) => 
                           negative_inputs_17_20_port, shift_out(19) => 
                           negative_inputs_17_19_port, shift_out(18) => 
                           negative_inputs_17_18_port, shift_out(17) => 
                           negative_inputs_17_17_port, shift_out(16) => 
                           negative_inputs_17_16_port, shift_out(15) => 
                           negative_inputs_17_15_port, shift_out(14) => 
                           negative_inputs_17_14_port, shift_out(13) => 
                           negative_inputs_17_13_port, shift_out(12) => 
                           negative_inputs_17_12_port, shift_out(11) => 
                           negative_inputs_17_11_port, shift_out(10) => 
                           negative_inputs_17_10_port, shift_out(9) => 
                           negative_inputs_17_9_port, shift_out(8) => 
                           negative_inputs_17_8_port, shift_out(7) => 
                           negative_inputs_17_7_port, shift_out(6) => 
                           negative_inputs_17_6_port, shift_out(5) => 
                           negative_inputs_17_5_port, shift_out(4) => 
                           negative_inputs_17_4_port, shift_out(3) => 
                           negative_inputs_17_3_port, shift_out(2) => 
                           negative_inputs_17_2_port, shift_out(1) => 
                           negative_inputs_17_1_port, shift_out(0) => n_1112);
   shifted_neg_18 : leftshifter_NbitShifter64_14 port map( shift_in(63) => 
                           negative_inputs_17_63_port, shift_in(62) => 
                           negative_inputs_17_62_port, shift_in(61) => 
                           negative_inputs_17_61_port, shift_in(60) => 
                           negative_inputs_17_60_port, shift_in(59) => 
                           negative_inputs_17_59_port, shift_in(58) => 
                           negative_inputs_17_58_port, shift_in(57) => 
                           negative_inputs_17_57_port, shift_in(56) => 
                           negative_inputs_17_56_port, shift_in(55) => 
                           negative_inputs_17_55_port, shift_in(54) => 
                           negative_inputs_17_54_port, shift_in(53) => 
                           negative_inputs_17_53_port, shift_in(52) => 
                           negative_inputs_17_52_port, shift_in(51) => 
                           negative_inputs_17_51_port, shift_in(50) => 
                           negative_inputs_17_50_port, shift_in(49) => 
                           negative_inputs_17_49_port, shift_in(48) => 
                           negative_inputs_17_48_port, shift_in(47) => 
                           negative_inputs_17_47_port, shift_in(46) => 
                           negative_inputs_17_46_port, shift_in(45) => 
                           negative_inputs_17_45_port, shift_in(44) => 
                           negative_inputs_17_44_port, shift_in(43) => 
                           negative_inputs_17_43_port, shift_in(42) => 
                           negative_inputs_17_42_port, shift_in(41) => 
                           negative_inputs_17_41_port, shift_in(40) => 
                           negative_inputs_17_40_port, shift_in(39) => 
                           negative_inputs_17_39_port, shift_in(38) => 
                           negative_inputs_17_38_port, shift_in(37) => 
                           negative_inputs_17_37_port, shift_in(36) => 
                           negative_inputs_17_36_port, shift_in(35) => 
                           negative_inputs_17_35_port, shift_in(34) => 
                           negative_inputs_17_34_port, shift_in(33) => 
                           negative_inputs_17_33_port, shift_in(32) => 
                           negative_inputs_17_32_port, shift_in(31) => 
                           negative_inputs_17_31_port, shift_in(30) => 
                           negative_inputs_17_30_port, shift_in(29) => 
                           negative_inputs_17_29_port, shift_in(28) => 
                           negative_inputs_17_28_port, shift_in(27) => 
                           negative_inputs_17_27_port, shift_in(26) => 
                           negative_inputs_17_26_port, shift_in(25) => 
                           negative_inputs_17_25_port, shift_in(24) => 
                           negative_inputs_17_24_port, shift_in(23) => 
                           negative_inputs_17_23_port, shift_in(22) => 
                           negative_inputs_17_22_port, shift_in(21) => 
                           negative_inputs_17_21_port, shift_in(20) => 
                           negative_inputs_17_20_port, shift_in(19) => 
                           negative_inputs_17_19_port, shift_in(18) => 
                           negative_inputs_17_18_port, shift_in(17) => 
                           negative_inputs_17_17_port, shift_in(16) => 
                           negative_inputs_17_16_port, shift_in(15) => 
                           negative_inputs_17_15_port, shift_in(14) => 
                           negative_inputs_17_14_port, shift_in(13) => 
                           negative_inputs_17_13_port, shift_in(12) => 
                           negative_inputs_17_12_port, shift_in(11) => 
                           negative_inputs_17_11_port, shift_in(10) => 
                           negative_inputs_17_10_port, shift_in(9) => 
                           negative_inputs_17_9_port, shift_in(8) => 
                           negative_inputs_17_8_port, shift_in(7) => 
                           negative_inputs_17_7_port, shift_in(6) => 
                           negative_inputs_17_6_port, shift_in(5) => 
                           negative_inputs_17_5_port, shift_in(4) => 
                           negative_inputs_17_4_port, shift_in(3) => 
                           negative_inputs_17_3_port, shift_in(2) => 
                           negative_inputs_17_2_port, shift_in(1) => 
                           negative_inputs_17_1_port, shift_in(0) => n9, 
                           shift_out(63) => negative_inputs_18_63_port, 
                           shift_out(62) => negative_inputs_18_62_port, 
                           shift_out(61) => negative_inputs_18_61_port, 
                           shift_out(60) => negative_inputs_18_60_port, 
                           shift_out(59) => negative_inputs_18_59_port, 
                           shift_out(58) => negative_inputs_18_58_port, 
                           shift_out(57) => negative_inputs_18_57_port, 
                           shift_out(56) => negative_inputs_18_56_port, 
                           shift_out(55) => negative_inputs_18_55_port, 
                           shift_out(54) => negative_inputs_18_54_port, 
                           shift_out(53) => negative_inputs_18_53_port, 
                           shift_out(52) => negative_inputs_18_52_port, 
                           shift_out(51) => negative_inputs_18_51_port, 
                           shift_out(50) => negative_inputs_18_50_port, 
                           shift_out(49) => negative_inputs_18_49_port, 
                           shift_out(48) => negative_inputs_18_48_port, 
                           shift_out(47) => negative_inputs_18_47_port, 
                           shift_out(46) => negative_inputs_18_46_port, 
                           shift_out(45) => negative_inputs_18_45_port, 
                           shift_out(44) => negative_inputs_18_44_port, 
                           shift_out(43) => negative_inputs_18_43_port, 
                           shift_out(42) => negative_inputs_18_42_port, 
                           shift_out(41) => negative_inputs_18_41_port, 
                           shift_out(40) => negative_inputs_18_40_port, 
                           shift_out(39) => negative_inputs_18_39_port, 
                           shift_out(38) => negative_inputs_18_38_port, 
                           shift_out(37) => negative_inputs_18_37_port, 
                           shift_out(36) => negative_inputs_18_36_port, 
                           shift_out(35) => negative_inputs_18_35_port, 
                           shift_out(34) => negative_inputs_18_34_port, 
                           shift_out(33) => negative_inputs_18_33_port, 
                           shift_out(32) => negative_inputs_18_32_port, 
                           shift_out(31) => negative_inputs_18_31_port, 
                           shift_out(30) => negative_inputs_18_30_port, 
                           shift_out(29) => negative_inputs_18_29_port, 
                           shift_out(28) => negative_inputs_18_28_port, 
                           shift_out(27) => negative_inputs_18_27_port, 
                           shift_out(26) => negative_inputs_18_26_port, 
                           shift_out(25) => negative_inputs_18_25_port, 
                           shift_out(24) => negative_inputs_18_24_port, 
                           shift_out(23) => negative_inputs_18_23_port, 
                           shift_out(22) => negative_inputs_18_22_port, 
                           shift_out(21) => negative_inputs_18_21_port, 
                           shift_out(20) => negative_inputs_18_20_port, 
                           shift_out(19) => negative_inputs_18_19_port, 
                           shift_out(18) => negative_inputs_18_18_port, 
                           shift_out(17) => negative_inputs_18_17_port, 
                           shift_out(16) => negative_inputs_18_16_port, 
                           shift_out(15) => negative_inputs_18_15_port, 
                           shift_out(14) => negative_inputs_18_14_port, 
                           shift_out(13) => negative_inputs_18_13_port, 
                           shift_out(12) => negative_inputs_18_12_port, 
                           shift_out(11) => negative_inputs_18_11_port, 
                           shift_out(10) => negative_inputs_18_10_port, 
                           shift_out(9) => negative_inputs_18_9_port, 
                           shift_out(8) => negative_inputs_18_8_port, 
                           shift_out(7) => negative_inputs_18_7_port, 
                           shift_out(6) => negative_inputs_18_6_port, 
                           shift_out(5) => negative_inputs_18_5_port, 
                           shift_out(4) => negative_inputs_18_4_port, 
                           shift_out(3) => negative_inputs_18_3_port, 
                           shift_out(2) => negative_inputs_18_2_port, 
                           shift_out(1) => negative_inputs_18_1_port, 
                           shift_out(0) => n_1113);
   shifted_neg_19 : leftshifter_NbitShifter64_13 port map( shift_in(63) => 
                           negative_inputs_18_63_port, shift_in(62) => 
                           negative_inputs_18_62_port, shift_in(61) => 
                           negative_inputs_18_61_port, shift_in(60) => 
                           negative_inputs_18_60_port, shift_in(59) => 
                           negative_inputs_18_59_port, shift_in(58) => 
                           negative_inputs_18_58_port, shift_in(57) => 
                           negative_inputs_18_57_port, shift_in(56) => 
                           negative_inputs_18_56_port, shift_in(55) => 
                           negative_inputs_18_55_port, shift_in(54) => 
                           negative_inputs_18_54_port, shift_in(53) => 
                           negative_inputs_18_53_port, shift_in(52) => 
                           negative_inputs_18_52_port, shift_in(51) => 
                           negative_inputs_18_51_port, shift_in(50) => 
                           negative_inputs_18_50_port, shift_in(49) => 
                           negative_inputs_18_49_port, shift_in(48) => 
                           negative_inputs_18_48_port, shift_in(47) => 
                           negative_inputs_18_47_port, shift_in(46) => 
                           negative_inputs_18_46_port, shift_in(45) => 
                           negative_inputs_18_45_port, shift_in(44) => 
                           negative_inputs_18_44_port, shift_in(43) => 
                           negative_inputs_18_43_port, shift_in(42) => 
                           negative_inputs_18_42_port, shift_in(41) => 
                           negative_inputs_18_41_port, shift_in(40) => 
                           negative_inputs_18_40_port, shift_in(39) => 
                           negative_inputs_18_39_port, shift_in(38) => 
                           negative_inputs_18_38_port, shift_in(37) => 
                           negative_inputs_18_37_port, shift_in(36) => 
                           negative_inputs_18_36_port, shift_in(35) => 
                           negative_inputs_18_35_port, shift_in(34) => 
                           negative_inputs_18_34_port, shift_in(33) => 
                           negative_inputs_18_33_port, shift_in(32) => 
                           negative_inputs_18_32_port, shift_in(31) => 
                           negative_inputs_18_31_port, shift_in(30) => 
                           negative_inputs_18_30_port, shift_in(29) => 
                           negative_inputs_18_29_port, shift_in(28) => 
                           negative_inputs_18_28_port, shift_in(27) => 
                           negative_inputs_18_27_port, shift_in(26) => 
                           negative_inputs_18_26_port, shift_in(25) => 
                           negative_inputs_18_25_port, shift_in(24) => 
                           negative_inputs_18_24_port, shift_in(23) => 
                           negative_inputs_18_23_port, shift_in(22) => 
                           negative_inputs_18_22_port, shift_in(21) => 
                           negative_inputs_18_21_port, shift_in(20) => 
                           negative_inputs_18_20_port, shift_in(19) => 
                           negative_inputs_18_19_port, shift_in(18) => 
                           negative_inputs_18_18_port, shift_in(17) => 
                           negative_inputs_18_17_port, shift_in(16) => 
                           negative_inputs_18_16_port, shift_in(15) => 
                           negative_inputs_18_15_port, shift_in(14) => 
                           negative_inputs_18_14_port, shift_in(13) => 
                           negative_inputs_18_13_port, shift_in(12) => 
                           negative_inputs_18_12_port, shift_in(11) => 
                           negative_inputs_18_11_port, shift_in(10) => 
                           negative_inputs_18_10_port, shift_in(9) => 
                           negative_inputs_18_9_port, shift_in(8) => 
                           negative_inputs_18_8_port, shift_in(7) => 
                           negative_inputs_18_7_port, shift_in(6) => 
                           negative_inputs_18_6_port, shift_in(5) => 
                           negative_inputs_18_5_port, shift_in(4) => 
                           negative_inputs_18_4_port, shift_in(3) => 
                           negative_inputs_18_3_port, shift_in(2) => 
                           negative_inputs_18_2_port, shift_in(1) => 
                           negative_inputs_18_1_port, shift_in(0) => n9, 
                           shift_out(63) => negative_inputs_19_63_port, 
                           shift_out(62) => negative_inputs_19_62_port, 
                           shift_out(61) => negative_inputs_19_61_port, 
                           shift_out(60) => negative_inputs_19_60_port, 
                           shift_out(59) => negative_inputs_19_59_port, 
                           shift_out(58) => negative_inputs_19_58_port, 
                           shift_out(57) => negative_inputs_19_57_port, 
                           shift_out(56) => negative_inputs_19_56_port, 
                           shift_out(55) => negative_inputs_19_55_port, 
                           shift_out(54) => negative_inputs_19_54_port, 
                           shift_out(53) => negative_inputs_19_53_port, 
                           shift_out(52) => negative_inputs_19_52_port, 
                           shift_out(51) => negative_inputs_19_51_port, 
                           shift_out(50) => negative_inputs_19_50_port, 
                           shift_out(49) => negative_inputs_19_49_port, 
                           shift_out(48) => negative_inputs_19_48_port, 
                           shift_out(47) => negative_inputs_19_47_port, 
                           shift_out(46) => negative_inputs_19_46_port, 
                           shift_out(45) => negative_inputs_19_45_port, 
                           shift_out(44) => negative_inputs_19_44_port, 
                           shift_out(43) => negative_inputs_19_43_port, 
                           shift_out(42) => negative_inputs_19_42_port, 
                           shift_out(41) => negative_inputs_19_41_port, 
                           shift_out(40) => negative_inputs_19_40_port, 
                           shift_out(39) => negative_inputs_19_39_port, 
                           shift_out(38) => negative_inputs_19_38_port, 
                           shift_out(37) => negative_inputs_19_37_port, 
                           shift_out(36) => negative_inputs_19_36_port, 
                           shift_out(35) => negative_inputs_19_35_port, 
                           shift_out(34) => negative_inputs_19_34_port, 
                           shift_out(33) => negative_inputs_19_33_port, 
                           shift_out(32) => negative_inputs_19_32_port, 
                           shift_out(31) => negative_inputs_19_31_port, 
                           shift_out(30) => negative_inputs_19_30_port, 
                           shift_out(29) => negative_inputs_19_29_port, 
                           shift_out(28) => negative_inputs_19_28_port, 
                           shift_out(27) => negative_inputs_19_27_port, 
                           shift_out(26) => negative_inputs_19_26_port, 
                           shift_out(25) => negative_inputs_19_25_port, 
                           shift_out(24) => negative_inputs_19_24_port, 
                           shift_out(23) => negative_inputs_19_23_port, 
                           shift_out(22) => negative_inputs_19_22_port, 
                           shift_out(21) => negative_inputs_19_21_port, 
                           shift_out(20) => negative_inputs_19_20_port, 
                           shift_out(19) => negative_inputs_19_19_port, 
                           shift_out(18) => negative_inputs_19_18_port, 
                           shift_out(17) => negative_inputs_19_17_port, 
                           shift_out(16) => negative_inputs_19_16_port, 
                           shift_out(15) => negative_inputs_19_15_port, 
                           shift_out(14) => negative_inputs_19_14_port, 
                           shift_out(13) => negative_inputs_19_13_port, 
                           shift_out(12) => negative_inputs_19_12_port, 
                           shift_out(11) => negative_inputs_19_11_port, 
                           shift_out(10) => negative_inputs_19_10_port, 
                           shift_out(9) => negative_inputs_19_9_port, 
                           shift_out(8) => negative_inputs_19_8_port, 
                           shift_out(7) => negative_inputs_19_7_port, 
                           shift_out(6) => negative_inputs_19_6_port, 
                           shift_out(5) => negative_inputs_19_5_port, 
                           shift_out(4) => negative_inputs_19_4_port, 
                           shift_out(3) => negative_inputs_19_3_port, 
                           shift_out(2) => negative_inputs_19_2_port, 
                           shift_out(1) => negative_inputs_19_1_port, 
                           shift_out(0) => n_1114);
   shifted_neg_20 : leftshifter_NbitShifter64_12 port map( shift_in(63) => 
                           negative_inputs_19_63_port, shift_in(62) => 
                           negative_inputs_19_62_port, shift_in(61) => 
                           negative_inputs_19_61_port, shift_in(60) => 
                           negative_inputs_19_60_port, shift_in(59) => 
                           negative_inputs_19_59_port, shift_in(58) => 
                           negative_inputs_19_58_port, shift_in(57) => 
                           negative_inputs_19_57_port, shift_in(56) => 
                           negative_inputs_19_56_port, shift_in(55) => 
                           negative_inputs_19_55_port, shift_in(54) => 
                           negative_inputs_19_54_port, shift_in(53) => 
                           negative_inputs_19_53_port, shift_in(52) => 
                           negative_inputs_19_52_port, shift_in(51) => 
                           negative_inputs_19_51_port, shift_in(50) => 
                           negative_inputs_19_50_port, shift_in(49) => 
                           negative_inputs_19_49_port, shift_in(48) => 
                           negative_inputs_19_48_port, shift_in(47) => 
                           negative_inputs_19_47_port, shift_in(46) => 
                           negative_inputs_19_46_port, shift_in(45) => 
                           negative_inputs_19_45_port, shift_in(44) => 
                           negative_inputs_19_44_port, shift_in(43) => 
                           negative_inputs_19_43_port, shift_in(42) => 
                           negative_inputs_19_42_port, shift_in(41) => 
                           negative_inputs_19_41_port, shift_in(40) => 
                           negative_inputs_19_40_port, shift_in(39) => 
                           negative_inputs_19_39_port, shift_in(38) => 
                           negative_inputs_19_38_port, shift_in(37) => 
                           negative_inputs_19_37_port, shift_in(36) => 
                           negative_inputs_19_36_port, shift_in(35) => 
                           negative_inputs_19_35_port, shift_in(34) => 
                           negative_inputs_19_34_port, shift_in(33) => 
                           negative_inputs_19_33_port, shift_in(32) => 
                           negative_inputs_19_32_port, shift_in(31) => 
                           negative_inputs_19_31_port, shift_in(30) => 
                           negative_inputs_19_30_port, shift_in(29) => 
                           negative_inputs_19_29_port, shift_in(28) => 
                           negative_inputs_19_28_port, shift_in(27) => 
                           negative_inputs_19_27_port, shift_in(26) => 
                           negative_inputs_19_26_port, shift_in(25) => 
                           negative_inputs_19_25_port, shift_in(24) => 
                           negative_inputs_19_24_port, shift_in(23) => 
                           negative_inputs_19_23_port, shift_in(22) => 
                           negative_inputs_19_22_port, shift_in(21) => 
                           negative_inputs_19_21_port, shift_in(20) => 
                           negative_inputs_19_20_port, shift_in(19) => 
                           negative_inputs_19_19_port, shift_in(18) => 
                           negative_inputs_19_18_port, shift_in(17) => 
                           negative_inputs_19_17_port, shift_in(16) => 
                           negative_inputs_19_16_port, shift_in(15) => 
                           negative_inputs_19_15_port, shift_in(14) => 
                           negative_inputs_19_14_port, shift_in(13) => 
                           negative_inputs_19_13_port, shift_in(12) => 
                           negative_inputs_19_12_port, shift_in(11) => 
                           negative_inputs_19_11_port, shift_in(10) => 
                           negative_inputs_19_10_port, shift_in(9) => 
                           negative_inputs_19_9_port, shift_in(8) => 
                           negative_inputs_19_8_port, shift_in(7) => 
                           negative_inputs_19_7_port, shift_in(6) => 
                           negative_inputs_19_6_port, shift_in(5) => 
                           negative_inputs_19_5_port, shift_in(4) => 
                           negative_inputs_19_4_port, shift_in(3) => 
                           negative_inputs_19_3_port, shift_in(2) => 
                           negative_inputs_19_2_port, shift_in(1) => 
                           negative_inputs_19_1_port, shift_in(0) => n9, 
                           shift_out(63) => negative_inputs_20_63_port, 
                           shift_out(62) => negative_inputs_20_62_port, 
                           shift_out(61) => negative_inputs_20_61_port, 
                           shift_out(60) => negative_inputs_20_60_port, 
                           shift_out(59) => negative_inputs_20_59_port, 
                           shift_out(58) => negative_inputs_20_58_port, 
                           shift_out(57) => negative_inputs_20_57_port, 
                           shift_out(56) => negative_inputs_20_56_port, 
                           shift_out(55) => negative_inputs_20_55_port, 
                           shift_out(54) => negative_inputs_20_54_port, 
                           shift_out(53) => negative_inputs_20_53_port, 
                           shift_out(52) => negative_inputs_20_52_port, 
                           shift_out(51) => negative_inputs_20_51_port, 
                           shift_out(50) => negative_inputs_20_50_port, 
                           shift_out(49) => negative_inputs_20_49_port, 
                           shift_out(48) => negative_inputs_20_48_port, 
                           shift_out(47) => negative_inputs_20_47_port, 
                           shift_out(46) => negative_inputs_20_46_port, 
                           shift_out(45) => negative_inputs_20_45_port, 
                           shift_out(44) => negative_inputs_20_44_port, 
                           shift_out(43) => negative_inputs_20_43_port, 
                           shift_out(42) => negative_inputs_20_42_port, 
                           shift_out(41) => negative_inputs_20_41_port, 
                           shift_out(40) => negative_inputs_20_40_port, 
                           shift_out(39) => negative_inputs_20_39_port, 
                           shift_out(38) => negative_inputs_20_38_port, 
                           shift_out(37) => negative_inputs_20_37_port, 
                           shift_out(36) => negative_inputs_20_36_port, 
                           shift_out(35) => negative_inputs_20_35_port, 
                           shift_out(34) => negative_inputs_20_34_port, 
                           shift_out(33) => negative_inputs_20_33_port, 
                           shift_out(32) => negative_inputs_20_32_port, 
                           shift_out(31) => negative_inputs_20_31_port, 
                           shift_out(30) => negative_inputs_20_30_port, 
                           shift_out(29) => negative_inputs_20_29_port, 
                           shift_out(28) => negative_inputs_20_28_port, 
                           shift_out(27) => negative_inputs_20_27_port, 
                           shift_out(26) => negative_inputs_20_26_port, 
                           shift_out(25) => negative_inputs_20_25_port, 
                           shift_out(24) => negative_inputs_20_24_port, 
                           shift_out(23) => negative_inputs_20_23_port, 
                           shift_out(22) => negative_inputs_20_22_port, 
                           shift_out(21) => negative_inputs_20_21_port, 
                           shift_out(20) => negative_inputs_20_20_port, 
                           shift_out(19) => negative_inputs_20_19_port, 
                           shift_out(18) => negative_inputs_20_18_port, 
                           shift_out(17) => negative_inputs_20_17_port, 
                           shift_out(16) => negative_inputs_20_16_port, 
                           shift_out(15) => negative_inputs_20_15_port, 
                           shift_out(14) => negative_inputs_20_14_port, 
                           shift_out(13) => negative_inputs_20_13_port, 
                           shift_out(12) => negative_inputs_20_12_port, 
                           shift_out(11) => negative_inputs_20_11_port, 
                           shift_out(10) => negative_inputs_20_10_port, 
                           shift_out(9) => negative_inputs_20_9_port, 
                           shift_out(8) => negative_inputs_20_8_port, 
                           shift_out(7) => negative_inputs_20_7_port, 
                           shift_out(6) => negative_inputs_20_6_port, 
                           shift_out(5) => negative_inputs_20_5_port, 
                           shift_out(4) => negative_inputs_20_4_port, 
                           shift_out(3) => negative_inputs_20_3_port, 
                           shift_out(2) => negative_inputs_20_2_port, 
                           shift_out(1) => negative_inputs_20_1_port, 
                           shift_out(0) => n_1115);
   shifted_neg_21 : leftshifter_NbitShifter64_11 port map( shift_in(63) => 
                           negative_inputs_20_63_port, shift_in(62) => 
                           negative_inputs_20_62_port, shift_in(61) => 
                           negative_inputs_20_61_port, shift_in(60) => 
                           negative_inputs_20_60_port, shift_in(59) => 
                           negative_inputs_20_59_port, shift_in(58) => 
                           negative_inputs_20_58_port, shift_in(57) => 
                           negative_inputs_20_57_port, shift_in(56) => 
                           negative_inputs_20_56_port, shift_in(55) => 
                           negative_inputs_20_55_port, shift_in(54) => 
                           negative_inputs_20_54_port, shift_in(53) => 
                           negative_inputs_20_53_port, shift_in(52) => 
                           negative_inputs_20_52_port, shift_in(51) => 
                           negative_inputs_20_51_port, shift_in(50) => 
                           negative_inputs_20_50_port, shift_in(49) => 
                           negative_inputs_20_49_port, shift_in(48) => 
                           negative_inputs_20_48_port, shift_in(47) => 
                           negative_inputs_20_47_port, shift_in(46) => 
                           negative_inputs_20_46_port, shift_in(45) => 
                           negative_inputs_20_45_port, shift_in(44) => 
                           negative_inputs_20_44_port, shift_in(43) => 
                           negative_inputs_20_43_port, shift_in(42) => 
                           negative_inputs_20_42_port, shift_in(41) => 
                           negative_inputs_20_41_port, shift_in(40) => 
                           negative_inputs_20_40_port, shift_in(39) => 
                           negative_inputs_20_39_port, shift_in(38) => 
                           negative_inputs_20_38_port, shift_in(37) => 
                           negative_inputs_20_37_port, shift_in(36) => 
                           negative_inputs_20_36_port, shift_in(35) => 
                           negative_inputs_20_35_port, shift_in(34) => 
                           negative_inputs_20_34_port, shift_in(33) => 
                           negative_inputs_20_33_port, shift_in(32) => 
                           negative_inputs_20_32_port, shift_in(31) => 
                           negative_inputs_20_31_port, shift_in(30) => 
                           negative_inputs_20_30_port, shift_in(29) => 
                           negative_inputs_20_29_port, shift_in(28) => 
                           negative_inputs_20_28_port, shift_in(27) => 
                           negative_inputs_20_27_port, shift_in(26) => 
                           negative_inputs_20_26_port, shift_in(25) => 
                           negative_inputs_20_25_port, shift_in(24) => 
                           negative_inputs_20_24_port, shift_in(23) => 
                           negative_inputs_20_23_port, shift_in(22) => 
                           negative_inputs_20_22_port, shift_in(21) => 
                           negative_inputs_20_21_port, shift_in(20) => 
                           negative_inputs_20_20_port, shift_in(19) => 
                           negative_inputs_20_19_port, shift_in(18) => 
                           negative_inputs_20_18_port, shift_in(17) => 
                           negative_inputs_20_17_port, shift_in(16) => 
                           negative_inputs_20_16_port, shift_in(15) => 
                           negative_inputs_20_15_port, shift_in(14) => 
                           negative_inputs_20_14_port, shift_in(13) => 
                           negative_inputs_20_13_port, shift_in(12) => 
                           negative_inputs_20_12_port, shift_in(11) => 
                           negative_inputs_20_11_port, shift_in(10) => 
                           negative_inputs_20_10_port, shift_in(9) => 
                           negative_inputs_20_9_port, shift_in(8) => 
                           negative_inputs_20_8_port, shift_in(7) => 
                           negative_inputs_20_7_port, shift_in(6) => 
                           negative_inputs_20_6_port, shift_in(5) => 
                           negative_inputs_20_5_port, shift_in(4) => 
                           negative_inputs_20_4_port, shift_in(3) => 
                           negative_inputs_20_3_port, shift_in(2) => 
                           negative_inputs_20_2_port, shift_in(1) => 
                           negative_inputs_20_1_port, shift_in(0) => n9, 
                           shift_out(63) => negative_inputs_21_63_port, 
                           shift_out(62) => negative_inputs_21_62_port, 
                           shift_out(61) => negative_inputs_21_61_port, 
                           shift_out(60) => negative_inputs_21_60_port, 
                           shift_out(59) => negative_inputs_21_59_port, 
                           shift_out(58) => negative_inputs_21_58_port, 
                           shift_out(57) => negative_inputs_21_57_port, 
                           shift_out(56) => negative_inputs_21_56_port, 
                           shift_out(55) => negative_inputs_21_55_port, 
                           shift_out(54) => negative_inputs_21_54_port, 
                           shift_out(53) => negative_inputs_21_53_port, 
                           shift_out(52) => negative_inputs_21_52_port, 
                           shift_out(51) => negative_inputs_21_51_port, 
                           shift_out(50) => negative_inputs_21_50_port, 
                           shift_out(49) => negative_inputs_21_49_port, 
                           shift_out(48) => negative_inputs_21_48_port, 
                           shift_out(47) => negative_inputs_21_47_port, 
                           shift_out(46) => negative_inputs_21_46_port, 
                           shift_out(45) => negative_inputs_21_45_port, 
                           shift_out(44) => negative_inputs_21_44_port, 
                           shift_out(43) => negative_inputs_21_43_port, 
                           shift_out(42) => negative_inputs_21_42_port, 
                           shift_out(41) => negative_inputs_21_41_port, 
                           shift_out(40) => negative_inputs_21_40_port, 
                           shift_out(39) => negative_inputs_21_39_port, 
                           shift_out(38) => negative_inputs_21_38_port, 
                           shift_out(37) => negative_inputs_21_37_port, 
                           shift_out(36) => negative_inputs_21_36_port, 
                           shift_out(35) => negative_inputs_21_35_port, 
                           shift_out(34) => negative_inputs_21_34_port, 
                           shift_out(33) => negative_inputs_21_33_port, 
                           shift_out(32) => negative_inputs_21_32_port, 
                           shift_out(31) => negative_inputs_21_31_port, 
                           shift_out(30) => negative_inputs_21_30_port, 
                           shift_out(29) => negative_inputs_21_29_port, 
                           shift_out(28) => negative_inputs_21_28_port, 
                           shift_out(27) => negative_inputs_21_27_port, 
                           shift_out(26) => negative_inputs_21_26_port, 
                           shift_out(25) => negative_inputs_21_25_port, 
                           shift_out(24) => negative_inputs_21_24_port, 
                           shift_out(23) => negative_inputs_21_23_port, 
                           shift_out(22) => negative_inputs_21_22_port, 
                           shift_out(21) => negative_inputs_21_21_port, 
                           shift_out(20) => negative_inputs_21_20_port, 
                           shift_out(19) => negative_inputs_21_19_port, 
                           shift_out(18) => negative_inputs_21_18_port, 
                           shift_out(17) => negative_inputs_21_17_port, 
                           shift_out(16) => negative_inputs_21_16_port, 
                           shift_out(15) => negative_inputs_21_15_port, 
                           shift_out(14) => negative_inputs_21_14_port, 
                           shift_out(13) => negative_inputs_21_13_port, 
                           shift_out(12) => negative_inputs_21_12_port, 
                           shift_out(11) => negative_inputs_21_11_port, 
                           shift_out(10) => negative_inputs_21_10_port, 
                           shift_out(9) => negative_inputs_21_9_port, 
                           shift_out(8) => negative_inputs_21_8_port, 
                           shift_out(7) => negative_inputs_21_7_port, 
                           shift_out(6) => negative_inputs_21_6_port, 
                           shift_out(5) => negative_inputs_21_5_port, 
                           shift_out(4) => negative_inputs_21_4_port, 
                           shift_out(3) => negative_inputs_21_3_port, 
                           shift_out(2) => negative_inputs_21_2_port, 
                           shift_out(1) => negative_inputs_21_1_port, 
                           shift_out(0) => n_1116);
   shifted_neg_22 : leftshifter_NbitShifter64_10 port map( shift_in(63) => 
                           negative_inputs_21_63_port, shift_in(62) => 
                           negative_inputs_21_62_port, shift_in(61) => 
                           negative_inputs_21_61_port, shift_in(60) => 
                           negative_inputs_21_60_port, shift_in(59) => 
                           negative_inputs_21_59_port, shift_in(58) => 
                           negative_inputs_21_58_port, shift_in(57) => 
                           negative_inputs_21_57_port, shift_in(56) => 
                           negative_inputs_21_56_port, shift_in(55) => 
                           negative_inputs_21_55_port, shift_in(54) => 
                           negative_inputs_21_54_port, shift_in(53) => 
                           negative_inputs_21_53_port, shift_in(52) => 
                           negative_inputs_21_52_port, shift_in(51) => 
                           negative_inputs_21_51_port, shift_in(50) => 
                           negative_inputs_21_50_port, shift_in(49) => 
                           negative_inputs_21_49_port, shift_in(48) => 
                           negative_inputs_21_48_port, shift_in(47) => 
                           negative_inputs_21_47_port, shift_in(46) => 
                           negative_inputs_21_46_port, shift_in(45) => 
                           negative_inputs_21_45_port, shift_in(44) => 
                           negative_inputs_21_44_port, shift_in(43) => 
                           negative_inputs_21_43_port, shift_in(42) => 
                           negative_inputs_21_42_port, shift_in(41) => 
                           negative_inputs_21_41_port, shift_in(40) => 
                           negative_inputs_21_40_port, shift_in(39) => 
                           negative_inputs_21_39_port, shift_in(38) => 
                           negative_inputs_21_38_port, shift_in(37) => 
                           negative_inputs_21_37_port, shift_in(36) => 
                           negative_inputs_21_36_port, shift_in(35) => 
                           negative_inputs_21_35_port, shift_in(34) => 
                           negative_inputs_21_34_port, shift_in(33) => 
                           negative_inputs_21_33_port, shift_in(32) => 
                           negative_inputs_21_32_port, shift_in(31) => 
                           negative_inputs_21_31_port, shift_in(30) => 
                           negative_inputs_21_30_port, shift_in(29) => 
                           negative_inputs_21_29_port, shift_in(28) => 
                           negative_inputs_21_28_port, shift_in(27) => 
                           negative_inputs_21_27_port, shift_in(26) => 
                           negative_inputs_21_26_port, shift_in(25) => 
                           negative_inputs_21_25_port, shift_in(24) => 
                           negative_inputs_21_24_port, shift_in(23) => 
                           negative_inputs_21_23_port, shift_in(22) => 
                           negative_inputs_21_22_port, shift_in(21) => 
                           negative_inputs_21_21_port, shift_in(20) => 
                           negative_inputs_21_20_port, shift_in(19) => 
                           negative_inputs_21_19_port, shift_in(18) => 
                           negative_inputs_21_18_port, shift_in(17) => 
                           negative_inputs_21_17_port, shift_in(16) => 
                           negative_inputs_21_16_port, shift_in(15) => 
                           negative_inputs_21_15_port, shift_in(14) => 
                           negative_inputs_21_14_port, shift_in(13) => 
                           negative_inputs_21_13_port, shift_in(12) => 
                           negative_inputs_21_12_port, shift_in(11) => 
                           negative_inputs_21_11_port, shift_in(10) => 
                           negative_inputs_21_10_port, shift_in(9) => 
                           negative_inputs_21_9_port, shift_in(8) => 
                           negative_inputs_21_8_port, shift_in(7) => 
                           negative_inputs_21_7_port, shift_in(6) => 
                           negative_inputs_21_6_port, shift_in(5) => 
                           negative_inputs_21_5_port, shift_in(4) => 
                           negative_inputs_21_4_port, shift_in(3) => 
                           negative_inputs_21_3_port, shift_in(2) => 
                           negative_inputs_21_2_port, shift_in(1) => 
                           negative_inputs_21_1_port, shift_in(0) => n9, 
                           shift_out(63) => negative_inputs_22_63_port, 
                           shift_out(62) => negative_inputs_22_62_port, 
                           shift_out(61) => negative_inputs_22_61_port, 
                           shift_out(60) => negative_inputs_22_60_port, 
                           shift_out(59) => negative_inputs_22_59_port, 
                           shift_out(58) => negative_inputs_22_58_port, 
                           shift_out(57) => negative_inputs_22_57_port, 
                           shift_out(56) => negative_inputs_22_56_port, 
                           shift_out(55) => negative_inputs_22_55_port, 
                           shift_out(54) => negative_inputs_22_54_port, 
                           shift_out(53) => negative_inputs_22_53_port, 
                           shift_out(52) => negative_inputs_22_52_port, 
                           shift_out(51) => negative_inputs_22_51_port, 
                           shift_out(50) => negative_inputs_22_50_port, 
                           shift_out(49) => negative_inputs_22_49_port, 
                           shift_out(48) => negative_inputs_22_48_port, 
                           shift_out(47) => negative_inputs_22_47_port, 
                           shift_out(46) => negative_inputs_22_46_port, 
                           shift_out(45) => negative_inputs_22_45_port, 
                           shift_out(44) => negative_inputs_22_44_port, 
                           shift_out(43) => negative_inputs_22_43_port, 
                           shift_out(42) => negative_inputs_22_42_port, 
                           shift_out(41) => negative_inputs_22_41_port, 
                           shift_out(40) => negative_inputs_22_40_port, 
                           shift_out(39) => negative_inputs_22_39_port, 
                           shift_out(38) => negative_inputs_22_38_port, 
                           shift_out(37) => negative_inputs_22_37_port, 
                           shift_out(36) => negative_inputs_22_36_port, 
                           shift_out(35) => negative_inputs_22_35_port, 
                           shift_out(34) => negative_inputs_22_34_port, 
                           shift_out(33) => negative_inputs_22_33_port, 
                           shift_out(32) => negative_inputs_22_32_port, 
                           shift_out(31) => negative_inputs_22_31_port, 
                           shift_out(30) => negative_inputs_22_30_port, 
                           shift_out(29) => negative_inputs_22_29_port, 
                           shift_out(28) => negative_inputs_22_28_port, 
                           shift_out(27) => negative_inputs_22_27_port, 
                           shift_out(26) => negative_inputs_22_26_port, 
                           shift_out(25) => negative_inputs_22_25_port, 
                           shift_out(24) => negative_inputs_22_24_port, 
                           shift_out(23) => negative_inputs_22_23_port, 
                           shift_out(22) => negative_inputs_22_22_port, 
                           shift_out(21) => negative_inputs_22_21_port, 
                           shift_out(20) => negative_inputs_22_20_port, 
                           shift_out(19) => negative_inputs_22_19_port, 
                           shift_out(18) => negative_inputs_22_18_port, 
                           shift_out(17) => negative_inputs_22_17_port, 
                           shift_out(16) => negative_inputs_22_16_port, 
                           shift_out(15) => negative_inputs_22_15_port, 
                           shift_out(14) => negative_inputs_22_14_port, 
                           shift_out(13) => negative_inputs_22_13_port, 
                           shift_out(12) => negative_inputs_22_12_port, 
                           shift_out(11) => negative_inputs_22_11_port, 
                           shift_out(10) => negative_inputs_22_10_port, 
                           shift_out(9) => negative_inputs_22_9_port, 
                           shift_out(8) => negative_inputs_22_8_port, 
                           shift_out(7) => negative_inputs_22_7_port, 
                           shift_out(6) => negative_inputs_22_6_port, 
                           shift_out(5) => negative_inputs_22_5_port, 
                           shift_out(4) => negative_inputs_22_4_port, 
                           shift_out(3) => negative_inputs_22_3_port, 
                           shift_out(2) => negative_inputs_22_2_port, 
                           shift_out(1) => negative_inputs_22_1_port, 
                           shift_out(0) => n_1117);
   shifted_neg_23 : leftshifter_NbitShifter64_9 port map( shift_in(63) => 
                           negative_inputs_22_63_port, shift_in(62) => 
                           negative_inputs_22_62_port, shift_in(61) => 
                           negative_inputs_22_61_port, shift_in(60) => 
                           negative_inputs_22_60_port, shift_in(59) => 
                           negative_inputs_22_59_port, shift_in(58) => 
                           negative_inputs_22_58_port, shift_in(57) => 
                           negative_inputs_22_57_port, shift_in(56) => 
                           negative_inputs_22_56_port, shift_in(55) => 
                           negative_inputs_22_55_port, shift_in(54) => 
                           negative_inputs_22_54_port, shift_in(53) => 
                           negative_inputs_22_53_port, shift_in(52) => 
                           negative_inputs_22_52_port, shift_in(51) => 
                           negative_inputs_22_51_port, shift_in(50) => 
                           negative_inputs_22_50_port, shift_in(49) => 
                           negative_inputs_22_49_port, shift_in(48) => 
                           negative_inputs_22_48_port, shift_in(47) => 
                           negative_inputs_22_47_port, shift_in(46) => 
                           negative_inputs_22_46_port, shift_in(45) => 
                           negative_inputs_22_45_port, shift_in(44) => 
                           negative_inputs_22_44_port, shift_in(43) => 
                           negative_inputs_22_43_port, shift_in(42) => 
                           negative_inputs_22_42_port, shift_in(41) => 
                           negative_inputs_22_41_port, shift_in(40) => 
                           negative_inputs_22_40_port, shift_in(39) => 
                           negative_inputs_22_39_port, shift_in(38) => 
                           negative_inputs_22_38_port, shift_in(37) => 
                           negative_inputs_22_37_port, shift_in(36) => 
                           negative_inputs_22_36_port, shift_in(35) => 
                           negative_inputs_22_35_port, shift_in(34) => 
                           negative_inputs_22_34_port, shift_in(33) => 
                           negative_inputs_22_33_port, shift_in(32) => 
                           negative_inputs_22_32_port, shift_in(31) => 
                           negative_inputs_22_31_port, shift_in(30) => 
                           negative_inputs_22_30_port, shift_in(29) => 
                           negative_inputs_22_29_port, shift_in(28) => 
                           negative_inputs_22_28_port, shift_in(27) => 
                           negative_inputs_22_27_port, shift_in(26) => 
                           negative_inputs_22_26_port, shift_in(25) => 
                           negative_inputs_22_25_port, shift_in(24) => 
                           negative_inputs_22_24_port, shift_in(23) => 
                           negative_inputs_22_23_port, shift_in(22) => 
                           negative_inputs_22_22_port, shift_in(21) => 
                           negative_inputs_22_21_port, shift_in(20) => 
                           negative_inputs_22_20_port, shift_in(19) => 
                           negative_inputs_22_19_port, shift_in(18) => 
                           negative_inputs_22_18_port, shift_in(17) => 
                           negative_inputs_22_17_port, shift_in(16) => 
                           negative_inputs_22_16_port, shift_in(15) => 
                           negative_inputs_22_15_port, shift_in(14) => 
                           negative_inputs_22_14_port, shift_in(13) => 
                           negative_inputs_22_13_port, shift_in(12) => 
                           negative_inputs_22_12_port, shift_in(11) => 
                           negative_inputs_22_11_port, shift_in(10) => 
                           negative_inputs_22_10_port, shift_in(9) => 
                           negative_inputs_22_9_port, shift_in(8) => 
                           negative_inputs_22_8_port, shift_in(7) => 
                           negative_inputs_22_7_port, shift_in(6) => 
                           negative_inputs_22_6_port, shift_in(5) => 
                           negative_inputs_22_5_port, shift_in(4) => 
                           negative_inputs_22_4_port, shift_in(3) => 
                           negative_inputs_22_3_port, shift_in(2) => 
                           negative_inputs_22_2_port, shift_in(1) => 
                           negative_inputs_22_1_port, shift_in(0) => n9, 
                           shift_out(63) => negative_inputs_23_63_port, 
                           shift_out(62) => negative_inputs_23_62_port, 
                           shift_out(61) => negative_inputs_23_61_port, 
                           shift_out(60) => negative_inputs_23_60_port, 
                           shift_out(59) => negative_inputs_23_59_port, 
                           shift_out(58) => negative_inputs_23_58_port, 
                           shift_out(57) => negative_inputs_23_57_port, 
                           shift_out(56) => negative_inputs_23_56_port, 
                           shift_out(55) => negative_inputs_23_55_port, 
                           shift_out(54) => negative_inputs_23_54_port, 
                           shift_out(53) => negative_inputs_23_53_port, 
                           shift_out(52) => negative_inputs_23_52_port, 
                           shift_out(51) => negative_inputs_23_51_port, 
                           shift_out(50) => negative_inputs_23_50_port, 
                           shift_out(49) => negative_inputs_23_49_port, 
                           shift_out(48) => negative_inputs_23_48_port, 
                           shift_out(47) => negative_inputs_23_47_port, 
                           shift_out(46) => negative_inputs_23_46_port, 
                           shift_out(45) => negative_inputs_23_45_port, 
                           shift_out(44) => negative_inputs_23_44_port, 
                           shift_out(43) => negative_inputs_23_43_port, 
                           shift_out(42) => negative_inputs_23_42_port, 
                           shift_out(41) => negative_inputs_23_41_port, 
                           shift_out(40) => negative_inputs_23_40_port, 
                           shift_out(39) => negative_inputs_23_39_port, 
                           shift_out(38) => negative_inputs_23_38_port, 
                           shift_out(37) => negative_inputs_23_37_port, 
                           shift_out(36) => negative_inputs_23_36_port, 
                           shift_out(35) => negative_inputs_23_35_port, 
                           shift_out(34) => negative_inputs_23_34_port, 
                           shift_out(33) => negative_inputs_23_33_port, 
                           shift_out(32) => negative_inputs_23_32_port, 
                           shift_out(31) => negative_inputs_23_31_port, 
                           shift_out(30) => negative_inputs_23_30_port, 
                           shift_out(29) => negative_inputs_23_29_port, 
                           shift_out(28) => negative_inputs_23_28_port, 
                           shift_out(27) => negative_inputs_23_27_port, 
                           shift_out(26) => negative_inputs_23_26_port, 
                           shift_out(25) => negative_inputs_23_25_port, 
                           shift_out(24) => negative_inputs_23_24_port, 
                           shift_out(23) => negative_inputs_23_23_port, 
                           shift_out(22) => negative_inputs_23_22_port, 
                           shift_out(21) => negative_inputs_23_21_port, 
                           shift_out(20) => negative_inputs_23_20_port, 
                           shift_out(19) => negative_inputs_23_19_port, 
                           shift_out(18) => negative_inputs_23_18_port, 
                           shift_out(17) => negative_inputs_23_17_port, 
                           shift_out(16) => negative_inputs_23_16_port, 
                           shift_out(15) => negative_inputs_23_15_port, 
                           shift_out(14) => negative_inputs_23_14_port, 
                           shift_out(13) => negative_inputs_23_13_port, 
                           shift_out(12) => negative_inputs_23_12_port, 
                           shift_out(11) => negative_inputs_23_11_port, 
                           shift_out(10) => negative_inputs_23_10_port, 
                           shift_out(9) => negative_inputs_23_9_port, 
                           shift_out(8) => negative_inputs_23_8_port, 
                           shift_out(7) => negative_inputs_23_7_port, 
                           shift_out(6) => negative_inputs_23_6_port, 
                           shift_out(5) => negative_inputs_23_5_port, 
                           shift_out(4) => negative_inputs_23_4_port, 
                           shift_out(3) => negative_inputs_23_3_port, 
                           shift_out(2) => negative_inputs_23_2_port, 
                           shift_out(1) => negative_inputs_23_1_port, 
                           shift_out(0) => n_1118);
   shifted_neg_24 : leftshifter_NbitShifter64_8 port map( shift_in(63) => 
                           negative_inputs_23_63_port, shift_in(62) => 
                           negative_inputs_23_62_port, shift_in(61) => 
                           negative_inputs_23_61_port, shift_in(60) => 
                           negative_inputs_23_60_port, shift_in(59) => 
                           negative_inputs_23_59_port, shift_in(58) => 
                           negative_inputs_23_58_port, shift_in(57) => 
                           negative_inputs_23_57_port, shift_in(56) => 
                           negative_inputs_23_56_port, shift_in(55) => 
                           negative_inputs_23_55_port, shift_in(54) => 
                           negative_inputs_23_54_port, shift_in(53) => 
                           negative_inputs_23_53_port, shift_in(52) => 
                           negative_inputs_23_52_port, shift_in(51) => 
                           negative_inputs_23_51_port, shift_in(50) => 
                           negative_inputs_23_50_port, shift_in(49) => 
                           negative_inputs_23_49_port, shift_in(48) => 
                           negative_inputs_23_48_port, shift_in(47) => 
                           negative_inputs_23_47_port, shift_in(46) => 
                           negative_inputs_23_46_port, shift_in(45) => 
                           negative_inputs_23_45_port, shift_in(44) => 
                           negative_inputs_23_44_port, shift_in(43) => 
                           negative_inputs_23_43_port, shift_in(42) => 
                           negative_inputs_23_42_port, shift_in(41) => 
                           negative_inputs_23_41_port, shift_in(40) => 
                           negative_inputs_23_40_port, shift_in(39) => 
                           negative_inputs_23_39_port, shift_in(38) => 
                           negative_inputs_23_38_port, shift_in(37) => 
                           negative_inputs_23_37_port, shift_in(36) => 
                           negative_inputs_23_36_port, shift_in(35) => 
                           negative_inputs_23_35_port, shift_in(34) => 
                           negative_inputs_23_34_port, shift_in(33) => 
                           negative_inputs_23_33_port, shift_in(32) => 
                           negative_inputs_23_32_port, shift_in(31) => 
                           negative_inputs_23_31_port, shift_in(30) => 
                           negative_inputs_23_30_port, shift_in(29) => 
                           negative_inputs_23_29_port, shift_in(28) => 
                           negative_inputs_23_28_port, shift_in(27) => 
                           negative_inputs_23_27_port, shift_in(26) => 
                           negative_inputs_23_26_port, shift_in(25) => 
                           negative_inputs_23_25_port, shift_in(24) => 
                           negative_inputs_23_24_port, shift_in(23) => 
                           negative_inputs_23_23_port, shift_in(22) => 
                           negative_inputs_23_22_port, shift_in(21) => 
                           negative_inputs_23_21_port, shift_in(20) => 
                           negative_inputs_23_20_port, shift_in(19) => 
                           negative_inputs_23_19_port, shift_in(18) => 
                           negative_inputs_23_18_port, shift_in(17) => 
                           negative_inputs_23_17_port, shift_in(16) => 
                           negative_inputs_23_16_port, shift_in(15) => 
                           negative_inputs_23_15_port, shift_in(14) => 
                           negative_inputs_23_14_port, shift_in(13) => 
                           negative_inputs_23_13_port, shift_in(12) => 
                           negative_inputs_23_12_port, shift_in(11) => 
                           negative_inputs_23_11_port, shift_in(10) => 
                           negative_inputs_23_10_port, shift_in(9) => 
                           negative_inputs_23_9_port, shift_in(8) => 
                           negative_inputs_23_8_port, shift_in(7) => 
                           negative_inputs_23_7_port, shift_in(6) => 
                           negative_inputs_23_6_port, shift_in(5) => 
                           negative_inputs_23_5_port, shift_in(4) => 
                           negative_inputs_23_4_port, shift_in(3) => 
                           negative_inputs_23_3_port, shift_in(2) => 
                           negative_inputs_23_2_port, shift_in(1) => 
                           negative_inputs_23_1_port, shift_in(0) => n9, 
                           shift_out(63) => negative_inputs_24_63_port, 
                           shift_out(62) => negative_inputs_24_62_port, 
                           shift_out(61) => negative_inputs_24_61_port, 
                           shift_out(60) => negative_inputs_24_60_port, 
                           shift_out(59) => negative_inputs_24_59_port, 
                           shift_out(58) => negative_inputs_24_58_port, 
                           shift_out(57) => negative_inputs_24_57_port, 
                           shift_out(56) => negative_inputs_24_56_port, 
                           shift_out(55) => negative_inputs_24_55_port, 
                           shift_out(54) => negative_inputs_24_54_port, 
                           shift_out(53) => negative_inputs_24_53_port, 
                           shift_out(52) => negative_inputs_24_52_port, 
                           shift_out(51) => negative_inputs_24_51_port, 
                           shift_out(50) => negative_inputs_24_50_port, 
                           shift_out(49) => negative_inputs_24_49_port, 
                           shift_out(48) => negative_inputs_24_48_port, 
                           shift_out(47) => negative_inputs_24_47_port, 
                           shift_out(46) => negative_inputs_24_46_port, 
                           shift_out(45) => negative_inputs_24_45_port, 
                           shift_out(44) => negative_inputs_24_44_port, 
                           shift_out(43) => negative_inputs_24_43_port, 
                           shift_out(42) => negative_inputs_24_42_port, 
                           shift_out(41) => negative_inputs_24_41_port, 
                           shift_out(40) => negative_inputs_24_40_port, 
                           shift_out(39) => negative_inputs_24_39_port, 
                           shift_out(38) => negative_inputs_24_38_port, 
                           shift_out(37) => negative_inputs_24_37_port, 
                           shift_out(36) => negative_inputs_24_36_port, 
                           shift_out(35) => negative_inputs_24_35_port, 
                           shift_out(34) => negative_inputs_24_34_port, 
                           shift_out(33) => negative_inputs_24_33_port, 
                           shift_out(32) => negative_inputs_24_32_port, 
                           shift_out(31) => negative_inputs_24_31_port, 
                           shift_out(30) => negative_inputs_24_30_port, 
                           shift_out(29) => negative_inputs_24_29_port, 
                           shift_out(28) => negative_inputs_24_28_port, 
                           shift_out(27) => negative_inputs_24_27_port, 
                           shift_out(26) => negative_inputs_24_26_port, 
                           shift_out(25) => negative_inputs_24_25_port, 
                           shift_out(24) => negative_inputs_24_24_port, 
                           shift_out(23) => negative_inputs_24_23_port, 
                           shift_out(22) => negative_inputs_24_22_port, 
                           shift_out(21) => negative_inputs_24_21_port, 
                           shift_out(20) => negative_inputs_24_20_port, 
                           shift_out(19) => negative_inputs_24_19_port, 
                           shift_out(18) => negative_inputs_24_18_port, 
                           shift_out(17) => negative_inputs_24_17_port, 
                           shift_out(16) => negative_inputs_24_16_port, 
                           shift_out(15) => negative_inputs_24_15_port, 
                           shift_out(14) => negative_inputs_24_14_port, 
                           shift_out(13) => negative_inputs_24_13_port, 
                           shift_out(12) => negative_inputs_24_12_port, 
                           shift_out(11) => negative_inputs_24_11_port, 
                           shift_out(10) => negative_inputs_24_10_port, 
                           shift_out(9) => negative_inputs_24_9_port, 
                           shift_out(8) => negative_inputs_24_8_port, 
                           shift_out(7) => negative_inputs_24_7_port, 
                           shift_out(6) => negative_inputs_24_6_port, 
                           shift_out(5) => negative_inputs_24_5_port, 
                           shift_out(4) => negative_inputs_24_4_port, 
                           shift_out(3) => negative_inputs_24_3_port, 
                           shift_out(2) => negative_inputs_24_2_port, 
                           shift_out(1) => negative_inputs_24_1_port, 
                           shift_out(0) => n_1119);
   shifted_neg_25 : leftshifter_NbitShifter64_7 port map( shift_in(63) => 
                           negative_inputs_24_63_port, shift_in(62) => 
                           negative_inputs_24_62_port, shift_in(61) => 
                           negative_inputs_24_61_port, shift_in(60) => 
                           negative_inputs_24_60_port, shift_in(59) => 
                           negative_inputs_24_59_port, shift_in(58) => 
                           negative_inputs_24_58_port, shift_in(57) => 
                           negative_inputs_24_57_port, shift_in(56) => 
                           negative_inputs_24_56_port, shift_in(55) => 
                           negative_inputs_24_55_port, shift_in(54) => 
                           negative_inputs_24_54_port, shift_in(53) => 
                           negative_inputs_24_53_port, shift_in(52) => 
                           negative_inputs_24_52_port, shift_in(51) => 
                           negative_inputs_24_51_port, shift_in(50) => 
                           negative_inputs_24_50_port, shift_in(49) => 
                           negative_inputs_24_49_port, shift_in(48) => 
                           negative_inputs_24_48_port, shift_in(47) => 
                           negative_inputs_24_47_port, shift_in(46) => 
                           negative_inputs_24_46_port, shift_in(45) => 
                           negative_inputs_24_45_port, shift_in(44) => 
                           negative_inputs_24_44_port, shift_in(43) => 
                           negative_inputs_24_43_port, shift_in(42) => 
                           negative_inputs_24_42_port, shift_in(41) => 
                           negative_inputs_24_41_port, shift_in(40) => 
                           negative_inputs_24_40_port, shift_in(39) => 
                           negative_inputs_24_39_port, shift_in(38) => 
                           negative_inputs_24_38_port, shift_in(37) => 
                           negative_inputs_24_37_port, shift_in(36) => 
                           negative_inputs_24_36_port, shift_in(35) => 
                           negative_inputs_24_35_port, shift_in(34) => 
                           negative_inputs_24_34_port, shift_in(33) => 
                           negative_inputs_24_33_port, shift_in(32) => 
                           negative_inputs_24_32_port, shift_in(31) => 
                           negative_inputs_24_31_port, shift_in(30) => 
                           negative_inputs_24_30_port, shift_in(29) => 
                           negative_inputs_24_29_port, shift_in(28) => 
                           negative_inputs_24_28_port, shift_in(27) => 
                           negative_inputs_24_27_port, shift_in(26) => 
                           negative_inputs_24_26_port, shift_in(25) => 
                           negative_inputs_24_25_port, shift_in(24) => 
                           negative_inputs_24_24_port, shift_in(23) => 
                           negative_inputs_24_23_port, shift_in(22) => 
                           negative_inputs_24_22_port, shift_in(21) => 
                           negative_inputs_24_21_port, shift_in(20) => 
                           negative_inputs_24_20_port, shift_in(19) => 
                           negative_inputs_24_19_port, shift_in(18) => 
                           negative_inputs_24_18_port, shift_in(17) => 
                           negative_inputs_24_17_port, shift_in(16) => 
                           negative_inputs_24_16_port, shift_in(15) => 
                           negative_inputs_24_15_port, shift_in(14) => 
                           negative_inputs_24_14_port, shift_in(13) => 
                           negative_inputs_24_13_port, shift_in(12) => 
                           negative_inputs_24_12_port, shift_in(11) => 
                           negative_inputs_24_11_port, shift_in(10) => 
                           negative_inputs_24_10_port, shift_in(9) => 
                           negative_inputs_24_9_port, shift_in(8) => 
                           negative_inputs_24_8_port, shift_in(7) => 
                           negative_inputs_24_7_port, shift_in(6) => 
                           negative_inputs_24_6_port, shift_in(5) => 
                           negative_inputs_24_5_port, shift_in(4) => 
                           negative_inputs_24_4_port, shift_in(3) => 
                           negative_inputs_24_3_port, shift_in(2) => 
                           negative_inputs_24_2_port, shift_in(1) => 
                           negative_inputs_24_1_port, shift_in(0) => n9, 
                           shift_out(63) => negative_inputs_25_63_port, 
                           shift_out(62) => negative_inputs_25_62_port, 
                           shift_out(61) => negative_inputs_25_61_port, 
                           shift_out(60) => negative_inputs_25_60_port, 
                           shift_out(59) => negative_inputs_25_59_port, 
                           shift_out(58) => negative_inputs_25_58_port, 
                           shift_out(57) => negative_inputs_25_57_port, 
                           shift_out(56) => negative_inputs_25_56_port, 
                           shift_out(55) => negative_inputs_25_55_port, 
                           shift_out(54) => negative_inputs_25_54_port, 
                           shift_out(53) => negative_inputs_25_53_port, 
                           shift_out(52) => negative_inputs_25_52_port, 
                           shift_out(51) => negative_inputs_25_51_port, 
                           shift_out(50) => negative_inputs_25_50_port, 
                           shift_out(49) => negative_inputs_25_49_port, 
                           shift_out(48) => negative_inputs_25_48_port, 
                           shift_out(47) => negative_inputs_25_47_port, 
                           shift_out(46) => negative_inputs_25_46_port, 
                           shift_out(45) => negative_inputs_25_45_port, 
                           shift_out(44) => negative_inputs_25_44_port, 
                           shift_out(43) => negative_inputs_25_43_port, 
                           shift_out(42) => negative_inputs_25_42_port, 
                           shift_out(41) => negative_inputs_25_41_port, 
                           shift_out(40) => negative_inputs_25_40_port, 
                           shift_out(39) => negative_inputs_25_39_port, 
                           shift_out(38) => negative_inputs_25_38_port, 
                           shift_out(37) => negative_inputs_25_37_port, 
                           shift_out(36) => negative_inputs_25_36_port, 
                           shift_out(35) => negative_inputs_25_35_port, 
                           shift_out(34) => negative_inputs_25_34_port, 
                           shift_out(33) => negative_inputs_25_33_port, 
                           shift_out(32) => negative_inputs_25_32_port, 
                           shift_out(31) => negative_inputs_25_31_port, 
                           shift_out(30) => negative_inputs_25_30_port, 
                           shift_out(29) => negative_inputs_25_29_port, 
                           shift_out(28) => negative_inputs_25_28_port, 
                           shift_out(27) => negative_inputs_25_27_port, 
                           shift_out(26) => negative_inputs_25_26_port, 
                           shift_out(25) => negative_inputs_25_25_port, 
                           shift_out(24) => negative_inputs_25_24_port, 
                           shift_out(23) => negative_inputs_25_23_port, 
                           shift_out(22) => negative_inputs_25_22_port, 
                           shift_out(21) => negative_inputs_25_21_port, 
                           shift_out(20) => negative_inputs_25_20_port, 
                           shift_out(19) => negative_inputs_25_19_port, 
                           shift_out(18) => negative_inputs_25_18_port, 
                           shift_out(17) => negative_inputs_25_17_port, 
                           shift_out(16) => negative_inputs_25_16_port, 
                           shift_out(15) => negative_inputs_25_15_port, 
                           shift_out(14) => negative_inputs_25_14_port, 
                           shift_out(13) => negative_inputs_25_13_port, 
                           shift_out(12) => negative_inputs_25_12_port, 
                           shift_out(11) => negative_inputs_25_11_port, 
                           shift_out(10) => negative_inputs_25_10_port, 
                           shift_out(9) => negative_inputs_25_9_port, 
                           shift_out(8) => negative_inputs_25_8_port, 
                           shift_out(7) => negative_inputs_25_7_port, 
                           shift_out(6) => negative_inputs_25_6_port, 
                           shift_out(5) => negative_inputs_25_5_port, 
                           shift_out(4) => negative_inputs_25_4_port, 
                           shift_out(3) => negative_inputs_25_3_port, 
                           shift_out(2) => negative_inputs_25_2_port, 
                           shift_out(1) => negative_inputs_25_1_port, 
                           shift_out(0) => n_1120);
   shifted_neg_26 : leftshifter_NbitShifter64_6 port map( shift_in(63) => 
                           negative_inputs_25_63_port, shift_in(62) => 
                           negative_inputs_25_62_port, shift_in(61) => 
                           negative_inputs_25_61_port, shift_in(60) => 
                           negative_inputs_25_60_port, shift_in(59) => 
                           negative_inputs_25_59_port, shift_in(58) => 
                           negative_inputs_25_58_port, shift_in(57) => 
                           negative_inputs_25_57_port, shift_in(56) => 
                           negative_inputs_25_56_port, shift_in(55) => 
                           negative_inputs_25_55_port, shift_in(54) => 
                           negative_inputs_25_54_port, shift_in(53) => 
                           negative_inputs_25_53_port, shift_in(52) => 
                           negative_inputs_25_52_port, shift_in(51) => 
                           negative_inputs_25_51_port, shift_in(50) => 
                           negative_inputs_25_50_port, shift_in(49) => 
                           negative_inputs_25_49_port, shift_in(48) => 
                           negative_inputs_25_48_port, shift_in(47) => 
                           negative_inputs_25_47_port, shift_in(46) => 
                           negative_inputs_25_46_port, shift_in(45) => 
                           negative_inputs_25_45_port, shift_in(44) => 
                           negative_inputs_25_44_port, shift_in(43) => 
                           negative_inputs_25_43_port, shift_in(42) => 
                           negative_inputs_25_42_port, shift_in(41) => 
                           negative_inputs_25_41_port, shift_in(40) => 
                           negative_inputs_25_40_port, shift_in(39) => 
                           negative_inputs_25_39_port, shift_in(38) => 
                           negative_inputs_25_38_port, shift_in(37) => 
                           negative_inputs_25_37_port, shift_in(36) => 
                           negative_inputs_25_36_port, shift_in(35) => 
                           negative_inputs_25_35_port, shift_in(34) => 
                           negative_inputs_25_34_port, shift_in(33) => 
                           negative_inputs_25_33_port, shift_in(32) => 
                           negative_inputs_25_32_port, shift_in(31) => 
                           negative_inputs_25_31_port, shift_in(30) => 
                           negative_inputs_25_30_port, shift_in(29) => 
                           negative_inputs_25_29_port, shift_in(28) => 
                           negative_inputs_25_28_port, shift_in(27) => 
                           negative_inputs_25_27_port, shift_in(26) => 
                           negative_inputs_25_26_port, shift_in(25) => 
                           negative_inputs_25_25_port, shift_in(24) => 
                           negative_inputs_25_24_port, shift_in(23) => 
                           negative_inputs_25_23_port, shift_in(22) => 
                           negative_inputs_25_22_port, shift_in(21) => 
                           negative_inputs_25_21_port, shift_in(20) => 
                           negative_inputs_25_20_port, shift_in(19) => 
                           negative_inputs_25_19_port, shift_in(18) => 
                           negative_inputs_25_18_port, shift_in(17) => 
                           negative_inputs_25_17_port, shift_in(16) => 
                           negative_inputs_25_16_port, shift_in(15) => 
                           negative_inputs_25_15_port, shift_in(14) => 
                           negative_inputs_25_14_port, shift_in(13) => 
                           negative_inputs_25_13_port, shift_in(12) => 
                           negative_inputs_25_12_port, shift_in(11) => 
                           negative_inputs_25_11_port, shift_in(10) => 
                           negative_inputs_25_10_port, shift_in(9) => 
                           negative_inputs_25_9_port, shift_in(8) => 
                           negative_inputs_25_8_port, shift_in(7) => 
                           negative_inputs_25_7_port, shift_in(6) => 
                           negative_inputs_25_6_port, shift_in(5) => 
                           negative_inputs_25_5_port, shift_in(4) => 
                           negative_inputs_25_4_port, shift_in(3) => 
                           negative_inputs_25_3_port, shift_in(2) => 
                           negative_inputs_25_2_port, shift_in(1) => 
                           negative_inputs_25_1_port, shift_in(0) => n9, 
                           shift_out(63) => negative_inputs_26_63_port, 
                           shift_out(62) => negative_inputs_26_62_port, 
                           shift_out(61) => negative_inputs_26_61_port, 
                           shift_out(60) => negative_inputs_26_60_port, 
                           shift_out(59) => negative_inputs_26_59_port, 
                           shift_out(58) => negative_inputs_26_58_port, 
                           shift_out(57) => negative_inputs_26_57_port, 
                           shift_out(56) => negative_inputs_26_56_port, 
                           shift_out(55) => negative_inputs_26_55_port, 
                           shift_out(54) => negative_inputs_26_54_port, 
                           shift_out(53) => negative_inputs_26_53_port, 
                           shift_out(52) => negative_inputs_26_52_port, 
                           shift_out(51) => negative_inputs_26_51_port, 
                           shift_out(50) => negative_inputs_26_50_port, 
                           shift_out(49) => negative_inputs_26_49_port, 
                           shift_out(48) => negative_inputs_26_48_port, 
                           shift_out(47) => negative_inputs_26_47_port, 
                           shift_out(46) => negative_inputs_26_46_port, 
                           shift_out(45) => negative_inputs_26_45_port, 
                           shift_out(44) => negative_inputs_26_44_port, 
                           shift_out(43) => negative_inputs_26_43_port, 
                           shift_out(42) => negative_inputs_26_42_port, 
                           shift_out(41) => negative_inputs_26_41_port, 
                           shift_out(40) => negative_inputs_26_40_port, 
                           shift_out(39) => negative_inputs_26_39_port, 
                           shift_out(38) => negative_inputs_26_38_port, 
                           shift_out(37) => negative_inputs_26_37_port, 
                           shift_out(36) => negative_inputs_26_36_port, 
                           shift_out(35) => negative_inputs_26_35_port, 
                           shift_out(34) => negative_inputs_26_34_port, 
                           shift_out(33) => negative_inputs_26_33_port, 
                           shift_out(32) => negative_inputs_26_32_port, 
                           shift_out(31) => negative_inputs_26_31_port, 
                           shift_out(30) => negative_inputs_26_30_port, 
                           shift_out(29) => negative_inputs_26_29_port, 
                           shift_out(28) => negative_inputs_26_28_port, 
                           shift_out(27) => negative_inputs_26_27_port, 
                           shift_out(26) => negative_inputs_26_26_port, 
                           shift_out(25) => negative_inputs_26_25_port, 
                           shift_out(24) => negative_inputs_26_24_port, 
                           shift_out(23) => negative_inputs_26_23_port, 
                           shift_out(22) => negative_inputs_26_22_port, 
                           shift_out(21) => negative_inputs_26_21_port, 
                           shift_out(20) => negative_inputs_26_20_port, 
                           shift_out(19) => negative_inputs_26_19_port, 
                           shift_out(18) => negative_inputs_26_18_port, 
                           shift_out(17) => negative_inputs_26_17_port, 
                           shift_out(16) => negative_inputs_26_16_port, 
                           shift_out(15) => negative_inputs_26_15_port, 
                           shift_out(14) => negative_inputs_26_14_port, 
                           shift_out(13) => negative_inputs_26_13_port, 
                           shift_out(12) => negative_inputs_26_12_port, 
                           shift_out(11) => negative_inputs_26_11_port, 
                           shift_out(10) => negative_inputs_26_10_port, 
                           shift_out(9) => negative_inputs_26_9_port, 
                           shift_out(8) => negative_inputs_26_8_port, 
                           shift_out(7) => negative_inputs_26_7_port, 
                           shift_out(6) => negative_inputs_26_6_port, 
                           shift_out(5) => negative_inputs_26_5_port, 
                           shift_out(4) => negative_inputs_26_4_port, 
                           shift_out(3) => negative_inputs_26_3_port, 
                           shift_out(2) => negative_inputs_26_2_port, 
                           shift_out(1) => negative_inputs_26_1_port, 
                           shift_out(0) => n_1121);
   shifted_neg_27 : leftshifter_NbitShifter64_5 port map( shift_in(63) => 
                           negative_inputs_26_63_port, shift_in(62) => 
                           negative_inputs_26_62_port, shift_in(61) => 
                           negative_inputs_26_61_port, shift_in(60) => 
                           negative_inputs_26_60_port, shift_in(59) => 
                           negative_inputs_26_59_port, shift_in(58) => 
                           negative_inputs_26_58_port, shift_in(57) => 
                           negative_inputs_26_57_port, shift_in(56) => 
                           negative_inputs_26_56_port, shift_in(55) => 
                           negative_inputs_26_55_port, shift_in(54) => 
                           negative_inputs_26_54_port, shift_in(53) => 
                           negative_inputs_26_53_port, shift_in(52) => 
                           negative_inputs_26_52_port, shift_in(51) => 
                           negative_inputs_26_51_port, shift_in(50) => 
                           negative_inputs_26_50_port, shift_in(49) => 
                           negative_inputs_26_49_port, shift_in(48) => 
                           negative_inputs_26_48_port, shift_in(47) => 
                           negative_inputs_26_47_port, shift_in(46) => 
                           negative_inputs_26_46_port, shift_in(45) => 
                           negative_inputs_26_45_port, shift_in(44) => 
                           negative_inputs_26_44_port, shift_in(43) => 
                           negative_inputs_26_43_port, shift_in(42) => 
                           negative_inputs_26_42_port, shift_in(41) => 
                           negative_inputs_26_41_port, shift_in(40) => 
                           negative_inputs_26_40_port, shift_in(39) => 
                           negative_inputs_26_39_port, shift_in(38) => 
                           negative_inputs_26_38_port, shift_in(37) => 
                           negative_inputs_26_37_port, shift_in(36) => 
                           negative_inputs_26_36_port, shift_in(35) => 
                           negative_inputs_26_35_port, shift_in(34) => 
                           negative_inputs_26_34_port, shift_in(33) => 
                           negative_inputs_26_33_port, shift_in(32) => 
                           negative_inputs_26_32_port, shift_in(31) => 
                           negative_inputs_26_31_port, shift_in(30) => 
                           negative_inputs_26_30_port, shift_in(29) => 
                           negative_inputs_26_29_port, shift_in(28) => 
                           negative_inputs_26_28_port, shift_in(27) => 
                           negative_inputs_26_27_port, shift_in(26) => 
                           negative_inputs_26_26_port, shift_in(25) => 
                           negative_inputs_26_25_port, shift_in(24) => 
                           negative_inputs_26_24_port, shift_in(23) => 
                           negative_inputs_26_23_port, shift_in(22) => 
                           negative_inputs_26_22_port, shift_in(21) => 
                           negative_inputs_26_21_port, shift_in(20) => 
                           negative_inputs_26_20_port, shift_in(19) => 
                           negative_inputs_26_19_port, shift_in(18) => 
                           negative_inputs_26_18_port, shift_in(17) => 
                           negative_inputs_26_17_port, shift_in(16) => 
                           negative_inputs_26_16_port, shift_in(15) => 
                           negative_inputs_26_15_port, shift_in(14) => 
                           negative_inputs_26_14_port, shift_in(13) => 
                           negative_inputs_26_13_port, shift_in(12) => 
                           negative_inputs_26_12_port, shift_in(11) => 
                           negative_inputs_26_11_port, shift_in(10) => 
                           negative_inputs_26_10_port, shift_in(9) => 
                           negative_inputs_26_9_port, shift_in(8) => 
                           negative_inputs_26_8_port, shift_in(7) => 
                           negative_inputs_26_7_port, shift_in(6) => 
                           negative_inputs_26_6_port, shift_in(5) => 
                           negative_inputs_26_5_port, shift_in(4) => 
                           negative_inputs_26_4_port, shift_in(3) => 
                           negative_inputs_26_3_port, shift_in(2) => 
                           negative_inputs_26_2_port, shift_in(1) => 
                           negative_inputs_26_1_port, shift_in(0) => n9, 
                           shift_out(63) => negative_inputs_27_63_port, 
                           shift_out(62) => negative_inputs_27_62_port, 
                           shift_out(61) => negative_inputs_27_61_port, 
                           shift_out(60) => negative_inputs_27_60_port, 
                           shift_out(59) => negative_inputs_27_59_port, 
                           shift_out(58) => negative_inputs_27_58_port, 
                           shift_out(57) => negative_inputs_27_57_port, 
                           shift_out(56) => negative_inputs_27_56_port, 
                           shift_out(55) => negative_inputs_27_55_port, 
                           shift_out(54) => negative_inputs_27_54_port, 
                           shift_out(53) => negative_inputs_27_53_port, 
                           shift_out(52) => negative_inputs_27_52_port, 
                           shift_out(51) => negative_inputs_27_51_port, 
                           shift_out(50) => negative_inputs_27_50_port, 
                           shift_out(49) => negative_inputs_27_49_port, 
                           shift_out(48) => negative_inputs_27_48_port, 
                           shift_out(47) => negative_inputs_27_47_port, 
                           shift_out(46) => negative_inputs_27_46_port, 
                           shift_out(45) => negative_inputs_27_45_port, 
                           shift_out(44) => negative_inputs_27_44_port, 
                           shift_out(43) => negative_inputs_27_43_port, 
                           shift_out(42) => negative_inputs_27_42_port, 
                           shift_out(41) => negative_inputs_27_41_port, 
                           shift_out(40) => negative_inputs_27_40_port, 
                           shift_out(39) => negative_inputs_27_39_port, 
                           shift_out(38) => negative_inputs_27_38_port, 
                           shift_out(37) => negative_inputs_27_37_port, 
                           shift_out(36) => negative_inputs_27_36_port, 
                           shift_out(35) => negative_inputs_27_35_port, 
                           shift_out(34) => negative_inputs_27_34_port, 
                           shift_out(33) => negative_inputs_27_33_port, 
                           shift_out(32) => negative_inputs_27_32_port, 
                           shift_out(31) => negative_inputs_27_31_port, 
                           shift_out(30) => negative_inputs_27_30_port, 
                           shift_out(29) => negative_inputs_27_29_port, 
                           shift_out(28) => negative_inputs_27_28_port, 
                           shift_out(27) => negative_inputs_27_27_port, 
                           shift_out(26) => negative_inputs_27_26_port, 
                           shift_out(25) => negative_inputs_27_25_port, 
                           shift_out(24) => negative_inputs_27_24_port, 
                           shift_out(23) => negative_inputs_27_23_port, 
                           shift_out(22) => negative_inputs_27_22_port, 
                           shift_out(21) => negative_inputs_27_21_port, 
                           shift_out(20) => negative_inputs_27_20_port, 
                           shift_out(19) => negative_inputs_27_19_port, 
                           shift_out(18) => negative_inputs_27_18_port, 
                           shift_out(17) => negative_inputs_27_17_port, 
                           shift_out(16) => negative_inputs_27_16_port, 
                           shift_out(15) => negative_inputs_27_15_port, 
                           shift_out(14) => negative_inputs_27_14_port, 
                           shift_out(13) => negative_inputs_27_13_port, 
                           shift_out(12) => negative_inputs_27_12_port, 
                           shift_out(11) => negative_inputs_27_11_port, 
                           shift_out(10) => negative_inputs_27_10_port, 
                           shift_out(9) => negative_inputs_27_9_port, 
                           shift_out(8) => negative_inputs_27_8_port, 
                           shift_out(7) => negative_inputs_27_7_port, 
                           shift_out(6) => negative_inputs_27_6_port, 
                           shift_out(5) => negative_inputs_27_5_port, 
                           shift_out(4) => negative_inputs_27_4_port, 
                           shift_out(3) => negative_inputs_27_3_port, 
                           shift_out(2) => negative_inputs_27_2_port, 
                           shift_out(1) => negative_inputs_27_1_port, 
                           shift_out(0) => n_1122);
   shifted_neg_28 : leftshifter_NbitShifter64_4 port map( shift_in(63) => 
                           negative_inputs_27_63_port, shift_in(62) => 
                           negative_inputs_27_62_port, shift_in(61) => 
                           negative_inputs_27_61_port, shift_in(60) => 
                           negative_inputs_27_60_port, shift_in(59) => 
                           negative_inputs_27_59_port, shift_in(58) => 
                           negative_inputs_27_58_port, shift_in(57) => 
                           negative_inputs_27_57_port, shift_in(56) => 
                           negative_inputs_27_56_port, shift_in(55) => 
                           negative_inputs_27_55_port, shift_in(54) => 
                           negative_inputs_27_54_port, shift_in(53) => 
                           negative_inputs_27_53_port, shift_in(52) => 
                           negative_inputs_27_52_port, shift_in(51) => 
                           negative_inputs_27_51_port, shift_in(50) => 
                           negative_inputs_27_50_port, shift_in(49) => 
                           negative_inputs_27_49_port, shift_in(48) => 
                           negative_inputs_27_48_port, shift_in(47) => 
                           negative_inputs_27_47_port, shift_in(46) => 
                           negative_inputs_27_46_port, shift_in(45) => 
                           negative_inputs_27_45_port, shift_in(44) => 
                           negative_inputs_27_44_port, shift_in(43) => 
                           negative_inputs_27_43_port, shift_in(42) => 
                           negative_inputs_27_42_port, shift_in(41) => 
                           negative_inputs_27_41_port, shift_in(40) => 
                           negative_inputs_27_40_port, shift_in(39) => 
                           negative_inputs_27_39_port, shift_in(38) => 
                           negative_inputs_27_38_port, shift_in(37) => 
                           negative_inputs_27_37_port, shift_in(36) => 
                           negative_inputs_27_36_port, shift_in(35) => 
                           negative_inputs_27_35_port, shift_in(34) => 
                           negative_inputs_27_34_port, shift_in(33) => 
                           negative_inputs_27_33_port, shift_in(32) => 
                           negative_inputs_27_32_port, shift_in(31) => 
                           negative_inputs_27_31_port, shift_in(30) => 
                           negative_inputs_27_30_port, shift_in(29) => 
                           negative_inputs_27_29_port, shift_in(28) => 
                           negative_inputs_27_28_port, shift_in(27) => 
                           negative_inputs_27_27_port, shift_in(26) => 
                           negative_inputs_27_26_port, shift_in(25) => 
                           negative_inputs_27_25_port, shift_in(24) => 
                           negative_inputs_27_24_port, shift_in(23) => 
                           negative_inputs_27_23_port, shift_in(22) => 
                           negative_inputs_27_22_port, shift_in(21) => 
                           negative_inputs_27_21_port, shift_in(20) => 
                           negative_inputs_27_20_port, shift_in(19) => 
                           negative_inputs_27_19_port, shift_in(18) => 
                           negative_inputs_27_18_port, shift_in(17) => 
                           negative_inputs_27_17_port, shift_in(16) => 
                           negative_inputs_27_16_port, shift_in(15) => 
                           negative_inputs_27_15_port, shift_in(14) => 
                           negative_inputs_27_14_port, shift_in(13) => 
                           negative_inputs_27_13_port, shift_in(12) => 
                           negative_inputs_27_12_port, shift_in(11) => 
                           negative_inputs_27_11_port, shift_in(10) => 
                           negative_inputs_27_10_port, shift_in(9) => 
                           negative_inputs_27_9_port, shift_in(8) => 
                           negative_inputs_27_8_port, shift_in(7) => 
                           negative_inputs_27_7_port, shift_in(6) => 
                           negative_inputs_27_6_port, shift_in(5) => 
                           negative_inputs_27_5_port, shift_in(4) => 
                           negative_inputs_27_4_port, shift_in(3) => 
                           negative_inputs_27_3_port, shift_in(2) => 
                           negative_inputs_27_2_port, shift_in(1) => 
                           negative_inputs_27_1_port, shift_in(0) => n9, 
                           shift_out(63) => negative_inputs_28_63_port, 
                           shift_out(62) => negative_inputs_28_62_port, 
                           shift_out(61) => negative_inputs_28_61_port, 
                           shift_out(60) => negative_inputs_28_60_port, 
                           shift_out(59) => negative_inputs_28_59_port, 
                           shift_out(58) => negative_inputs_28_58_port, 
                           shift_out(57) => negative_inputs_28_57_port, 
                           shift_out(56) => negative_inputs_28_56_port, 
                           shift_out(55) => negative_inputs_28_55_port, 
                           shift_out(54) => negative_inputs_28_54_port, 
                           shift_out(53) => negative_inputs_28_53_port, 
                           shift_out(52) => negative_inputs_28_52_port, 
                           shift_out(51) => negative_inputs_28_51_port, 
                           shift_out(50) => negative_inputs_28_50_port, 
                           shift_out(49) => negative_inputs_28_49_port, 
                           shift_out(48) => negative_inputs_28_48_port, 
                           shift_out(47) => negative_inputs_28_47_port, 
                           shift_out(46) => negative_inputs_28_46_port, 
                           shift_out(45) => negative_inputs_28_45_port, 
                           shift_out(44) => negative_inputs_28_44_port, 
                           shift_out(43) => negative_inputs_28_43_port, 
                           shift_out(42) => negative_inputs_28_42_port, 
                           shift_out(41) => negative_inputs_28_41_port, 
                           shift_out(40) => negative_inputs_28_40_port, 
                           shift_out(39) => negative_inputs_28_39_port, 
                           shift_out(38) => negative_inputs_28_38_port, 
                           shift_out(37) => negative_inputs_28_37_port, 
                           shift_out(36) => negative_inputs_28_36_port, 
                           shift_out(35) => negative_inputs_28_35_port, 
                           shift_out(34) => negative_inputs_28_34_port, 
                           shift_out(33) => negative_inputs_28_33_port, 
                           shift_out(32) => negative_inputs_28_32_port, 
                           shift_out(31) => negative_inputs_28_31_port, 
                           shift_out(30) => negative_inputs_28_30_port, 
                           shift_out(29) => negative_inputs_28_29_port, 
                           shift_out(28) => negative_inputs_28_28_port, 
                           shift_out(27) => negative_inputs_28_27_port, 
                           shift_out(26) => negative_inputs_28_26_port, 
                           shift_out(25) => negative_inputs_28_25_port, 
                           shift_out(24) => negative_inputs_28_24_port, 
                           shift_out(23) => negative_inputs_28_23_port, 
                           shift_out(22) => negative_inputs_28_22_port, 
                           shift_out(21) => negative_inputs_28_21_port, 
                           shift_out(20) => negative_inputs_28_20_port, 
                           shift_out(19) => negative_inputs_28_19_port, 
                           shift_out(18) => negative_inputs_28_18_port, 
                           shift_out(17) => negative_inputs_28_17_port, 
                           shift_out(16) => negative_inputs_28_16_port, 
                           shift_out(15) => negative_inputs_28_15_port, 
                           shift_out(14) => negative_inputs_28_14_port, 
                           shift_out(13) => negative_inputs_28_13_port, 
                           shift_out(12) => negative_inputs_28_12_port, 
                           shift_out(11) => negative_inputs_28_11_port, 
                           shift_out(10) => negative_inputs_28_10_port, 
                           shift_out(9) => negative_inputs_28_9_port, 
                           shift_out(8) => negative_inputs_28_8_port, 
                           shift_out(7) => negative_inputs_28_7_port, 
                           shift_out(6) => negative_inputs_28_6_port, 
                           shift_out(5) => negative_inputs_28_5_port, 
                           shift_out(4) => negative_inputs_28_4_port, 
                           shift_out(3) => negative_inputs_28_3_port, 
                           shift_out(2) => negative_inputs_28_2_port, 
                           shift_out(1) => negative_inputs_28_1_port, 
                           shift_out(0) => n_1123);
   shifted_neg_29 : leftshifter_NbitShifter64_3 port map( shift_in(63) => 
                           negative_inputs_28_63_port, shift_in(62) => 
                           negative_inputs_28_62_port, shift_in(61) => 
                           negative_inputs_28_61_port, shift_in(60) => 
                           negative_inputs_28_60_port, shift_in(59) => 
                           negative_inputs_28_59_port, shift_in(58) => 
                           negative_inputs_28_58_port, shift_in(57) => 
                           negative_inputs_28_57_port, shift_in(56) => 
                           negative_inputs_28_56_port, shift_in(55) => 
                           negative_inputs_28_55_port, shift_in(54) => 
                           negative_inputs_28_54_port, shift_in(53) => 
                           negative_inputs_28_53_port, shift_in(52) => 
                           negative_inputs_28_52_port, shift_in(51) => 
                           negative_inputs_28_51_port, shift_in(50) => 
                           negative_inputs_28_50_port, shift_in(49) => 
                           negative_inputs_28_49_port, shift_in(48) => 
                           negative_inputs_28_48_port, shift_in(47) => 
                           negative_inputs_28_47_port, shift_in(46) => 
                           negative_inputs_28_46_port, shift_in(45) => 
                           negative_inputs_28_45_port, shift_in(44) => 
                           negative_inputs_28_44_port, shift_in(43) => 
                           negative_inputs_28_43_port, shift_in(42) => 
                           negative_inputs_28_42_port, shift_in(41) => 
                           negative_inputs_28_41_port, shift_in(40) => 
                           negative_inputs_28_40_port, shift_in(39) => 
                           negative_inputs_28_39_port, shift_in(38) => 
                           negative_inputs_28_38_port, shift_in(37) => 
                           negative_inputs_28_37_port, shift_in(36) => 
                           negative_inputs_28_36_port, shift_in(35) => 
                           negative_inputs_28_35_port, shift_in(34) => 
                           negative_inputs_28_34_port, shift_in(33) => 
                           negative_inputs_28_33_port, shift_in(32) => 
                           negative_inputs_28_32_port, shift_in(31) => 
                           negative_inputs_28_31_port, shift_in(30) => 
                           negative_inputs_28_30_port, shift_in(29) => 
                           negative_inputs_28_29_port, shift_in(28) => 
                           negative_inputs_28_28_port, shift_in(27) => 
                           negative_inputs_28_27_port, shift_in(26) => 
                           negative_inputs_28_26_port, shift_in(25) => 
                           negative_inputs_28_25_port, shift_in(24) => 
                           negative_inputs_28_24_port, shift_in(23) => 
                           negative_inputs_28_23_port, shift_in(22) => 
                           negative_inputs_28_22_port, shift_in(21) => 
                           negative_inputs_28_21_port, shift_in(20) => 
                           negative_inputs_28_20_port, shift_in(19) => 
                           negative_inputs_28_19_port, shift_in(18) => 
                           negative_inputs_28_18_port, shift_in(17) => 
                           negative_inputs_28_17_port, shift_in(16) => 
                           negative_inputs_28_16_port, shift_in(15) => 
                           negative_inputs_28_15_port, shift_in(14) => 
                           negative_inputs_28_14_port, shift_in(13) => 
                           negative_inputs_28_13_port, shift_in(12) => 
                           negative_inputs_28_12_port, shift_in(11) => 
                           negative_inputs_28_11_port, shift_in(10) => 
                           negative_inputs_28_10_port, shift_in(9) => 
                           negative_inputs_28_9_port, shift_in(8) => 
                           negative_inputs_28_8_port, shift_in(7) => 
                           negative_inputs_28_7_port, shift_in(6) => 
                           negative_inputs_28_6_port, shift_in(5) => 
                           negative_inputs_28_5_port, shift_in(4) => 
                           negative_inputs_28_4_port, shift_in(3) => 
                           negative_inputs_28_3_port, shift_in(2) => 
                           negative_inputs_28_2_port, shift_in(1) => 
                           negative_inputs_28_1_port, shift_in(0) => n9, 
                           shift_out(63) => negative_inputs_29_63_port, 
                           shift_out(62) => negative_inputs_29_62_port, 
                           shift_out(61) => negative_inputs_29_61_port, 
                           shift_out(60) => negative_inputs_29_60_port, 
                           shift_out(59) => negative_inputs_29_59_port, 
                           shift_out(58) => negative_inputs_29_58_port, 
                           shift_out(57) => negative_inputs_29_57_port, 
                           shift_out(56) => negative_inputs_29_56_port, 
                           shift_out(55) => negative_inputs_29_55_port, 
                           shift_out(54) => negative_inputs_29_54_port, 
                           shift_out(53) => negative_inputs_29_53_port, 
                           shift_out(52) => negative_inputs_29_52_port, 
                           shift_out(51) => negative_inputs_29_51_port, 
                           shift_out(50) => negative_inputs_29_50_port, 
                           shift_out(49) => negative_inputs_29_49_port, 
                           shift_out(48) => negative_inputs_29_48_port, 
                           shift_out(47) => negative_inputs_29_47_port, 
                           shift_out(46) => negative_inputs_29_46_port, 
                           shift_out(45) => negative_inputs_29_45_port, 
                           shift_out(44) => negative_inputs_29_44_port, 
                           shift_out(43) => negative_inputs_29_43_port, 
                           shift_out(42) => negative_inputs_29_42_port, 
                           shift_out(41) => negative_inputs_29_41_port, 
                           shift_out(40) => negative_inputs_29_40_port, 
                           shift_out(39) => negative_inputs_29_39_port, 
                           shift_out(38) => negative_inputs_29_38_port, 
                           shift_out(37) => negative_inputs_29_37_port, 
                           shift_out(36) => negative_inputs_29_36_port, 
                           shift_out(35) => negative_inputs_29_35_port, 
                           shift_out(34) => negative_inputs_29_34_port, 
                           shift_out(33) => negative_inputs_29_33_port, 
                           shift_out(32) => negative_inputs_29_32_port, 
                           shift_out(31) => negative_inputs_29_31_port, 
                           shift_out(30) => negative_inputs_29_30_port, 
                           shift_out(29) => negative_inputs_29_29_port, 
                           shift_out(28) => negative_inputs_29_28_port, 
                           shift_out(27) => negative_inputs_29_27_port, 
                           shift_out(26) => negative_inputs_29_26_port, 
                           shift_out(25) => negative_inputs_29_25_port, 
                           shift_out(24) => negative_inputs_29_24_port, 
                           shift_out(23) => negative_inputs_29_23_port, 
                           shift_out(22) => negative_inputs_29_22_port, 
                           shift_out(21) => negative_inputs_29_21_port, 
                           shift_out(20) => negative_inputs_29_20_port, 
                           shift_out(19) => negative_inputs_29_19_port, 
                           shift_out(18) => negative_inputs_29_18_port, 
                           shift_out(17) => negative_inputs_29_17_port, 
                           shift_out(16) => negative_inputs_29_16_port, 
                           shift_out(15) => negative_inputs_29_15_port, 
                           shift_out(14) => negative_inputs_29_14_port, 
                           shift_out(13) => negative_inputs_29_13_port, 
                           shift_out(12) => negative_inputs_29_12_port, 
                           shift_out(11) => negative_inputs_29_11_port, 
                           shift_out(10) => negative_inputs_29_10_port, 
                           shift_out(9) => negative_inputs_29_9_port, 
                           shift_out(8) => negative_inputs_29_8_port, 
                           shift_out(7) => negative_inputs_29_7_port, 
                           shift_out(6) => negative_inputs_29_6_port, 
                           shift_out(5) => negative_inputs_29_5_port, 
                           shift_out(4) => negative_inputs_29_4_port, 
                           shift_out(3) => negative_inputs_29_3_port, 
                           shift_out(2) => negative_inputs_29_2_port, 
                           shift_out(1) => negative_inputs_29_1_port, 
                           shift_out(0) => n_1124);
   shifted_neg_30 : leftshifter_NbitShifter64_2 port map( shift_in(63) => 
                           negative_inputs_29_63_port, shift_in(62) => 
                           negative_inputs_29_62_port, shift_in(61) => 
                           negative_inputs_29_61_port, shift_in(60) => 
                           negative_inputs_29_60_port, shift_in(59) => 
                           negative_inputs_29_59_port, shift_in(58) => 
                           negative_inputs_29_58_port, shift_in(57) => 
                           negative_inputs_29_57_port, shift_in(56) => 
                           negative_inputs_29_56_port, shift_in(55) => 
                           negative_inputs_29_55_port, shift_in(54) => 
                           negative_inputs_29_54_port, shift_in(53) => 
                           negative_inputs_29_53_port, shift_in(52) => 
                           negative_inputs_29_52_port, shift_in(51) => 
                           negative_inputs_29_51_port, shift_in(50) => 
                           negative_inputs_29_50_port, shift_in(49) => 
                           negative_inputs_29_49_port, shift_in(48) => 
                           negative_inputs_29_48_port, shift_in(47) => 
                           negative_inputs_29_47_port, shift_in(46) => 
                           negative_inputs_29_46_port, shift_in(45) => 
                           negative_inputs_29_45_port, shift_in(44) => 
                           negative_inputs_29_44_port, shift_in(43) => 
                           negative_inputs_29_43_port, shift_in(42) => 
                           negative_inputs_29_42_port, shift_in(41) => 
                           negative_inputs_29_41_port, shift_in(40) => 
                           negative_inputs_29_40_port, shift_in(39) => 
                           negative_inputs_29_39_port, shift_in(38) => 
                           negative_inputs_29_38_port, shift_in(37) => 
                           negative_inputs_29_37_port, shift_in(36) => 
                           negative_inputs_29_36_port, shift_in(35) => 
                           negative_inputs_29_35_port, shift_in(34) => 
                           negative_inputs_29_34_port, shift_in(33) => 
                           negative_inputs_29_33_port, shift_in(32) => 
                           negative_inputs_29_32_port, shift_in(31) => 
                           negative_inputs_29_31_port, shift_in(30) => 
                           negative_inputs_29_30_port, shift_in(29) => 
                           negative_inputs_29_29_port, shift_in(28) => 
                           negative_inputs_29_28_port, shift_in(27) => 
                           negative_inputs_29_27_port, shift_in(26) => 
                           negative_inputs_29_26_port, shift_in(25) => 
                           negative_inputs_29_25_port, shift_in(24) => 
                           negative_inputs_29_24_port, shift_in(23) => 
                           negative_inputs_29_23_port, shift_in(22) => 
                           negative_inputs_29_22_port, shift_in(21) => 
                           negative_inputs_29_21_port, shift_in(20) => 
                           negative_inputs_29_20_port, shift_in(19) => 
                           negative_inputs_29_19_port, shift_in(18) => 
                           negative_inputs_29_18_port, shift_in(17) => 
                           negative_inputs_29_17_port, shift_in(16) => 
                           negative_inputs_29_16_port, shift_in(15) => 
                           negative_inputs_29_15_port, shift_in(14) => 
                           negative_inputs_29_14_port, shift_in(13) => 
                           negative_inputs_29_13_port, shift_in(12) => 
                           negative_inputs_29_12_port, shift_in(11) => 
                           negative_inputs_29_11_port, shift_in(10) => 
                           negative_inputs_29_10_port, shift_in(9) => 
                           negative_inputs_29_9_port, shift_in(8) => 
                           negative_inputs_29_8_port, shift_in(7) => 
                           negative_inputs_29_7_port, shift_in(6) => 
                           negative_inputs_29_6_port, shift_in(5) => 
                           negative_inputs_29_5_port, shift_in(4) => 
                           negative_inputs_29_4_port, shift_in(3) => 
                           negative_inputs_29_3_port, shift_in(2) => 
                           negative_inputs_29_2_port, shift_in(1) => 
                           negative_inputs_29_1_port, shift_in(0) => n9, 
                           shift_out(63) => negative_inputs_30_63_port, 
                           shift_out(62) => negative_inputs_30_62_port, 
                           shift_out(61) => negative_inputs_30_61_port, 
                           shift_out(60) => negative_inputs_30_60_port, 
                           shift_out(59) => negative_inputs_30_59_port, 
                           shift_out(58) => negative_inputs_30_58_port, 
                           shift_out(57) => negative_inputs_30_57_port, 
                           shift_out(56) => negative_inputs_30_56_port, 
                           shift_out(55) => negative_inputs_30_55_port, 
                           shift_out(54) => negative_inputs_30_54_port, 
                           shift_out(53) => negative_inputs_30_53_port, 
                           shift_out(52) => negative_inputs_30_52_port, 
                           shift_out(51) => negative_inputs_30_51_port, 
                           shift_out(50) => negative_inputs_30_50_port, 
                           shift_out(49) => negative_inputs_30_49_port, 
                           shift_out(48) => negative_inputs_30_48_port, 
                           shift_out(47) => negative_inputs_30_47_port, 
                           shift_out(46) => negative_inputs_30_46_port, 
                           shift_out(45) => negative_inputs_30_45_port, 
                           shift_out(44) => negative_inputs_30_44_port, 
                           shift_out(43) => negative_inputs_30_43_port, 
                           shift_out(42) => negative_inputs_30_42_port, 
                           shift_out(41) => negative_inputs_30_41_port, 
                           shift_out(40) => negative_inputs_30_40_port, 
                           shift_out(39) => negative_inputs_30_39_port, 
                           shift_out(38) => negative_inputs_30_38_port, 
                           shift_out(37) => negative_inputs_30_37_port, 
                           shift_out(36) => negative_inputs_30_36_port, 
                           shift_out(35) => negative_inputs_30_35_port, 
                           shift_out(34) => negative_inputs_30_34_port, 
                           shift_out(33) => negative_inputs_30_33_port, 
                           shift_out(32) => negative_inputs_30_32_port, 
                           shift_out(31) => negative_inputs_30_31_port, 
                           shift_out(30) => negative_inputs_30_30_port, 
                           shift_out(29) => negative_inputs_30_29_port, 
                           shift_out(28) => negative_inputs_30_28_port, 
                           shift_out(27) => negative_inputs_30_27_port, 
                           shift_out(26) => negative_inputs_30_26_port, 
                           shift_out(25) => negative_inputs_30_25_port, 
                           shift_out(24) => negative_inputs_30_24_port, 
                           shift_out(23) => negative_inputs_30_23_port, 
                           shift_out(22) => negative_inputs_30_22_port, 
                           shift_out(21) => negative_inputs_30_21_port, 
                           shift_out(20) => negative_inputs_30_20_port, 
                           shift_out(19) => negative_inputs_30_19_port, 
                           shift_out(18) => negative_inputs_30_18_port, 
                           shift_out(17) => negative_inputs_30_17_port, 
                           shift_out(16) => negative_inputs_30_16_port, 
                           shift_out(15) => negative_inputs_30_15_port, 
                           shift_out(14) => negative_inputs_30_14_port, 
                           shift_out(13) => negative_inputs_30_13_port, 
                           shift_out(12) => negative_inputs_30_12_port, 
                           shift_out(11) => negative_inputs_30_11_port, 
                           shift_out(10) => negative_inputs_30_10_port, 
                           shift_out(9) => negative_inputs_30_9_port, 
                           shift_out(8) => negative_inputs_30_8_port, 
                           shift_out(7) => negative_inputs_30_7_port, 
                           shift_out(6) => negative_inputs_30_6_port, 
                           shift_out(5) => negative_inputs_30_5_port, 
                           shift_out(4) => negative_inputs_30_4_port, 
                           shift_out(3) => negative_inputs_30_3_port, 
                           shift_out(2) => negative_inputs_30_2_port, 
                           shift_out(1) => negative_inputs_30_1_port, 
                           shift_out(0) => n_1125);
   shifted_neg_31 : leftshifter_NbitShifter64_1 port map( shift_in(63) => 
                           negative_inputs_30_63_port, shift_in(62) => 
                           negative_inputs_30_62_port, shift_in(61) => 
                           negative_inputs_30_61_port, shift_in(60) => 
                           negative_inputs_30_60_port, shift_in(59) => 
                           negative_inputs_30_59_port, shift_in(58) => 
                           negative_inputs_30_58_port, shift_in(57) => 
                           negative_inputs_30_57_port, shift_in(56) => 
                           negative_inputs_30_56_port, shift_in(55) => 
                           negative_inputs_30_55_port, shift_in(54) => 
                           negative_inputs_30_54_port, shift_in(53) => 
                           negative_inputs_30_53_port, shift_in(52) => 
                           negative_inputs_30_52_port, shift_in(51) => 
                           negative_inputs_30_51_port, shift_in(50) => 
                           negative_inputs_30_50_port, shift_in(49) => 
                           negative_inputs_30_49_port, shift_in(48) => 
                           negative_inputs_30_48_port, shift_in(47) => 
                           negative_inputs_30_47_port, shift_in(46) => 
                           negative_inputs_30_46_port, shift_in(45) => 
                           negative_inputs_30_45_port, shift_in(44) => 
                           negative_inputs_30_44_port, shift_in(43) => 
                           negative_inputs_30_43_port, shift_in(42) => 
                           negative_inputs_30_42_port, shift_in(41) => 
                           negative_inputs_30_41_port, shift_in(40) => 
                           negative_inputs_30_40_port, shift_in(39) => 
                           negative_inputs_30_39_port, shift_in(38) => 
                           negative_inputs_30_38_port, shift_in(37) => 
                           negative_inputs_30_37_port, shift_in(36) => 
                           negative_inputs_30_36_port, shift_in(35) => 
                           negative_inputs_30_35_port, shift_in(34) => 
                           negative_inputs_30_34_port, shift_in(33) => 
                           negative_inputs_30_33_port, shift_in(32) => 
                           negative_inputs_30_32_port, shift_in(31) => 
                           negative_inputs_30_31_port, shift_in(30) => 
                           negative_inputs_30_30_port, shift_in(29) => 
                           negative_inputs_30_29_port, shift_in(28) => 
                           negative_inputs_30_28_port, shift_in(27) => 
                           negative_inputs_30_27_port, shift_in(26) => 
                           negative_inputs_30_26_port, shift_in(25) => 
                           negative_inputs_30_25_port, shift_in(24) => 
                           negative_inputs_30_24_port, shift_in(23) => 
                           negative_inputs_30_23_port, shift_in(22) => 
                           negative_inputs_30_22_port, shift_in(21) => 
                           negative_inputs_30_21_port, shift_in(20) => 
                           negative_inputs_30_20_port, shift_in(19) => 
                           negative_inputs_30_19_port, shift_in(18) => 
                           negative_inputs_30_18_port, shift_in(17) => 
                           negative_inputs_30_17_port, shift_in(16) => 
                           negative_inputs_30_16_port, shift_in(15) => 
                           negative_inputs_30_15_port, shift_in(14) => 
                           negative_inputs_30_14_port, shift_in(13) => 
                           negative_inputs_30_13_port, shift_in(12) => 
                           negative_inputs_30_12_port, shift_in(11) => 
                           negative_inputs_30_11_port, shift_in(10) => 
                           negative_inputs_30_10_port, shift_in(9) => 
                           negative_inputs_30_9_port, shift_in(8) => 
                           negative_inputs_30_8_port, shift_in(7) => 
                           negative_inputs_30_7_port, shift_in(6) => 
                           negative_inputs_30_6_port, shift_in(5) => 
                           negative_inputs_30_5_port, shift_in(4) => 
                           negative_inputs_30_4_port, shift_in(3) => 
                           negative_inputs_30_3_port, shift_in(2) => 
                           negative_inputs_30_2_port, shift_in(1) => 
                           negative_inputs_30_1_port, shift_in(0) => n9, 
                           shift_out(63) => negative_inputs_31_63_port, 
                           shift_out(62) => negative_inputs_31_62_port, 
                           shift_out(61) => negative_inputs_31_61_port, 
                           shift_out(60) => negative_inputs_31_60_port, 
                           shift_out(59) => negative_inputs_31_59_port, 
                           shift_out(58) => negative_inputs_31_58_port, 
                           shift_out(57) => negative_inputs_31_57_port, 
                           shift_out(56) => negative_inputs_31_56_port, 
                           shift_out(55) => negative_inputs_31_55_port, 
                           shift_out(54) => negative_inputs_31_54_port, 
                           shift_out(53) => negative_inputs_31_53_port, 
                           shift_out(52) => negative_inputs_31_52_port, 
                           shift_out(51) => negative_inputs_31_51_port, 
                           shift_out(50) => negative_inputs_31_50_port, 
                           shift_out(49) => negative_inputs_31_49_port, 
                           shift_out(48) => negative_inputs_31_48_port, 
                           shift_out(47) => negative_inputs_31_47_port, 
                           shift_out(46) => negative_inputs_31_46_port, 
                           shift_out(45) => negative_inputs_31_45_port, 
                           shift_out(44) => negative_inputs_31_44_port, 
                           shift_out(43) => negative_inputs_31_43_port, 
                           shift_out(42) => negative_inputs_31_42_port, 
                           shift_out(41) => negative_inputs_31_41_port, 
                           shift_out(40) => negative_inputs_31_40_port, 
                           shift_out(39) => negative_inputs_31_39_port, 
                           shift_out(38) => negative_inputs_31_38_port, 
                           shift_out(37) => negative_inputs_31_37_port, 
                           shift_out(36) => negative_inputs_31_36_port, 
                           shift_out(35) => negative_inputs_31_35_port, 
                           shift_out(34) => negative_inputs_31_34_port, 
                           shift_out(33) => negative_inputs_31_33_port, 
                           shift_out(32) => negative_inputs_31_32_port, 
                           shift_out(31) => negative_inputs_31_31_port, 
                           shift_out(30) => negative_inputs_31_30_port, 
                           shift_out(29) => negative_inputs_31_29_port, 
                           shift_out(28) => negative_inputs_31_28_port, 
                           shift_out(27) => negative_inputs_31_27_port, 
                           shift_out(26) => negative_inputs_31_26_port, 
                           shift_out(25) => negative_inputs_31_25_port, 
                           shift_out(24) => negative_inputs_31_24_port, 
                           shift_out(23) => negative_inputs_31_23_port, 
                           shift_out(22) => negative_inputs_31_22_port, 
                           shift_out(21) => negative_inputs_31_21_port, 
                           shift_out(20) => negative_inputs_31_20_port, 
                           shift_out(19) => negative_inputs_31_19_port, 
                           shift_out(18) => negative_inputs_31_18_port, 
                           shift_out(17) => negative_inputs_31_17_port, 
                           shift_out(16) => negative_inputs_31_16_port, 
                           shift_out(15) => negative_inputs_31_15_port, 
                           shift_out(14) => negative_inputs_31_14_port, 
                           shift_out(13) => negative_inputs_31_13_port, 
                           shift_out(12) => negative_inputs_31_12_port, 
                           shift_out(11) => negative_inputs_31_11_port, 
                           shift_out(10) => negative_inputs_31_10_port, 
                           shift_out(9) => negative_inputs_31_9_port, 
                           shift_out(8) => negative_inputs_31_8_port, 
                           shift_out(7) => negative_inputs_31_7_port, 
                           shift_out(6) => negative_inputs_31_6_port, 
                           shift_out(5) => negative_inputs_31_5_port, 
                           shift_out(4) => negative_inputs_31_4_port, 
                           shift_out(3) => negative_inputs_31_3_port, 
                           shift_out(2) => negative_inputs_31_2_port, 
                           shift_out(1) => negative_inputs_31_1_port, 
                           shift_out(0) => n_1126);
   encoder0_0 : encoder_0 port map( pieceofB(2) => B(1), pieceofB(1) => B(0), 
                           pieceofB(0) => X_Logic0_port, sel(2) => sel_0_2_port
                           , sel(1) => sel_0_1_port, sel(0) => sel_0_0_port);
   MUX0_0 : MUX51_MuxNbit64_0 port map( zeroSignal(63) => X_Logic0_port, 
                           zeroSignal(62) => X_Logic0_port, zeroSignal(61) => 
                           X_Logic0_port, zeroSignal(60) => X_Logic0_port, 
                           zeroSignal(59) => X_Logic0_port, zeroSignal(58) => 
                           X_Logic0_port, zeroSignal(57) => X_Logic0_port, 
                           zeroSignal(56) => X_Logic0_port, zeroSignal(55) => 
                           X_Logic0_port, zeroSignal(54) => X_Logic0_port, 
                           zeroSignal(53) => X_Logic0_port, zeroSignal(52) => 
                           X_Logic0_port, zeroSignal(51) => X_Logic0_port, 
                           zeroSignal(50) => X_Logic0_port, zeroSignal(49) => 
                           X_Logic0_port, zeroSignal(48) => X_Logic0_port, 
                           zeroSignal(47) => X_Logic0_port, zeroSignal(46) => 
                           X_Logic0_port, zeroSignal(45) => X_Logic0_port, 
                           zeroSignal(44) => X_Logic0_port, zeroSignal(43) => 
                           X_Logic0_port, zeroSignal(42) => X_Logic0_port, 
                           zeroSignal(41) => X_Logic0_port, zeroSignal(40) => 
                           X_Logic0_port, zeroSignal(39) => X_Logic0_port, 
                           zeroSignal(38) => X_Logic0_port, zeroSignal(37) => 
                           X_Logic0_port, zeroSignal(36) => X_Logic0_port, 
                           zeroSignal(35) => X_Logic0_port, zeroSignal(34) => 
                           X_Logic0_port, zeroSignal(33) => X_Logic0_port, 
                           zeroSignal(32) => X_Logic0_port, zeroSignal(31) => 
                           X_Logic0_port, zeroSignal(30) => X_Logic0_port, 
                           zeroSignal(29) => X_Logic0_port, zeroSignal(28) => 
                           X_Logic0_port, zeroSignal(27) => X_Logic0_port, 
                           zeroSignal(26) => X_Logic0_port, zeroSignal(25) => 
                           X_Logic0_port, zeroSignal(24) => X_Logic0_port, 
                           zeroSignal(23) => X_Logic0_port, zeroSignal(22) => 
                           X_Logic0_port, zeroSignal(21) => X_Logic0_port, 
                           zeroSignal(20) => X_Logic0_port, zeroSignal(19) => 
                           X_Logic0_port, zeroSignal(18) => X_Logic0_port, 
                           zeroSignal(17) => X_Logic0_port, zeroSignal(16) => 
                           X_Logic0_port, zeroSignal(15) => X_Logic0_port, 
                           zeroSignal(14) => X_Logic0_port, zeroSignal(13) => 
                           X_Logic0_port, zeroSignal(12) => X_Logic0_port, 
                           zeroSignal(11) => X_Logic0_port, zeroSignal(10) => 
                           X_Logic0_port, zeroSignal(9) => X_Logic0_port, 
                           zeroSignal(8) => X_Logic0_port, zeroSignal(7) => 
                           X_Logic0_port, zeroSignal(6) => X_Logic0_port, 
                           zeroSignal(5) => X_Logic0_port, zeroSignal(4) => 
                           X_Logic0_port, zeroSignal(3) => X_Logic0_port, 
                           zeroSignal(2) => X_Logic0_port, zeroSignal(1) => 
                           X_Logic0_port, zeroSignal(0) => X_Logic0_port, 
                           A_signal(63) => A(31), A_signal(62) => A(31), 
                           A_signal(61) => A(31), A_signal(60) => A(31), 
                           A_signal(59) => A(31), A_signal(58) => A(31), 
                           A_signal(57) => A(31), A_signal(56) => A(31), 
                           A_signal(55) => A(31), A_signal(54) => A(31), 
                           A_signal(53) => A(31), A_signal(52) => A(31), 
                           A_signal(51) => A(31), A_signal(50) => A(31), 
                           A_signal(49) => A(31), A_signal(48) => A(31), 
                           A_signal(47) => A(31), A_signal(46) => A(31), 
                           A_signal(45) => A(31), A_signal(44) => A(31), 
                           A_signal(43) => A(31), A_signal(42) => A(31), 
                           A_signal(41) => A(31), A_signal(40) => A(31), 
                           A_signal(39) => A(31), A_signal(38) => A(31), 
                           A_signal(37) => A(31), A_signal(36) => A(31), 
                           A_signal(35) => A(31), A_signal(34) => A(31), 
                           A_signal(33) => A(31), A_signal(32) => A(31), 
                           A_signal(31) => A(31), A_signal(30) => A(30), 
                           A_signal(29) => A(29), A_signal(28) => A(28), 
                           A_signal(27) => A(27), A_signal(26) => A(26), 
                           A_signal(25) => A(25), A_signal(24) => A(24), 
                           A_signal(23) => A(23), A_signal(22) => A(22), 
                           A_signal(21) => A(21), A_signal(20) => A(20), 
                           A_signal(19) => A(19), A_signal(18) => A(18), 
                           A_signal(17) => A(17), A_signal(16) => A(16), 
                           A_signal(15) => A(15), A_signal(14) => A(14), 
                           A_signal(13) => A(13), A_signal(12) => A(12), 
                           A_signal(11) => A(11), A_signal(10) => A(10), 
                           A_signal(9) => A(9), A_signal(8) => A(8), 
                           A_signal(7) => A(7), A_signal(6) => A(6), 
                           A_signal(5) => A(5), A_signal(4) => A(4), 
                           A_signal(3) => A(3), A_signal(2) => A(2), 
                           A_signal(1) => n11, A_signal(0) => n72, A_neg(63) =>
                           negative_inputs_0_63_port, A_neg(62) => 
                           negative_inputs_0_62_port, A_neg(61) => 
                           negative_inputs_0_61_port, A_neg(60) => 
                           negative_inputs_0_60_port, A_neg(59) => 
                           negative_inputs_0_59_port, A_neg(58) => 
                           negative_inputs_0_58_port, A_neg(57) => 
                           negative_inputs_0_57_port, A_neg(56) => 
                           negative_inputs_0_56_port, A_neg(55) => 
                           negative_inputs_0_55_port, A_neg(54) => 
                           negative_inputs_0_54_port, A_neg(53) => 
                           negative_inputs_0_53_port, A_neg(52) => 
                           negative_inputs_0_52_port, A_neg(51) => 
                           negative_inputs_0_51_port, A_neg(50) => 
                           negative_inputs_0_50_port, A_neg(49) => 
                           negative_inputs_0_49_port, A_neg(48) => 
                           negative_inputs_0_48_port, A_neg(47) => 
                           negative_inputs_0_47_port, A_neg(46) => 
                           negative_inputs_0_46_port, A_neg(45) => 
                           negative_inputs_0_45_port, A_neg(44) => 
                           negative_inputs_0_44_port, A_neg(43) => 
                           negative_inputs_0_43_port, A_neg(42) => 
                           negative_inputs_0_42_port, A_neg(41) => 
                           negative_inputs_0_41_port, A_neg(40) => 
                           negative_inputs_0_40_port, A_neg(39) => 
                           negative_inputs_0_39_port, A_neg(38) => 
                           negative_inputs_0_38_port, A_neg(37) => 
                           negative_inputs_0_37_port, A_neg(36) => 
                           negative_inputs_0_36_port, A_neg(35) => 
                           negative_inputs_0_35_port, A_neg(34) => 
                           negative_inputs_0_34_port, A_neg(33) => 
                           negative_inputs_0_33_port, A_neg(32) => 
                           negative_inputs_0_32_port, A_neg(31) => 
                           negative_inputs_0_31_port, A_neg(30) => 
                           negative_inputs_0_30_port, A_neg(29) => 
                           negative_inputs_0_29_port, A_neg(28) => 
                           negative_inputs_0_28_port, A_neg(27) => 
                           negative_inputs_0_27_port, A_neg(26) => 
                           negative_inputs_0_26_port, A_neg(25) => 
                           negative_inputs_0_25_port, A_neg(24) => 
                           negative_inputs_0_24_port, A_neg(23) => 
                           negative_inputs_0_23_port, A_neg(22) => 
                           negative_inputs_0_22_port, A_neg(21) => 
                           negative_inputs_0_21_port, A_neg(20) => 
                           negative_inputs_0_20_port, A_neg(19) => 
                           negative_inputs_0_19_port, A_neg(18) => 
                           negative_inputs_0_18_port, A_neg(17) => 
                           negative_inputs_0_17_port, A_neg(16) => 
                           negative_inputs_0_16_port, A_neg(15) => 
                           negative_inputs_0_15_port, A_neg(14) => 
                           negative_inputs_0_14_port, A_neg(13) => 
                           negative_inputs_0_13_port, A_neg(12) => 
                           negative_inputs_0_12_port, A_neg(11) => 
                           negative_inputs_0_11_port, A_neg(10) => 
                           negative_inputs_0_10_port, A_neg(9) => 
                           negative_inputs_0_9_port, A_neg(8) => 
                           negative_inputs_0_8_port, A_neg(7) => 
                           negative_inputs_0_7_port, A_neg(6) => 
                           negative_inputs_0_6_port, A_neg(5) => 
                           negative_inputs_0_5_port, A_neg(4) => 
                           negative_inputs_0_4_port, A_neg(3) => 
                           negative_inputs_0_3_port, A_neg(2) => 
                           negative_inputs_0_2_port, A_neg(1) => 
                           negative_inputs_0_1_port, A_neg(0) => 
                           negative_inputs_0_0_port, A_shifted(63) => 
                           positive_inputs_1_63_port, A_shifted(62) => 
                           positive_inputs_1_62_port, A_shifted(61) => 
                           positive_inputs_1_61_port, A_shifted(60) => 
                           positive_inputs_1_60_port, A_shifted(59) => 
                           positive_inputs_1_59_port, A_shifted(58) => 
                           positive_inputs_1_58_port, A_shifted(57) => 
                           positive_inputs_1_57_port, A_shifted(56) => 
                           positive_inputs_1_56_port, A_shifted(55) => 
                           positive_inputs_1_55_port, A_shifted(54) => 
                           positive_inputs_1_54_port, A_shifted(53) => 
                           positive_inputs_1_53_port, A_shifted(52) => 
                           positive_inputs_1_52_port, A_shifted(51) => 
                           positive_inputs_1_51_port, A_shifted(50) => 
                           positive_inputs_1_50_port, A_shifted(49) => 
                           positive_inputs_1_49_port, A_shifted(48) => n70, 
                           A_shifted(47) => positive_inputs_1_47_port, 
                           A_shifted(46) => positive_inputs_1_46_port, 
                           A_shifted(45) => positive_inputs_1_45_port, 
                           A_shifted(44) => positive_inputs_1_44_port, 
                           A_shifted(43) => positive_inputs_1_43_port, 
                           A_shifted(42) => positive_inputs_1_42_port, 
                           A_shifted(41) => positive_inputs_1_41_port, 
                           A_shifted(40) => positive_inputs_1_40_port, 
                           A_shifted(39) => positive_inputs_1_39_port, 
                           A_shifted(38) => n50, A_shifted(37) => 
                           positive_inputs_1_37_port, A_shifted(36) => 
                           positive_inputs_1_36_port, A_shifted(35) => 
                           positive_inputs_1_35_port, A_shifted(34) => 
                           positive_inputs_1_34_port, A_shifted(33) => 
                           positive_inputs_1_33_port, A_shifted(32) => 
                           positive_inputs_1_32_port, A_shifted(31) => 
                           positive_inputs_1_31_port, A_shifted(30) => 
                           positive_inputs_1_30_port, A_shifted(29) => 
                           positive_inputs_1_29_port, A_shifted(28) => 
                           positive_inputs_1_28_port, A_shifted(27) => 
                           positive_inputs_1_27_port, A_shifted(26) => 
                           positive_inputs_1_26_port, A_shifted(25) => 
                           positive_inputs_1_25_port, A_shifted(24) => 
                           positive_inputs_1_24_port, A_shifted(23) => 
                           positive_inputs_1_23_port, A_shifted(22) => 
                           positive_inputs_1_22_port, A_shifted(21) => 
                           positive_inputs_1_21_port, A_shifted(20) => 
                           positive_inputs_1_20_port, A_shifted(19) => 
                           positive_inputs_1_19_port, A_shifted(18) => 
                           positive_inputs_1_18_port, A_shifted(17) => 
                           positive_inputs_1_17_port, A_shifted(16) => 
                           positive_inputs_1_16_port, A_shifted(15) => 
                           positive_inputs_1_15_port, A_shifted(14) => 
                           positive_inputs_1_14_port, A_shifted(13) => 
                           positive_inputs_1_13_port, A_shifted(12) => 
                           positive_inputs_1_12_port, A_shifted(11) => 
                           positive_inputs_1_11_port, A_shifted(10) => 
                           positive_inputs_1_10_port, A_shifted(9) => 
                           positive_inputs_1_9_port, A_shifted(8) => 
                           positive_inputs_1_8_port, A_shifted(7) => 
                           positive_inputs_1_7_port, A_shifted(6) => 
                           positive_inputs_1_6_port, A_shifted(5) => 
                           positive_inputs_1_5_port, A_shifted(4) => 
                           positive_inputs_1_4_port, A_shifted(3) => 
                           positive_inputs_1_3_port, A_shifted(2) => 
                           positive_inputs_1_2_port, A_shifted(1) => 
                           positive_inputs_1_1_port, A_shifted(0) => n9, 
                           A_neg_shifted(63) => negative_inputs_1_63_port, 
                           A_neg_shifted(62) => negative_inputs_1_62_port, 
                           A_neg_shifted(61) => negative_inputs_1_61_port, 
                           A_neg_shifted(60) => negative_inputs_1_60_port, 
                           A_neg_shifted(59) => negative_inputs_1_59_port, 
                           A_neg_shifted(58) => negative_inputs_1_58_port, 
                           A_neg_shifted(57) => negative_inputs_1_57_port, 
                           A_neg_shifted(56) => negative_inputs_1_56_port, 
                           A_neg_shifted(55) => negative_inputs_1_55_port, 
                           A_neg_shifted(54) => negative_inputs_1_54_port, 
                           A_neg_shifted(53) => negative_inputs_1_53_port, 
                           A_neg_shifted(52) => negative_inputs_1_52_port, 
                           A_neg_shifted(51) => negative_inputs_1_51_port, 
                           A_neg_shifted(50) => negative_inputs_1_50_port, 
                           A_neg_shifted(49) => negative_inputs_1_49_port, 
                           A_neg_shifted(48) => negative_inputs_1_48_port, 
                           A_neg_shifted(47) => negative_inputs_1_47_port, 
                           A_neg_shifted(46) => negative_inputs_1_46_port, 
                           A_neg_shifted(45) => negative_inputs_1_45_port, 
                           A_neg_shifted(44) => negative_inputs_1_44_port, 
                           A_neg_shifted(43) => negative_inputs_1_43_port, 
                           A_neg_shifted(42) => negative_inputs_1_42_port, 
                           A_neg_shifted(41) => negative_inputs_1_41_port, 
                           A_neg_shifted(40) => negative_inputs_1_40_port, 
                           A_neg_shifted(39) => n149, A_neg_shifted(38) => 
                           negative_inputs_1_38_port, A_neg_shifted(37) => 
                           negative_inputs_1_37_port, A_neg_shifted(36) => 
                           negative_inputs_1_36_port, A_neg_shifted(35) => 
                           negative_inputs_1_35_port, A_neg_shifted(34) => 
                           negative_inputs_1_34_port, A_neg_shifted(33) => 
                           negative_inputs_1_33_port, A_neg_shifted(32) => 
                           negative_inputs_1_32_port, A_neg_shifted(31) => 
                           negative_inputs_1_31_port, A_neg_shifted(30) => 
                           negative_inputs_1_30_port, A_neg_shifted(29) => 
                           negative_inputs_1_29_port, A_neg_shifted(28) => 
                           negative_inputs_1_28_port, A_neg_shifted(27) => 
                           negative_inputs_1_27_port, A_neg_shifted(26) => 
                           negative_inputs_1_26_port, A_neg_shifted(25) => 
                           negative_inputs_1_25_port, A_neg_shifted(24) => 
                           negative_inputs_1_24_port, A_neg_shifted(23) => 
                           negative_inputs_1_23_port, A_neg_shifted(22) => 
                           negative_inputs_1_22_port, A_neg_shifted(21) => 
                           negative_inputs_1_21_port, A_neg_shifted(20) => 
                           negative_inputs_1_20_port, A_neg_shifted(19) => 
                           negative_inputs_1_19_port, A_neg_shifted(18) => 
                           negative_inputs_1_18_port, A_neg_shifted(17) => 
                           negative_inputs_1_17_port, A_neg_shifted(16) => 
                           negative_inputs_1_16_port, A_neg_shifted(15) => 
                           negative_inputs_1_15_port, A_neg_shifted(14) => 
                           negative_inputs_1_14_port, A_neg_shifted(13) => 
                           negative_inputs_1_13_port, A_neg_shifted(12) => 
                           negative_inputs_1_12_port, A_neg_shifted(11) => 
                           negative_inputs_1_11_port, A_neg_shifted(10) => 
                           negative_inputs_1_10_port, A_neg_shifted(9) => 
                           negative_inputs_1_9_port, A_neg_shifted(8) => 
                           negative_inputs_1_8_port, A_neg_shifted(7) => 
                           negative_inputs_1_7_port, A_neg_shifted(6) => 
                           negative_inputs_1_6_port, A_neg_shifted(5) => 
                           negative_inputs_1_5_port, A_neg_shifted(4) => 
                           negative_inputs_1_4_port, A_neg_shifted(3) => 
                           negative_inputs_1_3_port, A_neg_shifted(2) => 
                           negative_inputs_1_2_port, A_neg_shifted(1) => 
                           negative_inputs_1_1_port, A_neg_shifted(0) => n9, 
                           Sel(2) => sel_0_2_port, Sel(1) => sel_0_1_port, 
                           Sel(0) => sel_0_0_port, Y(63) => 
                           MuxOutputs_0_63_port, Y(62) => MuxOutputs_0_62_port,
                           Y(61) => MuxOutputs_0_61_port, Y(60) => 
                           MuxOutputs_0_60_port, Y(59) => MuxOutputs_0_59_port,
                           Y(58) => MuxOutputs_0_58_port, Y(57) => 
                           MuxOutputs_0_57_port, Y(56) => MuxOutputs_0_56_port,
                           Y(55) => MuxOutputs_0_55_port, Y(54) => 
                           MuxOutputs_0_54_port, Y(53) => MuxOutputs_0_53_port,
                           Y(52) => MuxOutputs_0_52_port, Y(51) => 
                           MuxOutputs_0_51_port, Y(50) => MuxOutputs_0_50_port,
                           Y(49) => MuxOutputs_0_49_port, Y(48) => 
                           MuxOutputs_0_48_port, Y(47) => MuxOutputs_0_47_port,
                           Y(46) => MuxOutputs_0_46_port, Y(45) => 
                           MuxOutputs_0_45_port, Y(44) => MuxOutputs_0_44_port,
                           Y(43) => MuxOutputs_0_43_port, Y(42) => 
                           MuxOutputs_0_42_port, Y(41) => MuxOutputs_0_41_port,
                           Y(40) => MuxOutputs_0_40_port, Y(39) => 
                           MuxOutputs_0_39_port, Y(38) => MuxOutputs_0_38_port,
                           Y(37) => MuxOutputs_0_37_port, Y(36) => 
                           MuxOutputs_0_36_port, Y(35) => MuxOutputs_0_35_port,
                           Y(34) => MuxOutputs_0_34_port, Y(33) => 
                           MuxOutputs_0_33_port, Y(32) => MuxOutputs_0_32_port,
                           Y(31) => MuxOutputs_0_31_port, Y(30) => 
                           MuxOutputs_0_30_port, Y(29) => MuxOutputs_0_29_port,
                           Y(28) => MuxOutputs_0_28_port, Y(27) => 
                           MuxOutputs_0_27_port, Y(26) => MuxOutputs_0_26_port,
                           Y(25) => MuxOutputs_0_25_port, Y(24) => 
                           MuxOutputs_0_24_port, Y(23) => MuxOutputs_0_23_port,
                           Y(22) => MuxOutputs_0_22_port, Y(21) => 
                           MuxOutputs_0_21_port, Y(20) => MuxOutputs_0_20_port,
                           Y(19) => MuxOutputs_0_19_port, Y(18) => 
                           MuxOutputs_0_18_port, Y(17) => MuxOutputs_0_17_port,
                           Y(16) => MuxOutputs_0_16_port, Y(15) => 
                           MuxOutputs_0_15_port, Y(14) => MuxOutputs_0_14_port,
                           Y(13) => MuxOutputs_0_13_port, Y(12) => 
                           MuxOutputs_0_12_port, Y(11) => MuxOutputs_0_11_port,
                           Y(10) => MuxOutputs_0_10_port, Y(9) => 
                           MuxOutputs_0_9_port, Y(8) => MuxOutputs_0_8_port, 
                           Y(7) => MuxOutputs_0_7_port, Y(6) => 
                           MuxOutputs_0_6_port, Y(5) => MuxOutputs_0_5_port, 
                           Y(4) => MuxOutputs_0_4_port, Y(3) => 
                           MuxOutputs_0_3_port, Y(2) => MuxOutputs_0_2_port, 
                           Y(1) => MuxOutputs_0_1_port, Y(0) => 
                           MuxOutputs_0_0_port);
   encoderI_1 : encoder_15 port map( pieceofB(2) => B(3), pieceofB(1) => B(2), 
                           pieceofB(0) => B(1), sel(2) => sel_1_2_port, sel(1) 
                           => sel_1_1_port, sel(0) => sel_1_0_port);
   MUXI_1 : MUX51_MuxNbit64_15 port map( zeroSignal(63) => X_Logic0_port, 
                           zeroSignal(62) => X_Logic0_port, zeroSignal(61) => 
                           X_Logic0_port, zeroSignal(60) => X_Logic0_port, 
                           zeroSignal(59) => X_Logic0_port, zeroSignal(58) => 
                           X_Logic0_port, zeroSignal(57) => X_Logic0_port, 
                           zeroSignal(56) => X_Logic0_port, zeroSignal(55) => 
                           X_Logic0_port, zeroSignal(54) => X_Logic0_port, 
                           zeroSignal(53) => X_Logic0_port, zeroSignal(52) => 
                           X_Logic0_port, zeroSignal(51) => X_Logic0_port, 
                           zeroSignal(50) => X_Logic0_port, zeroSignal(49) => 
                           X_Logic0_port, zeroSignal(48) => X_Logic0_port, 
                           zeroSignal(47) => X_Logic0_port, zeroSignal(46) => 
                           X_Logic0_port, zeroSignal(45) => X_Logic0_port, 
                           zeroSignal(44) => X_Logic0_port, zeroSignal(43) => 
                           X_Logic0_port, zeroSignal(42) => X_Logic0_port, 
                           zeroSignal(41) => X_Logic0_port, zeroSignal(40) => 
                           X_Logic0_port, zeroSignal(39) => X_Logic0_port, 
                           zeroSignal(38) => X_Logic0_port, zeroSignal(37) => 
                           X_Logic0_port, zeroSignal(36) => X_Logic0_port, 
                           zeroSignal(35) => X_Logic0_port, zeroSignal(34) => 
                           X_Logic0_port, zeroSignal(33) => X_Logic0_port, 
                           zeroSignal(32) => X_Logic0_port, zeroSignal(31) => 
                           X_Logic0_port, zeroSignal(30) => X_Logic0_port, 
                           zeroSignal(29) => X_Logic0_port, zeroSignal(28) => 
                           X_Logic0_port, zeroSignal(27) => X_Logic0_port, 
                           zeroSignal(26) => X_Logic0_port, zeroSignal(25) => 
                           X_Logic0_port, zeroSignal(24) => X_Logic0_port, 
                           zeroSignal(23) => X_Logic0_port, zeroSignal(22) => 
                           X_Logic0_port, zeroSignal(21) => X_Logic0_port, 
                           zeroSignal(20) => X_Logic0_port, zeroSignal(19) => 
                           X_Logic0_port, zeroSignal(18) => X_Logic0_port, 
                           zeroSignal(17) => X_Logic0_port, zeroSignal(16) => 
                           X_Logic0_port, zeroSignal(15) => X_Logic0_port, 
                           zeroSignal(14) => X_Logic0_port, zeroSignal(13) => 
                           X_Logic0_port, zeroSignal(12) => X_Logic0_port, 
                           zeroSignal(11) => X_Logic0_port, zeroSignal(10) => 
                           X_Logic0_port, zeroSignal(9) => X_Logic0_port, 
                           zeroSignal(8) => X_Logic0_port, zeroSignal(7) => 
                           X_Logic0_port, zeroSignal(6) => X_Logic0_port, 
                           zeroSignal(5) => X_Logic0_port, zeroSignal(4) => 
                           X_Logic0_port, zeroSignal(3) => X_Logic0_port, 
                           zeroSignal(2) => X_Logic0_port, zeroSignal(1) => 
                           X_Logic0_port, zeroSignal(0) => X_Logic0_port, 
                           A_signal(63) => positive_inputs_2_63_port, 
                           A_signal(62) => positive_inputs_2_62_port, 
                           A_signal(61) => positive_inputs_2_61_port, 
                           A_signal(60) => positive_inputs_2_60_port, 
                           A_signal(59) => positive_inputs_2_59_port, 
                           A_signal(58) => positive_inputs_2_58_port, 
                           A_signal(57) => positive_inputs_2_57_port, 
                           A_signal(56) => positive_inputs_2_56_port, 
                           A_signal(55) => positive_inputs_2_55_port, 
                           A_signal(54) => positive_inputs_2_54_port, 
                           A_signal(53) => positive_inputs_2_53_port, 
                           A_signal(52) => positive_inputs_2_52_port, 
                           A_signal(51) => positive_inputs_2_51_port, 
                           A_signal(50) => positive_inputs_2_50_port, 
                           A_signal(49) => positive_inputs_2_49_port, 
                           A_signal(48) => n69, A_signal(47) => 
                           positive_inputs_2_47_port, A_signal(46) => 
                           positive_inputs_2_46_port, A_signal(45) => 
                           positive_inputs_2_45_port, A_signal(44) => 
                           positive_inputs_2_44_port, A_signal(43) => 
                           positive_inputs_2_43_port, A_signal(42) => 
                           positive_inputs_2_42_port, A_signal(41) => 
                           positive_inputs_2_41_port, A_signal(40) => 
                           positive_inputs_2_40_port, A_signal(39) => 
                           positive_inputs_2_39_port, A_signal(38) => n49, 
                           A_signal(37) => positive_inputs_2_37_port, 
                           A_signal(36) => positive_inputs_2_36_port, 
                           A_signal(35) => positive_inputs_2_35_port, 
                           A_signal(34) => positive_inputs_2_34_port, 
                           A_signal(33) => positive_inputs_2_33_port, 
                           A_signal(32) => positive_inputs_2_32_port, 
                           A_signal(31) => positive_inputs_2_31_port, 
                           A_signal(30) => positive_inputs_2_30_port, 
                           A_signal(29) => positive_inputs_2_29_port, 
                           A_signal(28) => positive_inputs_2_28_port, 
                           A_signal(27) => positive_inputs_2_27_port, 
                           A_signal(26) => positive_inputs_2_26_port, 
                           A_signal(25) => positive_inputs_2_25_port, 
                           A_signal(24) => positive_inputs_2_24_port, 
                           A_signal(23) => positive_inputs_2_23_port, 
                           A_signal(22) => positive_inputs_2_22_port, 
                           A_signal(21) => positive_inputs_2_21_port, 
                           A_signal(20) => positive_inputs_2_20_port, 
                           A_signal(19) => positive_inputs_2_19_port, 
                           A_signal(18) => positive_inputs_2_18_port, 
                           A_signal(17) => positive_inputs_2_17_port, 
                           A_signal(16) => positive_inputs_2_16_port, 
                           A_signal(15) => positive_inputs_2_15_port, 
                           A_signal(14) => positive_inputs_2_14_port, 
                           A_signal(13) => positive_inputs_2_13_port, 
                           A_signal(12) => positive_inputs_2_12_port, 
                           A_signal(11) => positive_inputs_2_11_port, 
                           A_signal(10) => positive_inputs_2_10_port, 
                           A_signal(9) => positive_inputs_2_9_port, A_signal(8)
                           => positive_inputs_2_8_port, A_signal(7) => 
                           positive_inputs_2_7_port, A_signal(6) => 
                           positive_inputs_2_6_port, A_signal(5) => 
                           positive_inputs_2_5_port, A_signal(4) => 
                           positive_inputs_2_4_port, A_signal(3) => 
                           positive_inputs_2_3_port, A_signal(2) => 
                           positive_inputs_2_2_port, A_signal(1) => 
                           positive_inputs_2_1_port, A_signal(0) => n9, 
                           A_neg(63) => negative_inputs_2_63_port, A_neg(62) =>
                           negative_inputs_2_62_port, A_neg(61) => 
                           negative_inputs_2_61_port, A_neg(60) => 
                           negative_inputs_2_60_port, A_neg(59) => 
                           negative_inputs_2_59_port, A_neg(58) => 
                           negative_inputs_2_58_port, A_neg(57) => 
                           negative_inputs_2_57_port, A_neg(56) => 
                           negative_inputs_2_56_port, A_neg(55) => 
                           negative_inputs_2_55_port, A_neg(54) => 
                           negative_inputs_2_54_port, A_neg(53) => 
                           negative_inputs_2_53_port, A_neg(52) => 
                           negative_inputs_2_52_port, A_neg(51) => 
                           negative_inputs_2_51_port, A_neg(50) => 
                           negative_inputs_2_50_port, A_neg(49) => 
                           negative_inputs_2_49_port, A_neg(48) => 
                           negative_inputs_2_48_port, A_neg(47) => 
                           negative_inputs_2_47_port, A_neg(46) => 
                           negative_inputs_2_46_port, A_neg(45) => 
                           negative_inputs_2_45_port, A_neg(44) => 
                           negative_inputs_2_44_port, A_neg(43) => 
                           negative_inputs_2_43_port, A_neg(42) => 
                           negative_inputs_2_42_port, A_neg(41) => 
                           negative_inputs_2_41_port, A_neg(40) => 
                           negative_inputs_2_40_port, A_neg(39) => n147, 
                           A_neg(38) => negative_inputs_2_38_port, A_neg(37) =>
                           negative_inputs_2_37_port, A_neg(36) => 
                           negative_inputs_2_36_port, A_neg(35) => 
                           negative_inputs_2_35_port, A_neg(34) => 
                           negative_inputs_2_34_port, A_neg(33) => 
                           negative_inputs_2_33_port, A_neg(32) => 
                           negative_inputs_2_32_port, A_neg(31) => 
                           negative_inputs_2_31_port, A_neg(30) => 
                           negative_inputs_2_30_port, A_neg(29) => 
                           negative_inputs_2_29_port, A_neg(28) => 
                           negative_inputs_2_28_port, A_neg(27) => 
                           negative_inputs_2_27_port, A_neg(26) => 
                           negative_inputs_2_26_port, A_neg(25) => 
                           negative_inputs_2_25_port, A_neg(24) => 
                           negative_inputs_2_24_port, A_neg(23) => 
                           negative_inputs_2_23_port, A_neg(22) => 
                           negative_inputs_2_22_port, A_neg(21) => 
                           negative_inputs_2_21_port, A_neg(20) => 
                           negative_inputs_2_20_port, A_neg(19) => 
                           negative_inputs_2_19_port, A_neg(18) => 
                           negative_inputs_2_18_port, A_neg(17) => 
                           negative_inputs_2_17_port, A_neg(16) => 
                           negative_inputs_2_16_port, A_neg(15) => 
                           negative_inputs_2_15_port, A_neg(14) => 
                           negative_inputs_2_14_port, A_neg(13) => 
                           negative_inputs_2_13_port, A_neg(12) => 
                           negative_inputs_2_12_port, A_neg(11) => 
                           negative_inputs_2_11_port, A_neg(10) => 
                           negative_inputs_2_10_port, A_neg(9) => 
                           negative_inputs_2_9_port, A_neg(8) => 
                           negative_inputs_2_8_port, A_neg(7) => 
                           negative_inputs_2_7_port, A_neg(6) => 
                           negative_inputs_2_6_port, A_neg(5) => 
                           negative_inputs_2_5_port, A_neg(4) => 
                           negative_inputs_2_4_port, A_neg(3) => 
                           negative_inputs_2_3_port, A_neg(2) => 
                           negative_inputs_2_2_port, A_neg(1) => 
                           negative_inputs_2_1_port, A_neg(0) => n9, 
                           A_shifted(63) => positive_inputs_3_63_port, 
                           A_shifted(62) => positive_inputs_3_62_port, 
                           A_shifted(61) => positive_inputs_3_61_port, 
                           A_shifted(60) => positive_inputs_3_60_port, 
                           A_shifted(59) => positive_inputs_3_59_port, 
                           A_shifted(58) => positive_inputs_3_58_port, 
                           A_shifted(57) => positive_inputs_3_57_port, 
                           A_shifted(56) => positive_inputs_3_56_port, 
                           A_shifted(55) => positive_inputs_3_55_port, 
                           A_shifted(54) => positive_inputs_3_54_port, 
                           A_shifted(53) => positive_inputs_3_53_port, 
                           A_shifted(52) => positive_inputs_3_52_port, 
                           A_shifted(51) => positive_inputs_3_51_port, 
                           A_shifted(50) => positive_inputs_3_50_port, 
                           A_shifted(49) => positive_inputs_3_49_port, 
                           A_shifted(48) => positive_inputs_3_48_port, 
                           A_shifted(47) => positive_inputs_3_47_port, 
                           A_shifted(46) => positive_inputs_3_46_port, 
                           A_shifted(45) => positive_inputs_3_45_port, 
                           A_shifted(44) => positive_inputs_3_44_port, 
                           A_shifted(43) => positive_inputs_3_43_port, 
                           A_shifted(42) => positive_inputs_3_42_port, 
                           A_shifted(41) => positive_inputs_3_41_port, 
                           A_shifted(40) => positive_inputs_3_40_port, 
                           A_shifted(39) => positive_inputs_3_39_port, 
                           A_shifted(38) => positive_inputs_3_38_port, 
                           A_shifted(37) => positive_inputs_3_37_port, 
                           A_shifted(36) => positive_inputs_3_36_port, 
                           A_shifted(35) => positive_inputs_3_35_port, 
                           A_shifted(34) => positive_inputs_3_34_port, 
                           A_shifted(33) => positive_inputs_3_33_port, 
                           A_shifted(32) => positive_inputs_3_32_port, 
                           A_shifted(31) => positive_inputs_3_31_port, 
                           A_shifted(30) => positive_inputs_3_30_port, 
                           A_shifted(29) => positive_inputs_3_29_port, 
                           A_shifted(28) => positive_inputs_3_28_port, 
                           A_shifted(27) => positive_inputs_3_27_port, 
                           A_shifted(26) => positive_inputs_3_26_port, 
                           A_shifted(25) => positive_inputs_3_25_port, 
                           A_shifted(24) => positive_inputs_3_24_port, 
                           A_shifted(23) => positive_inputs_3_23_port, 
                           A_shifted(22) => positive_inputs_3_22_port, 
                           A_shifted(21) => positive_inputs_3_21_port, 
                           A_shifted(20) => positive_inputs_3_20_port, 
                           A_shifted(19) => positive_inputs_3_19_port, 
                           A_shifted(18) => positive_inputs_3_18_port, 
                           A_shifted(17) => positive_inputs_3_17_port, 
                           A_shifted(16) => positive_inputs_3_16_port, 
                           A_shifted(15) => positive_inputs_3_15_port, 
                           A_shifted(14) => positive_inputs_3_14_port, 
                           A_shifted(13) => positive_inputs_3_13_port, 
                           A_shifted(12) => positive_inputs_3_12_port, 
                           A_shifted(11) => positive_inputs_3_11_port, 
                           A_shifted(10) => positive_inputs_3_10_port, 
                           A_shifted(9) => positive_inputs_3_9_port, 
                           A_shifted(8) => positive_inputs_3_8_port, 
                           A_shifted(7) => positive_inputs_3_7_port, 
                           A_shifted(6) => positive_inputs_3_6_port, 
                           A_shifted(5) => positive_inputs_3_5_port, 
                           A_shifted(4) => positive_inputs_3_4_port, 
                           A_shifted(3) => positive_inputs_3_3_port, 
                           A_shifted(2) => positive_inputs_3_2_port, 
                           A_shifted(1) => positive_inputs_3_1_port, 
                           A_shifted(0) => n9, A_neg_shifted(63) => 
                           negative_inputs_3_63_port, A_neg_shifted(62) => 
                           negative_inputs_3_62_port, A_neg_shifted(61) => 
                           negative_inputs_3_61_port, A_neg_shifted(60) => 
                           negative_inputs_3_60_port, A_neg_shifted(59) => 
                           negative_inputs_3_59_port, A_neg_shifted(58) => 
                           negative_inputs_3_58_port, A_neg_shifted(57) => 
                           negative_inputs_3_57_port, A_neg_shifted(56) => 
                           negative_inputs_3_56_port, A_neg_shifted(55) => 
                           negative_inputs_3_55_port, A_neg_shifted(54) => 
                           negative_inputs_3_54_port, A_neg_shifted(53) => 
                           negative_inputs_3_53_port, A_neg_shifted(52) => 
                           negative_inputs_3_52_port, A_neg_shifted(51) => 
                           negative_inputs_3_51_port, A_neg_shifted(50) => 
                           negative_inputs_3_50_port, A_neg_shifted(49) => 
                           negative_inputs_3_49_port, A_neg_shifted(48) => 
                           negative_inputs_3_48_port, A_neg_shifted(47) => 
                           negative_inputs_3_47_port, A_neg_shifted(46) => 
                           negative_inputs_3_46_port, A_neg_shifted(45) => 
                           negative_inputs_3_45_port, A_neg_shifted(44) => 
                           negative_inputs_3_44_port, A_neg_shifted(43) => 
                           negative_inputs_3_43_port, A_neg_shifted(42) => 
                           negative_inputs_3_42_port, A_neg_shifted(41) => 
                           negative_inputs_3_41_port, A_neg_shifted(40) => 
                           negative_inputs_3_40_port, A_neg_shifted(39) => n145
                           , A_neg_shifted(38) => negative_inputs_3_38_port, 
                           A_neg_shifted(37) => negative_inputs_3_37_port, 
                           A_neg_shifted(36) => negative_inputs_3_36_port, 
                           A_neg_shifted(35) => negative_inputs_3_35_port, 
                           A_neg_shifted(34) => negative_inputs_3_34_port, 
                           A_neg_shifted(33) => negative_inputs_3_33_port, 
                           A_neg_shifted(32) => negative_inputs_3_32_port, 
                           A_neg_shifted(31) => negative_inputs_3_31_port, 
                           A_neg_shifted(30) => negative_inputs_3_30_port, 
                           A_neg_shifted(29) => negative_inputs_3_29_port, 
                           A_neg_shifted(28) => negative_inputs_3_28_port, 
                           A_neg_shifted(27) => negative_inputs_3_27_port, 
                           A_neg_shifted(26) => negative_inputs_3_26_port, 
                           A_neg_shifted(25) => negative_inputs_3_25_port, 
                           A_neg_shifted(24) => negative_inputs_3_24_port, 
                           A_neg_shifted(23) => negative_inputs_3_23_port, 
                           A_neg_shifted(22) => negative_inputs_3_22_port, 
                           A_neg_shifted(21) => negative_inputs_3_21_port, 
                           A_neg_shifted(20) => negative_inputs_3_20_port, 
                           A_neg_shifted(19) => negative_inputs_3_19_port, 
                           A_neg_shifted(18) => negative_inputs_3_18_port, 
                           A_neg_shifted(17) => negative_inputs_3_17_port, 
                           A_neg_shifted(16) => negative_inputs_3_16_port, 
                           A_neg_shifted(15) => negative_inputs_3_15_port, 
                           A_neg_shifted(14) => negative_inputs_3_14_port, 
                           A_neg_shifted(13) => negative_inputs_3_13_port, 
                           A_neg_shifted(12) => negative_inputs_3_12_port, 
                           A_neg_shifted(11) => negative_inputs_3_11_port, 
                           A_neg_shifted(10) => negative_inputs_3_10_port, 
                           A_neg_shifted(9) => negative_inputs_3_9_port, 
                           A_neg_shifted(8) => negative_inputs_3_8_port, 
                           A_neg_shifted(7) => negative_inputs_3_7_port, 
                           A_neg_shifted(6) => negative_inputs_3_6_port, 
                           A_neg_shifted(5) => negative_inputs_3_5_port, 
                           A_neg_shifted(4) => negative_inputs_3_4_port, 
                           A_neg_shifted(3) => negative_inputs_3_3_port, 
                           A_neg_shifted(2) => negative_inputs_3_2_port, 
                           A_neg_shifted(1) => negative_inputs_3_1_port, 
                           A_neg_shifted(0) => n9, Sel(2) => sel_1_2_port, 
                           Sel(1) => sel_1_1_port, Sel(0) => sel_1_0_port, 
                           Y(63) => MuxOutputs_1_63_port, Y(62) => 
                           MuxOutputs_1_62_port, Y(61) => MuxOutputs_1_61_port,
                           Y(60) => MuxOutputs_1_60_port, Y(59) => 
                           MuxOutputs_1_59_port, Y(58) => MuxOutputs_1_58_port,
                           Y(57) => MuxOutputs_1_57_port, Y(56) => 
                           MuxOutputs_1_56_port, Y(55) => MuxOutputs_1_55_port,
                           Y(54) => MuxOutputs_1_54_port, Y(53) => 
                           MuxOutputs_1_53_port, Y(52) => MuxOutputs_1_52_port,
                           Y(51) => MuxOutputs_1_51_port, Y(50) => 
                           MuxOutputs_1_50_port, Y(49) => MuxOutputs_1_49_port,
                           Y(48) => MuxOutputs_1_48_port, Y(47) => 
                           MuxOutputs_1_47_port, Y(46) => MuxOutputs_1_46_port,
                           Y(45) => MuxOutputs_1_45_port, Y(44) => 
                           MuxOutputs_1_44_port, Y(43) => MuxOutputs_1_43_port,
                           Y(42) => MuxOutputs_1_42_port, Y(41) => 
                           MuxOutputs_1_41_port, Y(40) => MuxOutputs_1_40_port,
                           Y(39) => MuxOutputs_1_39_port, Y(38) => 
                           MuxOutputs_1_38_port, Y(37) => MuxOutputs_1_37_port,
                           Y(36) => MuxOutputs_1_36_port, Y(35) => 
                           MuxOutputs_1_35_port, Y(34) => MuxOutputs_1_34_port,
                           Y(33) => MuxOutputs_1_33_port, Y(32) => 
                           MuxOutputs_1_32_port, Y(31) => MuxOutputs_1_31_port,
                           Y(30) => MuxOutputs_1_30_port, Y(29) => 
                           MuxOutputs_1_29_port, Y(28) => MuxOutputs_1_28_port,
                           Y(27) => MuxOutputs_1_27_port, Y(26) => 
                           MuxOutputs_1_26_port, Y(25) => MuxOutputs_1_25_port,
                           Y(24) => MuxOutputs_1_24_port, Y(23) => 
                           MuxOutputs_1_23_port, Y(22) => MuxOutputs_1_22_port,
                           Y(21) => MuxOutputs_1_21_port, Y(20) => 
                           MuxOutputs_1_20_port, Y(19) => MuxOutputs_1_19_port,
                           Y(18) => MuxOutputs_1_18_port, Y(17) => 
                           MuxOutputs_1_17_port, Y(16) => MuxOutputs_1_16_port,
                           Y(15) => MuxOutputs_1_15_port, Y(14) => 
                           MuxOutputs_1_14_port, Y(13) => MuxOutputs_1_13_port,
                           Y(12) => MuxOutputs_1_12_port, Y(11) => 
                           MuxOutputs_1_11_port, Y(10) => MuxOutputs_1_10_port,
                           Y(9) => MuxOutputs_1_9_port, Y(8) => 
                           MuxOutputs_1_8_port, Y(7) => MuxOutputs_1_7_port, 
                           Y(6) => MuxOutputs_1_6_port, Y(5) => 
                           MuxOutputs_1_5_port, Y(4) => MuxOutputs_1_4_port, 
                           Y(3) => MuxOutputs_1_3_port, Y(2) => 
                           MuxOutputs_1_2_port, Y(1) => MuxOutputs_1_1_port, 
                           Y(0) => MuxOutputs_1_0_port);
   encoderI_2 : encoder_14 port map( pieceofB(2) => B(5), pieceofB(1) => B(4), 
                           pieceofB(0) => B(3), sel(2) => sel_2_2_port, sel(1) 
                           => sel_2_1_port, sel(0) => sel_2_0_port);
   MUXI_2 : MUX51_MuxNbit64_14 port map( zeroSignal(63) => X_Logic0_port, 
                           zeroSignal(62) => X_Logic0_port, zeroSignal(61) => 
                           X_Logic0_port, zeroSignal(60) => X_Logic0_port, 
                           zeroSignal(59) => X_Logic0_port, zeroSignal(58) => 
                           X_Logic0_port, zeroSignal(57) => X_Logic0_port, 
                           zeroSignal(56) => X_Logic0_port, zeroSignal(55) => 
                           X_Logic0_port, zeroSignal(54) => X_Logic0_port, 
                           zeroSignal(53) => X_Logic0_port, zeroSignal(52) => 
                           X_Logic0_port, zeroSignal(51) => X_Logic0_port, 
                           zeroSignal(50) => X_Logic0_port, zeroSignal(49) => 
                           X_Logic0_port, zeroSignal(48) => X_Logic0_port, 
                           zeroSignal(47) => X_Logic0_port, zeroSignal(46) => 
                           X_Logic0_port, zeroSignal(45) => X_Logic0_port, 
                           zeroSignal(44) => X_Logic0_port, zeroSignal(43) => 
                           X_Logic0_port, zeroSignal(42) => X_Logic0_port, 
                           zeroSignal(41) => X_Logic0_port, zeroSignal(40) => 
                           X_Logic0_port, zeroSignal(39) => X_Logic0_port, 
                           zeroSignal(38) => X_Logic0_port, zeroSignal(37) => 
                           X_Logic0_port, zeroSignal(36) => X_Logic0_port, 
                           zeroSignal(35) => X_Logic0_port, zeroSignal(34) => 
                           X_Logic0_port, zeroSignal(33) => X_Logic0_port, 
                           zeroSignal(32) => X_Logic0_port, zeroSignal(31) => 
                           X_Logic0_port, zeroSignal(30) => X_Logic0_port, 
                           zeroSignal(29) => X_Logic0_port, zeroSignal(28) => 
                           X_Logic0_port, zeroSignal(27) => X_Logic0_port, 
                           zeroSignal(26) => X_Logic0_port, zeroSignal(25) => 
                           X_Logic0_port, zeroSignal(24) => X_Logic0_port, 
                           zeroSignal(23) => X_Logic0_port, zeroSignal(22) => 
                           X_Logic0_port, zeroSignal(21) => X_Logic0_port, 
                           zeroSignal(20) => X_Logic0_port, zeroSignal(19) => 
                           X_Logic0_port, zeroSignal(18) => X_Logic0_port, 
                           zeroSignal(17) => X_Logic0_port, zeroSignal(16) => 
                           X_Logic0_port, zeroSignal(15) => X_Logic0_port, 
                           zeroSignal(14) => X_Logic0_port, zeroSignal(13) => 
                           X_Logic0_port, zeroSignal(12) => X_Logic0_port, 
                           zeroSignal(11) => X_Logic0_port, zeroSignal(10) => 
                           X_Logic0_port, zeroSignal(9) => X_Logic0_port, 
                           zeroSignal(8) => X_Logic0_port, zeroSignal(7) => 
                           X_Logic0_port, zeroSignal(6) => X_Logic0_port, 
                           zeroSignal(5) => X_Logic0_port, zeroSignal(4) => 
                           X_Logic0_port, zeroSignal(3) => X_Logic0_port, 
                           zeroSignal(2) => X_Logic0_port, zeroSignal(1) => 
                           X_Logic0_port, zeroSignal(0) => X_Logic0_port, 
                           A_signal(63) => positive_inputs_4_63_port, 
                           A_signal(62) => positive_inputs_4_62_port, 
                           A_signal(61) => positive_inputs_4_61_port, 
                           A_signal(60) => positive_inputs_4_60_port, 
                           A_signal(59) => positive_inputs_4_59_port, 
                           A_signal(58) => positive_inputs_4_58_port, 
                           A_signal(57) => positive_inputs_4_57_port, 
                           A_signal(56) => positive_inputs_4_56_port, 
                           A_signal(55) => positive_inputs_4_55_port, 
                           A_signal(54) => positive_inputs_4_54_port, 
                           A_signal(53) => positive_inputs_4_53_port, 
                           A_signal(52) => positive_inputs_4_52_port, 
                           A_signal(51) => positive_inputs_4_51_port, 
                           A_signal(50) => positive_inputs_4_50_port, 
                           A_signal(49) => positive_inputs_4_49_port, 
                           A_signal(48) => n68, A_signal(47) => 
                           positive_inputs_4_47_port, A_signal(46) => 
                           positive_inputs_4_46_port, A_signal(45) => 
                           positive_inputs_4_45_port, A_signal(44) => 
                           positive_inputs_4_44_port, A_signal(43) => 
                           positive_inputs_4_43_port, A_signal(42) => 
                           positive_inputs_4_42_port, A_signal(41) => 
                           positive_inputs_4_41_port, A_signal(40) => 
                           positive_inputs_4_40_port, A_signal(39) => n55, 
                           A_signal(38) => positive_inputs_4_38_port, 
                           A_signal(37) => positive_inputs_4_37_port, 
                           A_signal(36) => positive_inputs_4_36_port, 
                           A_signal(35) => positive_inputs_4_35_port, 
                           A_signal(34) => positive_inputs_4_34_port, 
                           A_signal(33) => positive_inputs_4_33_port, 
                           A_signal(32) => positive_inputs_4_32_port, 
                           A_signal(31) => positive_inputs_4_31_port, 
                           A_signal(30) => positive_inputs_4_30_port, 
                           A_signal(29) => positive_inputs_4_29_port, 
                           A_signal(28) => positive_inputs_4_28_port, 
                           A_signal(27) => positive_inputs_4_27_port, 
                           A_signal(26) => positive_inputs_4_26_port, 
                           A_signal(25) => positive_inputs_4_25_port, 
                           A_signal(24) => positive_inputs_4_24_port, 
                           A_signal(23) => positive_inputs_4_23_port, 
                           A_signal(22) => positive_inputs_4_22_port, 
                           A_signal(21) => positive_inputs_4_21_port, 
                           A_signal(20) => positive_inputs_4_20_port, 
                           A_signal(19) => positive_inputs_4_19_port, 
                           A_signal(18) => positive_inputs_4_18_port, 
                           A_signal(17) => positive_inputs_4_17_port, 
                           A_signal(16) => positive_inputs_4_16_port, 
                           A_signal(15) => positive_inputs_4_15_port, 
                           A_signal(14) => positive_inputs_4_14_port, 
                           A_signal(13) => positive_inputs_4_13_port, 
                           A_signal(12) => positive_inputs_4_12_port, 
                           A_signal(11) => positive_inputs_4_11_port, 
                           A_signal(10) => positive_inputs_4_10_port, 
                           A_signal(9) => positive_inputs_4_9_port, A_signal(8)
                           => positive_inputs_4_8_port, A_signal(7) => 
                           positive_inputs_4_7_port, A_signal(6) => 
                           positive_inputs_4_6_port, A_signal(5) => 
                           positive_inputs_4_5_port, A_signal(4) => 
                           positive_inputs_4_4_port, A_signal(3) => 
                           positive_inputs_4_3_port, A_signal(2) => 
                           positive_inputs_4_2_port, A_signal(1) => 
                           positive_inputs_4_1_port, A_signal(0) => n9, 
                           A_neg(63) => negative_inputs_4_63_port, A_neg(62) =>
                           negative_inputs_4_62_port, A_neg(61) => 
                           negative_inputs_4_61_port, A_neg(60) => 
                           negative_inputs_4_60_port, A_neg(59) => 
                           negative_inputs_4_59_port, A_neg(58) => 
                           negative_inputs_4_58_port, A_neg(57) => 
                           negative_inputs_4_57_port, A_neg(56) => 
                           negative_inputs_4_56_port, A_neg(55) => 
                           negative_inputs_4_55_port, A_neg(54) => 
                           negative_inputs_4_54_port, A_neg(53) => 
                           negative_inputs_4_53_port, A_neg(52) => 
                           negative_inputs_4_52_port, A_neg(51) => 
                           negative_inputs_4_51_port, A_neg(50) => 
                           negative_inputs_4_50_port, A_neg(49) => 
                           negative_inputs_4_49_port, A_neg(48) => 
                           negative_inputs_4_48_port, A_neg(47) => 
                           negative_inputs_4_47_port, A_neg(46) => 
                           negative_inputs_4_46_port, A_neg(45) => 
                           negative_inputs_4_45_port, A_neg(44) => 
                           negative_inputs_4_44_port, A_neg(43) => 
                           negative_inputs_4_43_port, A_neg(42) => 
                           negative_inputs_4_42_port, A_neg(41) => 
                           negative_inputs_4_41_port, A_neg(40) => 
                           negative_inputs_4_40_port, A_neg(39) => n143, 
                           A_neg(38) => negative_inputs_4_38_port, A_neg(37) =>
                           negative_inputs_4_37_port, A_neg(36) => 
                           negative_inputs_4_36_port, A_neg(35) => 
                           negative_inputs_4_35_port, A_neg(34) => 
                           negative_inputs_4_34_port, A_neg(33) => 
                           negative_inputs_4_33_port, A_neg(32) => 
                           negative_inputs_4_32_port, A_neg(31) => 
                           negative_inputs_4_31_port, A_neg(30) => 
                           negative_inputs_4_30_port, A_neg(29) => 
                           negative_inputs_4_29_port, A_neg(28) => 
                           negative_inputs_4_28_port, A_neg(27) => 
                           negative_inputs_4_27_port, A_neg(26) => 
                           negative_inputs_4_26_port, A_neg(25) => 
                           negative_inputs_4_25_port, A_neg(24) => 
                           negative_inputs_4_24_port, A_neg(23) => 
                           negative_inputs_4_23_port, A_neg(22) => 
                           negative_inputs_4_22_port, A_neg(21) => 
                           negative_inputs_4_21_port, A_neg(20) => 
                           negative_inputs_4_20_port, A_neg(19) => 
                           negative_inputs_4_19_port, A_neg(18) => 
                           negative_inputs_4_18_port, A_neg(17) => 
                           negative_inputs_4_17_port, A_neg(16) => 
                           negative_inputs_4_16_port, A_neg(15) => 
                           negative_inputs_4_15_port, A_neg(14) => 
                           negative_inputs_4_14_port, A_neg(13) => 
                           negative_inputs_4_13_port, A_neg(12) => 
                           negative_inputs_4_12_port, A_neg(11) => 
                           negative_inputs_4_11_port, A_neg(10) => 
                           negative_inputs_4_10_port, A_neg(9) => 
                           negative_inputs_4_9_port, A_neg(8) => 
                           negative_inputs_4_8_port, A_neg(7) => 
                           negative_inputs_4_7_port, A_neg(6) => 
                           negative_inputs_4_6_port, A_neg(5) => 
                           negative_inputs_4_5_port, A_neg(4) => 
                           negative_inputs_4_4_port, A_neg(3) => 
                           negative_inputs_4_3_port, A_neg(2) => 
                           negative_inputs_4_2_port, A_neg(1) => 
                           negative_inputs_4_1_port, A_neg(0) => n9, 
                           A_shifted(63) => positive_inputs_5_63_port, 
                           A_shifted(62) => positive_inputs_5_62_port, 
                           A_shifted(61) => positive_inputs_5_61_port, 
                           A_shifted(60) => positive_inputs_5_60_port, 
                           A_shifted(59) => positive_inputs_5_59_port, 
                           A_shifted(58) => positive_inputs_5_58_port, 
                           A_shifted(57) => positive_inputs_5_57_port, 
                           A_shifted(56) => positive_inputs_5_56_port, 
                           A_shifted(55) => positive_inputs_5_55_port, 
                           A_shifted(54) => positive_inputs_5_54_port, 
                           A_shifted(53) => positive_inputs_5_53_port, 
                           A_shifted(52) => positive_inputs_5_52_port, 
                           A_shifted(51) => positive_inputs_5_51_port, 
                           A_shifted(50) => positive_inputs_5_50_port, 
                           A_shifted(49) => positive_inputs_5_49_port, 
                           A_shifted(48) => n67, A_shifted(47) => 
                           positive_inputs_5_47_port, A_shifted(46) => 
                           positive_inputs_5_46_port, A_shifted(45) => 
                           positive_inputs_5_45_port, A_shifted(44) => 
                           positive_inputs_5_44_port, A_shifted(43) => 
                           positive_inputs_5_43_port, A_shifted(42) => 
                           positive_inputs_5_42_port, A_shifted(41) => 
                           positive_inputs_5_41_port, A_shifted(40) => 
                           positive_inputs_5_40_port, A_shifted(39) => n54, 
                           A_shifted(38) => positive_inputs_5_38_port, 
                           A_shifted(37) => positive_inputs_5_37_port, 
                           A_shifted(36) => positive_inputs_5_36_port, 
                           A_shifted(35) => positive_inputs_5_35_port, 
                           A_shifted(34) => positive_inputs_5_34_port, 
                           A_shifted(33) => positive_inputs_5_33_port, 
                           A_shifted(32) => positive_inputs_5_32_port, 
                           A_shifted(31) => positive_inputs_5_31_port, 
                           A_shifted(30) => positive_inputs_5_30_port, 
                           A_shifted(29) => positive_inputs_5_29_port, 
                           A_shifted(28) => positive_inputs_5_28_port, 
                           A_shifted(27) => positive_inputs_5_27_port, 
                           A_shifted(26) => positive_inputs_5_26_port, 
                           A_shifted(25) => positive_inputs_5_25_port, 
                           A_shifted(24) => positive_inputs_5_24_port, 
                           A_shifted(23) => positive_inputs_5_23_port, 
                           A_shifted(22) => positive_inputs_5_22_port, 
                           A_shifted(21) => positive_inputs_5_21_port, 
                           A_shifted(20) => positive_inputs_5_20_port, 
                           A_shifted(19) => positive_inputs_5_19_port, 
                           A_shifted(18) => positive_inputs_5_18_port, 
                           A_shifted(17) => positive_inputs_5_17_port, 
                           A_shifted(16) => positive_inputs_5_16_port, 
                           A_shifted(15) => positive_inputs_5_15_port, 
                           A_shifted(14) => positive_inputs_5_14_port, 
                           A_shifted(13) => positive_inputs_5_13_port, 
                           A_shifted(12) => positive_inputs_5_12_port, 
                           A_shifted(11) => positive_inputs_5_11_port, 
                           A_shifted(10) => positive_inputs_5_10_port, 
                           A_shifted(9) => positive_inputs_5_9_port, 
                           A_shifted(8) => positive_inputs_5_8_port, 
                           A_shifted(7) => positive_inputs_5_7_port, 
                           A_shifted(6) => positive_inputs_5_6_port, 
                           A_shifted(5) => positive_inputs_5_5_port, 
                           A_shifted(4) => positive_inputs_5_4_port, 
                           A_shifted(3) => positive_inputs_5_3_port, 
                           A_shifted(2) => positive_inputs_5_2_port, 
                           A_shifted(1) => positive_inputs_5_1_port, 
                           A_shifted(0) => n9, A_neg_shifted(63) => 
                           negative_inputs_5_63_port, A_neg_shifted(62) => 
                           negative_inputs_5_62_port, A_neg_shifted(61) => 
                           negative_inputs_5_61_port, A_neg_shifted(60) => 
                           negative_inputs_5_60_port, A_neg_shifted(59) => 
                           negative_inputs_5_59_port, A_neg_shifted(58) => 
                           negative_inputs_5_58_port, A_neg_shifted(57) => 
                           negative_inputs_5_57_port, A_neg_shifted(56) => 
                           negative_inputs_5_56_port, A_neg_shifted(55) => 
                           negative_inputs_5_55_port, A_neg_shifted(54) => 
                           negative_inputs_5_54_port, A_neg_shifted(53) => 
                           negative_inputs_5_53_port, A_neg_shifted(52) => 
                           negative_inputs_5_52_port, A_neg_shifted(51) => 
                           negative_inputs_5_51_port, A_neg_shifted(50) => 
                           negative_inputs_5_50_port, A_neg_shifted(49) => 
                           negative_inputs_5_49_port, A_neg_shifted(48) => 
                           negative_inputs_5_48_port, A_neg_shifted(47) => 
                           negative_inputs_5_47_port, A_neg_shifted(46) => 
                           negative_inputs_5_46_port, A_neg_shifted(45) => 
                           negative_inputs_5_45_port, A_neg_shifted(44) => 
                           negative_inputs_5_44_port, A_neg_shifted(43) => 
                           negative_inputs_5_43_port, A_neg_shifted(42) => 
                           negative_inputs_5_42_port, A_neg_shifted(41) => 
                           negative_inputs_5_41_port, A_neg_shifted(40) => 
                           negative_inputs_5_40_port, A_neg_shifted(39) => n141
                           , A_neg_shifted(38) => negative_inputs_5_38_port, 
                           A_neg_shifted(37) => negative_inputs_5_37_port, 
                           A_neg_shifted(36) => negative_inputs_5_36_port, 
                           A_neg_shifted(35) => negative_inputs_5_35_port, 
                           A_neg_shifted(34) => negative_inputs_5_34_port, 
                           A_neg_shifted(33) => negative_inputs_5_33_port, 
                           A_neg_shifted(32) => negative_inputs_5_32_port, 
                           A_neg_shifted(31) => negative_inputs_5_31_port, 
                           A_neg_shifted(30) => negative_inputs_5_30_port, 
                           A_neg_shifted(29) => negative_inputs_5_29_port, 
                           A_neg_shifted(28) => negative_inputs_5_28_port, 
                           A_neg_shifted(27) => negative_inputs_5_27_port, 
                           A_neg_shifted(26) => negative_inputs_5_26_port, 
                           A_neg_shifted(25) => negative_inputs_5_25_port, 
                           A_neg_shifted(24) => negative_inputs_5_24_port, 
                           A_neg_shifted(23) => negative_inputs_5_23_port, 
                           A_neg_shifted(22) => negative_inputs_5_22_port, 
                           A_neg_shifted(21) => negative_inputs_5_21_port, 
                           A_neg_shifted(20) => negative_inputs_5_20_port, 
                           A_neg_shifted(19) => negative_inputs_5_19_port, 
                           A_neg_shifted(18) => negative_inputs_5_18_port, 
                           A_neg_shifted(17) => negative_inputs_5_17_port, 
                           A_neg_shifted(16) => negative_inputs_5_16_port, 
                           A_neg_shifted(15) => negative_inputs_5_15_port, 
                           A_neg_shifted(14) => negative_inputs_5_14_port, 
                           A_neg_shifted(13) => negative_inputs_5_13_port, 
                           A_neg_shifted(12) => negative_inputs_5_12_port, 
                           A_neg_shifted(11) => negative_inputs_5_11_port, 
                           A_neg_shifted(10) => negative_inputs_5_10_port, 
                           A_neg_shifted(9) => negative_inputs_5_9_port, 
                           A_neg_shifted(8) => negative_inputs_5_8_port, 
                           A_neg_shifted(7) => negative_inputs_5_7_port, 
                           A_neg_shifted(6) => negative_inputs_5_6_port, 
                           A_neg_shifted(5) => negative_inputs_5_5_port, 
                           A_neg_shifted(4) => negative_inputs_5_4_port, 
                           A_neg_shifted(3) => negative_inputs_5_3_port, 
                           A_neg_shifted(2) => negative_inputs_5_2_port, 
                           A_neg_shifted(1) => negative_inputs_5_1_port, 
                           A_neg_shifted(0) => n9, Sel(2) => sel_2_2_port, 
                           Sel(1) => sel_2_1_port, Sel(0) => sel_2_0_port, 
                           Y(63) => MuxOutputs_2_63_port, Y(62) => 
                           MuxOutputs_2_62_port, Y(61) => MuxOutputs_2_61_port,
                           Y(60) => MuxOutputs_2_60_port, Y(59) => 
                           MuxOutputs_2_59_port, Y(58) => MuxOutputs_2_58_port,
                           Y(57) => MuxOutputs_2_57_port, Y(56) => 
                           MuxOutputs_2_56_port, Y(55) => MuxOutputs_2_55_port,
                           Y(54) => MuxOutputs_2_54_port, Y(53) => 
                           MuxOutputs_2_53_port, Y(52) => MuxOutputs_2_52_port,
                           Y(51) => MuxOutputs_2_51_port, Y(50) => 
                           MuxOutputs_2_50_port, Y(49) => MuxOutputs_2_49_port,
                           Y(48) => MuxOutputs_2_48_port, Y(47) => 
                           MuxOutputs_2_47_port, Y(46) => MuxOutputs_2_46_port,
                           Y(45) => MuxOutputs_2_45_port, Y(44) => 
                           MuxOutputs_2_44_port, Y(43) => MuxOutputs_2_43_port,
                           Y(42) => MuxOutputs_2_42_port, Y(41) => 
                           MuxOutputs_2_41_port, Y(40) => MuxOutputs_2_40_port,
                           Y(39) => MuxOutputs_2_39_port, Y(38) => 
                           MuxOutputs_2_38_port, Y(37) => MuxOutputs_2_37_port,
                           Y(36) => MuxOutputs_2_36_port, Y(35) => 
                           MuxOutputs_2_35_port, Y(34) => MuxOutputs_2_34_port,
                           Y(33) => MuxOutputs_2_33_port, Y(32) => 
                           MuxOutputs_2_32_port, Y(31) => MuxOutputs_2_31_port,
                           Y(30) => MuxOutputs_2_30_port, Y(29) => 
                           MuxOutputs_2_29_port, Y(28) => MuxOutputs_2_28_port,
                           Y(27) => MuxOutputs_2_27_port, Y(26) => 
                           MuxOutputs_2_26_port, Y(25) => MuxOutputs_2_25_port,
                           Y(24) => MuxOutputs_2_24_port, Y(23) => 
                           MuxOutputs_2_23_port, Y(22) => MuxOutputs_2_22_port,
                           Y(21) => MuxOutputs_2_21_port, Y(20) => 
                           MuxOutputs_2_20_port, Y(19) => MuxOutputs_2_19_port,
                           Y(18) => MuxOutputs_2_18_port, Y(17) => 
                           MuxOutputs_2_17_port, Y(16) => MuxOutputs_2_16_port,
                           Y(15) => MuxOutputs_2_15_port, Y(14) => 
                           MuxOutputs_2_14_port, Y(13) => MuxOutputs_2_13_port,
                           Y(12) => MuxOutputs_2_12_port, Y(11) => 
                           MuxOutputs_2_11_port, Y(10) => MuxOutputs_2_10_port,
                           Y(9) => MuxOutputs_2_9_port, Y(8) => 
                           MuxOutputs_2_8_port, Y(7) => MuxOutputs_2_7_port, 
                           Y(6) => MuxOutputs_2_6_port, Y(5) => 
                           MuxOutputs_2_5_port, Y(4) => MuxOutputs_2_4_port, 
                           Y(3) => MuxOutputs_2_3_port, Y(2) => 
                           MuxOutputs_2_2_port, Y(1) => MuxOutputs_2_1_port, 
                           Y(0) => MuxOutputs_2_0_port);
   encoderI_3 : encoder_13 port map( pieceofB(2) => B(7), pieceofB(1) => B(6), 
                           pieceofB(0) => B(5), sel(2) => sel_3_2_port, sel(1) 
                           => sel_3_1_port, sel(0) => sel_3_0_port);
   MUXI_3 : MUX51_MuxNbit64_13 port map( zeroSignal(63) => X_Logic0_port, 
                           zeroSignal(62) => X_Logic0_port, zeroSignal(61) => 
                           X_Logic0_port, zeroSignal(60) => X_Logic0_port, 
                           zeroSignal(59) => X_Logic0_port, zeroSignal(58) => 
                           X_Logic0_port, zeroSignal(57) => X_Logic0_port, 
                           zeroSignal(56) => X_Logic0_port, zeroSignal(55) => 
                           X_Logic0_port, zeroSignal(54) => X_Logic0_port, 
                           zeroSignal(53) => X_Logic0_port, zeroSignal(52) => 
                           X_Logic0_port, zeroSignal(51) => X_Logic0_port, 
                           zeroSignal(50) => X_Logic0_port, zeroSignal(49) => 
                           X_Logic0_port, zeroSignal(48) => X_Logic0_port, 
                           zeroSignal(47) => X_Logic0_port, zeroSignal(46) => 
                           X_Logic0_port, zeroSignal(45) => X_Logic0_port, 
                           zeroSignal(44) => X_Logic0_port, zeroSignal(43) => 
                           X_Logic0_port, zeroSignal(42) => X_Logic0_port, 
                           zeroSignal(41) => X_Logic0_port, zeroSignal(40) => 
                           X_Logic0_port, zeroSignal(39) => X_Logic0_port, 
                           zeroSignal(38) => X_Logic0_port, zeroSignal(37) => 
                           X_Logic0_port, zeroSignal(36) => X_Logic0_port, 
                           zeroSignal(35) => X_Logic0_port, zeroSignal(34) => 
                           X_Logic0_port, zeroSignal(33) => X_Logic0_port, 
                           zeroSignal(32) => X_Logic0_port, zeroSignal(31) => 
                           X_Logic0_port, zeroSignal(30) => X_Logic0_port, 
                           zeroSignal(29) => X_Logic0_port, zeroSignal(28) => 
                           X_Logic0_port, zeroSignal(27) => X_Logic0_port, 
                           zeroSignal(26) => X_Logic0_port, zeroSignal(25) => 
                           X_Logic0_port, zeroSignal(24) => X_Logic0_port, 
                           zeroSignal(23) => X_Logic0_port, zeroSignal(22) => 
                           X_Logic0_port, zeroSignal(21) => X_Logic0_port, 
                           zeroSignal(20) => X_Logic0_port, zeroSignal(19) => 
                           X_Logic0_port, zeroSignal(18) => X_Logic0_port, 
                           zeroSignal(17) => X_Logic0_port, zeroSignal(16) => 
                           X_Logic0_port, zeroSignal(15) => X_Logic0_port, 
                           zeroSignal(14) => X_Logic0_port, zeroSignal(13) => 
                           X_Logic0_port, zeroSignal(12) => X_Logic0_port, 
                           zeroSignal(11) => X_Logic0_port, zeroSignal(10) => 
                           X_Logic0_port, zeroSignal(9) => X_Logic0_port, 
                           zeroSignal(8) => X_Logic0_port, zeroSignal(7) => 
                           X_Logic0_port, zeroSignal(6) => X_Logic0_port, 
                           zeroSignal(5) => X_Logic0_port, zeroSignal(4) => 
                           X_Logic0_port, zeroSignal(3) => X_Logic0_port, 
                           zeroSignal(2) => X_Logic0_port, zeroSignal(1) => 
                           X_Logic0_port, zeroSignal(0) => X_Logic0_port, 
                           A_signal(63) => positive_inputs_6_63_port, 
                           A_signal(62) => positive_inputs_6_62_port, 
                           A_signal(61) => positive_inputs_6_61_port, 
                           A_signal(60) => positive_inputs_6_60_port, 
                           A_signal(59) => positive_inputs_6_59_port, 
                           A_signal(58) => positive_inputs_6_58_port, 
                           A_signal(57) => positive_inputs_6_57_port, 
                           A_signal(56) => positive_inputs_6_56_port, 
                           A_signal(55) => positive_inputs_6_55_port, 
                           A_signal(54) => positive_inputs_6_54_port, 
                           A_signal(53) => positive_inputs_6_53_port, 
                           A_signal(52) => positive_inputs_6_52_port, 
                           A_signal(51) => positive_inputs_6_51_port, 
                           A_signal(50) => positive_inputs_6_50_port, 
                           A_signal(49) => positive_inputs_6_49_port, 
                           A_signal(48) => positive_inputs_6_48_port, 
                           A_signal(47) => positive_inputs_6_47_port, 
                           A_signal(46) => positive_inputs_6_46_port, 
                           A_signal(45) => positive_inputs_6_45_port, 
                           A_signal(44) => positive_inputs_6_44_port, 
                           A_signal(43) => positive_inputs_6_43_port, 
                           A_signal(42) => positive_inputs_6_42_port, 
                           A_signal(41) => positive_inputs_6_41_port, 
                           A_signal(40) => positive_inputs_6_40_port, 
                           A_signal(39) => n53, A_signal(38) => 
                           positive_inputs_6_38_port, A_signal(37) => 
                           positive_inputs_6_37_port, A_signal(36) => 
                           positive_inputs_6_36_port, A_signal(35) => 
                           positive_inputs_6_35_port, A_signal(34) => 
                           positive_inputs_6_34_port, A_signal(33) => 
                           positive_inputs_6_33_port, A_signal(32) => 
                           positive_inputs_6_32_port, A_signal(31) => 
                           positive_inputs_6_31_port, A_signal(30) => 
                           positive_inputs_6_30_port, A_signal(29) => 
                           positive_inputs_6_29_port, A_signal(28) => 
                           positive_inputs_6_28_port, A_signal(27) => 
                           positive_inputs_6_27_port, A_signal(26) => 
                           positive_inputs_6_26_port, A_signal(25) => 
                           positive_inputs_6_25_port, A_signal(24) => 
                           positive_inputs_6_24_port, A_signal(23) => 
                           positive_inputs_6_23_port, A_signal(22) => 
                           positive_inputs_6_22_port, A_signal(21) => 
                           positive_inputs_6_21_port, A_signal(20) => 
                           positive_inputs_6_20_port, A_signal(19) => 
                           positive_inputs_6_19_port, A_signal(18) => 
                           positive_inputs_6_18_port, A_signal(17) => 
                           positive_inputs_6_17_port, A_signal(16) => 
                           positive_inputs_6_16_port, A_signal(15) => 
                           positive_inputs_6_15_port, A_signal(14) => 
                           positive_inputs_6_14_port, A_signal(13) => 
                           positive_inputs_6_13_port, A_signal(12) => 
                           positive_inputs_6_12_port, A_signal(11) => 
                           positive_inputs_6_11_port, A_signal(10) => 
                           positive_inputs_6_10_port, A_signal(9) => 
                           positive_inputs_6_9_port, A_signal(8) => 
                           positive_inputs_6_8_port, A_signal(7) => 
                           positive_inputs_6_7_port, A_signal(6) => 
                           positive_inputs_6_6_port, A_signal(5) => 
                           positive_inputs_6_5_port, A_signal(4) => 
                           positive_inputs_6_4_port, A_signal(3) => 
                           positive_inputs_6_3_port, A_signal(2) => 
                           positive_inputs_6_2_port, A_signal(1) => 
                           positive_inputs_6_1_port, A_signal(0) => n9, 
                           A_neg(63) => negative_inputs_6_63_port, A_neg(62) =>
                           negative_inputs_6_62_port, A_neg(61) => 
                           negative_inputs_6_61_port, A_neg(60) => 
                           negative_inputs_6_60_port, A_neg(59) => 
                           negative_inputs_6_59_port, A_neg(58) => 
                           negative_inputs_6_58_port, A_neg(57) => 
                           negative_inputs_6_57_port, A_neg(56) => 
                           negative_inputs_6_56_port, A_neg(55) => 
                           negative_inputs_6_55_port, A_neg(54) => 
                           negative_inputs_6_54_port, A_neg(53) => 
                           negative_inputs_6_53_port, A_neg(52) => 
                           negative_inputs_6_52_port, A_neg(51) => 
                           negative_inputs_6_51_port, A_neg(50) => 
                           negative_inputs_6_50_port, A_neg(49) => 
                           negative_inputs_6_49_port, A_neg(48) => 
                           negative_inputs_6_48_port, A_neg(47) => 
                           negative_inputs_6_47_port, A_neg(46) => 
                           negative_inputs_6_46_port, A_neg(45) => 
                           negative_inputs_6_45_port, A_neg(44) => 
                           negative_inputs_6_44_port, A_neg(43) => 
                           negative_inputs_6_43_port, A_neg(42) => 
                           negative_inputs_6_42_port, A_neg(41) => 
                           negative_inputs_6_41_port, A_neg(40) => 
                           negative_inputs_6_40_port, A_neg(39) => n139, 
                           A_neg(38) => negative_inputs_6_38_port, A_neg(37) =>
                           negative_inputs_6_37_port, A_neg(36) => 
                           negative_inputs_6_36_port, A_neg(35) => 
                           negative_inputs_6_35_port, A_neg(34) => 
                           negative_inputs_6_34_port, A_neg(33) => 
                           negative_inputs_6_33_port, A_neg(32) => 
                           negative_inputs_6_32_port, A_neg(31) => 
                           negative_inputs_6_31_port, A_neg(30) => 
                           negative_inputs_6_30_port, A_neg(29) => 
                           negative_inputs_6_29_port, A_neg(28) => 
                           negative_inputs_6_28_port, A_neg(27) => 
                           negative_inputs_6_27_port, A_neg(26) => 
                           negative_inputs_6_26_port, A_neg(25) => 
                           negative_inputs_6_25_port, A_neg(24) => 
                           negative_inputs_6_24_port, A_neg(23) => 
                           negative_inputs_6_23_port, A_neg(22) => 
                           negative_inputs_6_22_port, A_neg(21) => 
                           negative_inputs_6_21_port, A_neg(20) => 
                           negative_inputs_6_20_port, A_neg(19) => 
                           negative_inputs_6_19_port, A_neg(18) => 
                           negative_inputs_6_18_port, A_neg(17) => 
                           negative_inputs_6_17_port, A_neg(16) => 
                           negative_inputs_6_16_port, A_neg(15) => 
                           negative_inputs_6_15_port, A_neg(14) => 
                           negative_inputs_6_14_port, A_neg(13) => 
                           negative_inputs_6_13_port, A_neg(12) => 
                           negative_inputs_6_12_port, A_neg(11) => 
                           negative_inputs_6_11_port, A_neg(10) => 
                           negative_inputs_6_10_port, A_neg(9) => 
                           negative_inputs_6_9_port, A_neg(8) => 
                           negative_inputs_6_8_port, A_neg(7) => 
                           negative_inputs_6_7_port, A_neg(6) => 
                           negative_inputs_6_6_port, A_neg(5) => 
                           negative_inputs_6_5_port, A_neg(4) => 
                           negative_inputs_6_4_port, A_neg(3) => 
                           negative_inputs_6_3_port, A_neg(2) => 
                           negative_inputs_6_2_port, A_neg(1) => 
                           negative_inputs_6_1_port, A_neg(0) => n9, 
                           A_shifted(63) => positive_inputs_7_63_port, 
                           A_shifted(62) => positive_inputs_7_62_port, 
                           A_shifted(61) => positive_inputs_7_61_port, 
                           A_shifted(60) => positive_inputs_7_60_port, 
                           A_shifted(59) => positive_inputs_7_59_port, 
                           A_shifted(58) => positive_inputs_7_58_port, 
                           A_shifted(57) => positive_inputs_7_57_port, 
                           A_shifted(56) => positive_inputs_7_56_port, 
                           A_shifted(55) => positive_inputs_7_55_port, 
                           A_shifted(54) => positive_inputs_7_54_port, 
                           A_shifted(53) => positive_inputs_7_53_port, 
                           A_shifted(52) => positive_inputs_7_52_port, 
                           A_shifted(51) => positive_inputs_7_51_port, 
                           A_shifted(50) => positive_inputs_7_50_port, 
                           A_shifted(49) => positive_inputs_7_49_port, 
                           A_shifted(48) => n66, A_shifted(47) => 
                           positive_inputs_7_47_port, A_shifted(46) => 
                           positive_inputs_7_46_port, A_shifted(45) => 
                           positive_inputs_7_45_port, A_shifted(44) => 
                           positive_inputs_7_44_port, A_shifted(43) => 
                           positive_inputs_7_43_port, A_shifted(42) => 
                           positive_inputs_7_42_port, A_shifted(41) => 
                           positive_inputs_7_41_port, A_shifted(40) => 
                           positive_inputs_7_40_port, A_shifted(39) => n52, 
                           A_shifted(38) => n51, A_shifted(37) => n214, 
                           A_shifted(36) => n212, A_shifted(35) => n210, 
                           A_shifted(34) => n208, A_shifted(33) => n206, 
                           A_shifted(32) => n204, A_shifted(31) => n202, 
                           A_shifted(30) => n200, A_shifted(29) => n198, 
                           A_shifted(28) => n196, A_shifted(27) => n194, 
                           A_shifted(26) => n192, A_shifted(25) => n190, 
                           A_shifted(24) => n188, A_shifted(23) => n186, 
                           A_shifted(22) => n184, A_shifted(21) => n182, 
                           A_shifted(20) => n180, A_shifted(19) => n178, 
                           A_shifted(18) => n176, A_shifted(17) => n174, 
                           A_shifted(16) => n172, A_shifted(15) => n170, 
                           A_shifted(14) => n168, A_shifted(13) => n166, 
                           A_shifted(12) => n164, A_shifted(11) => n162, 
                           A_shifted(10) => n160, A_shifted(9) => n158, 
                           A_shifted(8) => n156, A_shifted(7) => n154, 
                           A_shifted(6) => positive_inputs_7_6_port, 
                           A_shifted(5) => positive_inputs_7_5_port, 
                           A_shifted(4) => positive_inputs_7_4_port, 
                           A_shifted(3) => positive_inputs_7_3_port, 
                           A_shifted(2) => positive_inputs_7_2_port, 
                           A_shifted(1) => positive_inputs_7_1_port, 
                           A_shifted(0) => n9, A_neg_shifted(63) => 
                           negative_inputs_7_63_port, A_neg_shifted(62) => 
                           negative_inputs_7_62_port, A_neg_shifted(61) => 
                           negative_inputs_7_61_port, A_neg_shifted(60) => 
                           negative_inputs_7_60_port, A_neg_shifted(59) => 
                           negative_inputs_7_59_port, A_neg_shifted(58) => 
                           negative_inputs_7_58_port, A_neg_shifted(57) => 
                           negative_inputs_7_57_port, A_neg_shifted(56) => 
                           negative_inputs_7_56_port, A_neg_shifted(55) => 
                           negative_inputs_7_55_port, A_neg_shifted(54) => 
                           negative_inputs_7_54_port, A_neg_shifted(53) => 
                           negative_inputs_7_53_port, A_neg_shifted(52) => 
                           negative_inputs_7_52_port, A_neg_shifted(51) => 
                           negative_inputs_7_51_port, A_neg_shifted(50) => 
                           negative_inputs_7_50_port, A_neg_shifted(49) => 
                           negative_inputs_7_49_port, A_neg_shifted(48) => 
                           negative_inputs_7_48_port, A_neg_shifted(47) => 
                           negative_inputs_7_47_port, A_neg_shifted(46) => 
                           negative_inputs_7_46_port, A_neg_shifted(45) => 
                           negative_inputs_7_45_port, A_neg_shifted(44) => 
                           negative_inputs_7_44_port, A_neg_shifted(43) => 
                           negative_inputs_7_43_port, A_neg_shifted(42) => 
                           negative_inputs_7_42_port, A_neg_shifted(41) => 
                           negative_inputs_7_41_port, A_neg_shifted(40) => 
                           negative_inputs_7_40_port, A_neg_shifted(39) => n137
                           , A_neg_shifted(38) => n135, A_neg_shifted(37) => 
                           n133, A_neg_shifted(36) => n131, A_neg_shifted(35) 
                           => n129, A_neg_shifted(34) => n127, 
                           A_neg_shifted(33) => n125, A_neg_shifted(32) => n123
                           , A_neg_shifted(31) => n121, A_neg_shifted(30) => 
                           n119, A_neg_shifted(29) => n117, A_neg_shifted(28) 
                           => n115, A_neg_shifted(27) => n113, 
                           A_neg_shifted(26) => n111, A_neg_shifted(25) => n109
                           , A_neg_shifted(24) => n107, A_neg_shifted(23) => 
                           n105, A_neg_shifted(22) => n103, A_neg_shifted(21) 
                           => n101, A_neg_shifted(20) => n99, A_neg_shifted(19)
                           => n97, A_neg_shifted(18) => n95, A_neg_shifted(17) 
                           => n93, A_neg_shifted(16) => n91, A_neg_shifted(15) 
                           => n89, A_neg_shifted(14) => n87, A_neg_shifted(13) 
                           => n85, A_neg_shifted(12) => n83, A_neg_shifted(11) 
                           => n81, A_neg_shifted(10) => n79, A_neg_shifted(9) 
                           => n77, A_neg_shifted(8) => n75, A_neg_shifted(7) =>
                           n73, A_neg_shifted(6) => negative_inputs_7_6_port, 
                           A_neg_shifted(5) => negative_inputs_7_5_port, 
                           A_neg_shifted(4) => negative_inputs_7_4_port, 
                           A_neg_shifted(3) => negative_inputs_7_3_port, 
                           A_neg_shifted(2) => negative_inputs_7_2_port, 
                           A_neg_shifted(1) => negative_inputs_7_1_port, 
                           A_neg_shifted(0) => n9, Sel(2) => sel_3_2_port, 
                           Sel(1) => sel_3_1_port, Sel(0) => sel_3_0_port, 
                           Y(63) => MuxOutputs_3_63_port, Y(62) => 
                           MuxOutputs_3_62_port, Y(61) => MuxOutputs_3_61_port,
                           Y(60) => MuxOutputs_3_60_port, Y(59) => 
                           MuxOutputs_3_59_port, Y(58) => MuxOutputs_3_58_port,
                           Y(57) => MuxOutputs_3_57_port, Y(56) => 
                           MuxOutputs_3_56_port, Y(55) => MuxOutputs_3_55_port,
                           Y(54) => MuxOutputs_3_54_port, Y(53) => 
                           MuxOutputs_3_53_port, Y(52) => MuxOutputs_3_52_port,
                           Y(51) => MuxOutputs_3_51_port, Y(50) => 
                           MuxOutputs_3_50_port, Y(49) => MuxOutputs_3_49_port,
                           Y(48) => MuxOutputs_3_48_port, Y(47) => 
                           MuxOutputs_3_47_port, Y(46) => MuxOutputs_3_46_port,
                           Y(45) => MuxOutputs_3_45_port, Y(44) => 
                           MuxOutputs_3_44_port, Y(43) => MuxOutputs_3_43_port,
                           Y(42) => MuxOutputs_3_42_port, Y(41) => 
                           MuxOutputs_3_41_port, Y(40) => MuxOutputs_3_40_port,
                           Y(39) => MuxOutputs_3_39_port, Y(38) => 
                           MuxOutputs_3_38_port, Y(37) => MuxOutputs_3_37_port,
                           Y(36) => MuxOutputs_3_36_port, Y(35) => 
                           MuxOutputs_3_35_port, Y(34) => MuxOutputs_3_34_port,
                           Y(33) => MuxOutputs_3_33_port, Y(32) => 
                           MuxOutputs_3_32_port, Y(31) => MuxOutputs_3_31_port,
                           Y(30) => MuxOutputs_3_30_port, Y(29) => 
                           MuxOutputs_3_29_port, Y(28) => MuxOutputs_3_28_port,
                           Y(27) => MuxOutputs_3_27_port, Y(26) => 
                           MuxOutputs_3_26_port, Y(25) => MuxOutputs_3_25_port,
                           Y(24) => MuxOutputs_3_24_port, Y(23) => 
                           MuxOutputs_3_23_port, Y(22) => MuxOutputs_3_22_port,
                           Y(21) => MuxOutputs_3_21_port, Y(20) => 
                           MuxOutputs_3_20_port, Y(19) => MuxOutputs_3_19_port,
                           Y(18) => MuxOutputs_3_18_port, Y(17) => 
                           MuxOutputs_3_17_port, Y(16) => MuxOutputs_3_16_port,
                           Y(15) => MuxOutputs_3_15_port, Y(14) => 
                           MuxOutputs_3_14_port, Y(13) => MuxOutputs_3_13_port,
                           Y(12) => MuxOutputs_3_12_port, Y(11) => 
                           MuxOutputs_3_11_port, Y(10) => MuxOutputs_3_10_port,
                           Y(9) => MuxOutputs_3_9_port, Y(8) => 
                           MuxOutputs_3_8_port, Y(7) => MuxOutputs_3_7_port, 
                           Y(6) => MuxOutputs_3_6_port, Y(5) => 
                           MuxOutputs_3_5_port, Y(4) => MuxOutputs_3_4_port, 
                           Y(3) => MuxOutputs_3_3_port, Y(2) => 
                           MuxOutputs_3_2_port, Y(1) => MuxOutputs_3_1_port, 
                           Y(0) => MuxOutputs_3_0_port);
   encoderI_4 : encoder_12 port map( pieceofB(2) => B(9), pieceofB(1) => B(8), 
                           pieceofB(0) => B(7), sel(2) => sel_4_2_port, sel(1) 
                           => sel_4_1_port, sel(0) => sel_4_0_port);
   MUXI_4 : MUX51_MuxNbit64_12 port map( zeroSignal(63) => X_Logic0_port, 
                           zeroSignal(62) => X_Logic0_port, zeroSignal(61) => 
                           X_Logic0_port, zeroSignal(60) => X_Logic0_port, 
                           zeroSignal(59) => X_Logic0_port, zeroSignal(58) => 
                           X_Logic0_port, zeroSignal(57) => X_Logic0_port, 
                           zeroSignal(56) => X_Logic0_port, zeroSignal(55) => 
                           X_Logic0_port, zeroSignal(54) => X_Logic0_port, 
                           zeroSignal(53) => X_Logic0_port, zeroSignal(52) => 
                           X_Logic0_port, zeroSignal(51) => X_Logic0_port, 
                           zeroSignal(50) => X_Logic0_port, zeroSignal(49) => 
                           X_Logic0_port, zeroSignal(48) => X_Logic0_port, 
                           zeroSignal(47) => X_Logic0_port, zeroSignal(46) => 
                           X_Logic0_port, zeroSignal(45) => X_Logic0_port, 
                           zeroSignal(44) => X_Logic0_port, zeroSignal(43) => 
                           X_Logic0_port, zeroSignal(42) => X_Logic0_port, 
                           zeroSignal(41) => X_Logic0_port, zeroSignal(40) => 
                           X_Logic0_port, zeroSignal(39) => X_Logic0_port, 
                           zeroSignal(38) => X_Logic0_port, zeroSignal(37) => 
                           X_Logic0_port, zeroSignal(36) => X_Logic0_port, 
                           zeroSignal(35) => X_Logic0_port, zeroSignal(34) => 
                           X_Logic0_port, zeroSignal(33) => X_Logic0_port, 
                           zeroSignal(32) => X_Logic0_port, zeroSignal(31) => 
                           X_Logic0_port, zeroSignal(30) => X_Logic0_port, 
                           zeroSignal(29) => X_Logic0_port, zeroSignal(28) => 
                           X_Logic0_port, zeroSignal(27) => X_Logic0_port, 
                           zeroSignal(26) => X_Logic0_port, zeroSignal(25) => 
                           X_Logic0_port, zeroSignal(24) => X_Logic0_port, 
                           zeroSignal(23) => X_Logic0_port, zeroSignal(22) => 
                           X_Logic0_port, zeroSignal(21) => X_Logic0_port, 
                           zeroSignal(20) => X_Logic0_port, zeroSignal(19) => 
                           X_Logic0_port, zeroSignal(18) => X_Logic0_port, 
                           zeroSignal(17) => X_Logic0_port, zeroSignal(16) => 
                           X_Logic0_port, zeroSignal(15) => X_Logic0_port, 
                           zeroSignal(14) => X_Logic0_port, zeroSignal(13) => 
                           X_Logic0_port, zeroSignal(12) => X_Logic0_port, 
                           zeroSignal(11) => X_Logic0_port, zeroSignal(10) => 
                           X_Logic0_port, zeroSignal(9) => X_Logic0_port, 
                           zeroSignal(8) => X_Logic0_port, zeroSignal(7) => 
                           X_Logic0_port, zeroSignal(6) => X_Logic0_port, 
                           zeroSignal(5) => X_Logic0_port, zeroSignal(4) => 
                           X_Logic0_port, zeroSignal(3) => X_Logic0_port, 
                           zeroSignal(2) => X_Logic0_port, zeroSignal(1) => 
                           X_Logic0_port, zeroSignal(0) => X_Logic0_port, 
                           A_signal(63) => positive_inputs_8_63_port, 
                           A_signal(62) => positive_inputs_8_62_port, 
                           A_signal(61) => positive_inputs_8_61_port, 
                           A_signal(60) => positive_inputs_8_60_port, 
                           A_signal(59) => positive_inputs_8_59_port, 
                           A_signal(58) => positive_inputs_8_58_port, 
                           A_signal(57) => positive_inputs_8_57_port, 
                           A_signal(56) => positive_inputs_8_56_port, 
                           A_signal(55) => positive_inputs_8_55_port, 
                           A_signal(54) => positive_inputs_8_54_port, 
                           A_signal(53) => positive_inputs_8_53_port, 
                           A_signal(52) => positive_inputs_8_52_port, 
                           A_signal(51) => positive_inputs_8_51_port, 
                           A_signal(50) => positive_inputs_8_50_port, 
                           A_signal(49) => positive_inputs_8_49_port, 
                           A_signal(48) => n65, A_signal(47) => 
                           positive_inputs_8_47_port, A_signal(46) => 
                           positive_inputs_8_46_port, A_signal(45) => 
                           positive_inputs_8_45_port, A_signal(44) => 
                           positive_inputs_8_44_port, A_signal(43) => 
                           positive_inputs_8_43_port, A_signal(42) => 
                           positive_inputs_8_42_port, A_signal(41) => 
                           positive_inputs_8_41_port, A_signal(40) => 
                           positive_inputs_8_40_port, A_signal(39) => 
                           positive_inputs_8_39_port, A_signal(38) => 
                           positive_inputs_8_38_port, A_signal(37) => 
                           positive_inputs_8_37_port, A_signal(36) => 
                           positive_inputs_8_36_port, A_signal(35) => 
                           positive_inputs_8_35_port, A_signal(34) => 
                           positive_inputs_8_34_port, A_signal(33) => 
                           positive_inputs_8_33_port, A_signal(32) => 
                           positive_inputs_8_32_port, A_signal(31) => 
                           positive_inputs_8_31_port, A_signal(30) => 
                           positive_inputs_8_30_port, A_signal(29) => 
                           positive_inputs_8_29_port, A_signal(28) => 
                           positive_inputs_8_28_port, A_signal(27) => 
                           positive_inputs_8_27_port, A_signal(26) => 
                           positive_inputs_8_26_port, A_signal(25) => 
                           positive_inputs_8_25_port, A_signal(24) => 
                           positive_inputs_8_24_port, A_signal(23) => 
                           positive_inputs_8_23_port, A_signal(22) => 
                           positive_inputs_8_22_port, A_signal(21) => 
                           positive_inputs_8_21_port, A_signal(20) => 
                           positive_inputs_8_20_port, A_signal(19) => 
                           positive_inputs_8_19_port, A_signal(18) => 
                           positive_inputs_8_18_port, A_signal(17) => 
                           positive_inputs_8_17_port, A_signal(16) => 
                           positive_inputs_8_16_port, A_signal(15) => 
                           positive_inputs_8_15_port, A_signal(14) => 
                           positive_inputs_8_14_port, A_signal(13) => 
                           positive_inputs_8_13_port, A_signal(12) => 
                           positive_inputs_8_12_port, A_signal(11) => 
                           positive_inputs_8_11_port, A_signal(10) => 
                           positive_inputs_8_10_port, A_signal(9) => 
                           positive_inputs_8_9_port, A_signal(8) => 
                           positive_inputs_8_8_port, A_signal(7) => 
                           positive_inputs_8_7_port, A_signal(6) => 
                           positive_inputs_8_6_port, A_signal(5) => 
                           positive_inputs_8_5_port, A_signal(4) => 
                           positive_inputs_8_4_port, A_signal(3) => 
                           positive_inputs_8_3_port, A_signal(2) => 
                           positive_inputs_8_2_port, A_signal(1) => 
                           positive_inputs_8_1_port, A_signal(0) => n9, 
                           A_neg(63) => negative_inputs_8_63_port, A_neg(62) =>
                           negative_inputs_8_62_port, A_neg(61) => 
                           negative_inputs_8_61_port, A_neg(60) => 
                           negative_inputs_8_60_port, A_neg(59) => 
                           negative_inputs_8_59_port, A_neg(58) => 
                           negative_inputs_8_58_port, A_neg(57) => 
                           negative_inputs_8_57_port, A_neg(56) => 
                           negative_inputs_8_56_port, A_neg(55) => 
                           negative_inputs_8_55_port, A_neg(54) => 
                           negative_inputs_8_54_port, A_neg(53) => 
                           negative_inputs_8_53_port, A_neg(52) => 
                           negative_inputs_8_52_port, A_neg(51) => 
                           negative_inputs_8_51_port, A_neg(50) => 
                           negative_inputs_8_50_port, A_neg(49) => 
                           negative_inputs_8_49_port, A_neg(48) => n153, 
                           A_neg(47) => negative_inputs_8_47_port, A_neg(46) =>
                           negative_inputs_8_46_port, A_neg(45) => 
                           negative_inputs_8_45_port, A_neg(44) => 
                           negative_inputs_8_44_port, A_neg(43) => 
                           negative_inputs_8_43_port, A_neg(42) => 
                           negative_inputs_8_42_port, A_neg(41) => 
                           negative_inputs_8_41_port, A_neg(40) => 
                           negative_inputs_8_40_port, A_neg(39) => 
                           negative_inputs_8_39_port, A_neg(38) => 
                           negative_inputs_8_38_port, A_neg(37) => 
                           negative_inputs_8_37_port, A_neg(36) => 
                           negative_inputs_8_36_port, A_neg(35) => 
                           negative_inputs_8_35_port, A_neg(34) => 
                           negative_inputs_8_34_port, A_neg(33) => 
                           negative_inputs_8_33_port, A_neg(32) => 
                           negative_inputs_8_32_port, A_neg(31) => 
                           negative_inputs_8_31_port, A_neg(30) => 
                           negative_inputs_8_30_port, A_neg(29) => 
                           negative_inputs_8_29_port, A_neg(28) => 
                           negative_inputs_8_28_port, A_neg(27) => 
                           negative_inputs_8_27_port, A_neg(26) => 
                           negative_inputs_8_26_port, A_neg(25) => 
                           negative_inputs_8_25_port, A_neg(24) => 
                           negative_inputs_8_24_port, A_neg(23) => 
                           negative_inputs_8_23_port, A_neg(22) => 
                           negative_inputs_8_22_port, A_neg(21) => 
                           negative_inputs_8_21_port, A_neg(20) => 
                           negative_inputs_8_20_port, A_neg(19) => 
                           negative_inputs_8_19_port, A_neg(18) => 
                           negative_inputs_8_18_port, A_neg(17) => 
                           negative_inputs_8_17_port, A_neg(16) => 
                           negative_inputs_8_16_port, A_neg(15) => 
                           negative_inputs_8_15_port, A_neg(14) => 
                           negative_inputs_8_14_port, A_neg(13) => 
                           negative_inputs_8_13_port, A_neg(12) => 
                           negative_inputs_8_12_port, A_neg(11) => 
                           negative_inputs_8_11_port, A_neg(10) => 
                           negative_inputs_8_10_port, A_neg(9) => 
                           negative_inputs_8_9_port, A_neg(8) => 
                           negative_inputs_8_8_port, A_neg(7) => 
                           negative_inputs_8_7_port, A_neg(6) => 
                           negative_inputs_8_6_port, A_neg(5) => 
                           negative_inputs_8_5_port, A_neg(4) => 
                           negative_inputs_8_4_port, A_neg(3) => 
                           negative_inputs_8_3_port, A_neg(2) => 
                           negative_inputs_8_2_port, A_neg(1) => 
                           negative_inputs_8_1_port, A_neg(0) => n9, 
                           A_shifted(63) => positive_inputs_9_63_port, 
                           A_shifted(62) => positive_inputs_9_62_port, 
                           A_shifted(61) => positive_inputs_9_61_port, 
                           A_shifted(60) => positive_inputs_9_60_port, 
                           A_shifted(59) => positive_inputs_9_59_port, 
                           A_shifted(58) => positive_inputs_9_58_port, 
                           A_shifted(57) => positive_inputs_9_57_port, 
                           A_shifted(56) => positive_inputs_9_56_port, 
                           A_shifted(55) => positive_inputs_9_55_port, 
                           A_shifted(54) => positive_inputs_9_54_port, 
                           A_shifted(53) => positive_inputs_9_53_port, 
                           A_shifted(52) => positive_inputs_9_52_port, 
                           A_shifted(51) => positive_inputs_9_51_port, 
                           A_shifted(50) => positive_inputs_9_50_port, 
                           A_shifted(49) => positive_inputs_9_49_port, 
                           A_shifted(48) => n64, A_shifted(47) => 
                           positive_inputs_9_47_port, A_shifted(46) => 
                           positive_inputs_9_46_port, A_shifted(45) => 
                           positive_inputs_9_45_port, A_shifted(44) => 
                           positive_inputs_9_44_port, A_shifted(43) => 
                           positive_inputs_9_43_port, A_shifted(42) => 
                           positive_inputs_9_42_port, A_shifted(41) => 
                           positive_inputs_9_41_port, A_shifted(40) => 
                           positive_inputs_9_40_port, A_shifted(39) => 
                           positive_inputs_9_39_port, A_shifted(38) => 
                           positive_inputs_9_38_port, A_shifted(37) => 
                           positive_inputs_9_37_port, A_shifted(36) => 
                           positive_inputs_9_36_port, A_shifted(35) => 
                           positive_inputs_9_35_port, A_shifted(34) => 
                           positive_inputs_9_34_port, A_shifted(33) => 
                           positive_inputs_9_33_port, A_shifted(32) => 
                           positive_inputs_9_32_port, A_shifted(31) => 
                           positive_inputs_9_31_port, A_shifted(30) => 
                           positive_inputs_9_30_port, A_shifted(29) => 
                           positive_inputs_9_29_port, A_shifted(28) => 
                           positive_inputs_9_28_port, A_shifted(27) => 
                           positive_inputs_9_27_port, A_shifted(26) => 
                           positive_inputs_9_26_port, A_shifted(25) => 
                           positive_inputs_9_25_port, A_shifted(24) => 
                           positive_inputs_9_24_port, A_shifted(23) => 
                           positive_inputs_9_23_port, A_shifted(22) => 
                           positive_inputs_9_22_port, A_shifted(21) => 
                           positive_inputs_9_21_port, A_shifted(20) => 
                           positive_inputs_9_20_port, A_shifted(19) => 
                           positive_inputs_9_19_port, A_shifted(18) => 
                           positive_inputs_9_18_port, A_shifted(17) => 
                           positive_inputs_9_17_port, A_shifted(16) => 
                           positive_inputs_9_16_port, A_shifted(15) => 
                           positive_inputs_9_15_port, A_shifted(14) => 
                           positive_inputs_9_14_port, A_shifted(13) => 
                           positive_inputs_9_13_port, A_shifted(12) => 
                           positive_inputs_9_12_port, A_shifted(11) => 
                           positive_inputs_9_11_port, A_shifted(10) => 
                           positive_inputs_9_10_port, A_shifted(9) => 
                           positive_inputs_9_9_port, A_shifted(8) => 
                           positive_inputs_9_8_port, A_shifted(7) => 
                           positive_inputs_9_7_port, A_shifted(6) => 
                           positive_inputs_9_6_port, A_shifted(5) => 
                           positive_inputs_9_5_port, A_shifted(4) => 
                           positive_inputs_9_4_port, A_shifted(3) => 
                           positive_inputs_9_3_port, A_shifted(2) => 
                           positive_inputs_9_2_port, A_shifted(1) => 
                           positive_inputs_9_1_port, A_shifted(0) => n9, 
                           A_neg_shifted(63) => negative_inputs_9_63_port, 
                           A_neg_shifted(62) => negative_inputs_9_62_port, 
                           A_neg_shifted(61) => negative_inputs_9_61_port, 
                           A_neg_shifted(60) => negative_inputs_9_60_port, 
                           A_neg_shifted(59) => negative_inputs_9_59_port, 
                           A_neg_shifted(58) => negative_inputs_9_58_port, 
                           A_neg_shifted(57) => negative_inputs_9_57_port, 
                           A_neg_shifted(56) => negative_inputs_9_56_port, 
                           A_neg_shifted(55) => negative_inputs_9_55_port, 
                           A_neg_shifted(54) => negative_inputs_9_54_port, 
                           A_neg_shifted(53) => negative_inputs_9_53_port, 
                           A_neg_shifted(52) => negative_inputs_9_52_port, 
                           A_neg_shifted(51) => negative_inputs_9_51_port, 
                           A_neg_shifted(50) => negative_inputs_9_50_port, 
                           A_neg_shifted(49) => negative_inputs_9_49_port, 
                           A_neg_shifted(48) => n152, A_neg_shifted(47) => 
                           negative_inputs_9_47_port, A_neg_shifted(46) => 
                           negative_inputs_9_46_port, A_neg_shifted(45) => 
                           negative_inputs_9_45_port, A_neg_shifted(44) => 
                           negative_inputs_9_44_port, A_neg_shifted(43) => 
                           negative_inputs_9_43_port, A_neg_shifted(42) => 
                           negative_inputs_9_42_port, A_neg_shifted(41) => 
                           negative_inputs_9_41_port, A_neg_shifted(40) => 
                           negative_inputs_9_40_port, A_neg_shifted(39) => 
                           negative_inputs_9_39_port, A_neg_shifted(38) => 
                           negative_inputs_9_38_port, A_neg_shifted(37) => 
                           negative_inputs_9_37_port, A_neg_shifted(36) => 
                           negative_inputs_9_36_port, A_neg_shifted(35) => 
                           negative_inputs_9_35_port, A_neg_shifted(34) => 
                           negative_inputs_9_34_port, A_neg_shifted(33) => 
                           negative_inputs_9_33_port, A_neg_shifted(32) => 
                           negative_inputs_9_32_port, A_neg_shifted(31) => 
                           negative_inputs_9_31_port, A_neg_shifted(30) => 
                           negative_inputs_9_30_port, A_neg_shifted(29) => 
                           negative_inputs_9_29_port, A_neg_shifted(28) => 
                           negative_inputs_9_28_port, A_neg_shifted(27) => 
                           negative_inputs_9_27_port, A_neg_shifted(26) => 
                           negative_inputs_9_26_port, A_neg_shifted(25) => 
                           negative_inputs_9_25_port, A_neg_shifted(24) => 
                           negative_inputs_9_24_port, A_neg_shifted(23) => 
                           negative_inputs_9_23_port, A_neg_shifted(22) => 
                           negative_inputs_9_22_port, A_neg_shifted(21) => 
                           negative_inputs_9_21_port, A_neg_shifted(20) => 
                           negative_inputs_9_20_port, A_neg_shifted(19) => 
                           negative_inputs_9_19_port, A_neg_shifted(18) => 
                           negative_inputs_9_18_port, A_neg_shifted(17) => 
                           negative_inputs_9_17_port, A_neg_shifted(16) => 
                           negative_inputs_9_16_port, A_neg_shifted(15) => 
                           negative_inputs_9_15_port, A_neg_shifted(14) => 
                           negative_inputs_9_14_port, A_neg_shifted(13) => 
                           negative_inputs_9_13_port, A_neg_shifted(12) => 
                           negative_inputs_9_12_port, A_neg_shifted(11) => 
                           negative_inputs_9_11_port, A_neg_shifted(10) => 
                           negative_inputs_9_10_port, A_neg_shifted(9) => 
                           negative_inputs_9_9_port, A_neg_shifted(8) => 
                           negative_inputs_9_8_port, A_neg_shifted(7) => 
                           negative_inputs_9_7_port, A_neg_shifted(6) => 
                           negative_inputs_9_6_port, A_neg_shifted(5) => 
                           negative_inputs_9_5_port, A_neg_shifted(4) => 
                           negative_inputs_9_4_port, A_neg_shifted(3) => 
                           negative_inputs_9_3_port, A_neg_shifted(2) => 
                           negative_inputs_9_2_port, A_neg_shifted(1) => 
                           negative_inputs_9_1_port, A_neg_shifted(0) => n9, 
                           Sel(2) => sel_4_2_port, Sel(1) => sel_4_1_port, 
                           Sel(0) => sel_4_0_port, Y(63) => 
                           MuxOutputs_4_63_port, Y(62) => MuxOutputs_4_62_port,
                           Y(61) => MuxOutputs_4_61_port, Y(60) => 
                           MuxOutputs_4_60_port, Y(59) => MuxOutputs_4_59_port,
                           Y(58) => MuxOutputs_4_58_port, Y(57) => 
                           MuxOutputs_4_57_port, Y(56) => MuxOutputs_4_56_port,
                           Y(55) => MuxOutputs_4_55_port, Y(54) => 
                           MuxOutputs_4_54_port, Y(53) => MuxOutputs_4_53_port,
                           Y(52) => MuxOutputs_4_52_port, Y(51) => 
                           MuxOutputs_4_51_port, Y(50) => MuxOutputs_4_50_port,
                           Y(49) => MuxOutputs_4_49_port, Y(48) => 
                           MuxOutputs_4_48_port, Y(47) => MuxOutputs_4_47_port,
                           Y(46) => MuxOutputs_4_46_port, Y(45) => 
                           MuxOutputs_4_45_port, Y(44) => MuxOutputs_4_44_port,
                           Y(43) => MuxOutputs_4_43_port, Y(42) => 
                           MuxOutputs_4_42_port, Y(41) => MuxOutputs_4_41_port,
                           Y(40) => MuxOutputs_4_40_port, Y(39) => 
                           MuxOutputs_4_39_port, Y(38) => MuxOutputs_4_38_port,
                           Y(37) => MuxOutputs_4_37_port, Y(36) => 
                           MuxOutputs_4_36_port, Y(35) => MuxOutputs_4_35_port,
                           Y(34) => MuxOutputs_4_34_port, Y(33) => 
                           MuxOutputs_4_33_port, Y(32) => MuxOutputs_4_32_port,
                           Y(31) => MuxOutputs_4_31_port, Y(30) => 
                           MuxOutputs_4_30_port, Y(29) => MuxOutputs_4_29_port,
                           Y(28) => MuxOutputs_4_28_port, Y(27) => 
                           MuxOutputs_4_27_port, Y(26) => MuxOutputs_4_26_port,
                           Y(25) => MuxOutputs_4_25_port, Y(24) => 
                           MuxOutputs_4_24_port, Y(23) => MuxOutputs_4_23_port,
                           Y(22) => MuxOutputs_4_22_port, Y(21) => 
                           MuxOutputs_4_21_port, Y(20) => MuxOutputs_4_20_port,
                           Y(19) => MuxOutputs_4_19_port, Y(18) => 
                           MuxOutputs_4_18_port, Y(17) => MuxOutputs_4_17_port,
                           Y(16) => MuxOutputs_4_16_port, Y(15) => 
                           MuxOutputs_4_15_port, Y(14) => MuxOutputs_4_14_port,
                           Y(13) => MuxOutputs_4_13_port, Y(12) => 
                           MuxOutputs_4_12_port, Y(11) => MuxOutputs_4_11_port,
                           Y(10) => MuxOutputs_4_10_port, Y(9) => 
                           MuxOutputs_4_9_port, Y(8) => MuxOutputs_4_8_port, 
                           Y(7) => MuxOutputs_4_7_port, Y(6) => 
                           MuxOutputs_4_6_port, Y(5) => MuxOutputs_4_5_port, 
                           Y(4) => MuxOutputs_4_4_port, Y(3) => 
                           MuxOutputs_4_3_port, Y(2) => MuxOutputs_4_2_port, 
                           Y(1) => MuxOutputs_4_1_port, Y(0) => 
                           MuxOutputs_4_0_port);
   encoderI_5 : encoder_11 port map( pieceofB(2) => B(11), pieceofB(1) => B(10)
                           , pieceofB(0) => B(9), sel(2) => sel_5_2_port, 
                           sel(1) => sel_5_1_port, sel(0) => sel_5_0_port);
   MUXI_5 : MUX51_MuxNbit64_11 port map( zeroSignal(63) => X_Logic0_port, 
                           zeroSignal(62) => X_Logic0_port, zeroSignal(61) => 
                           X_Logic0_port, zeroSignal(60) => X_Logic0_port, 
                           zeroSignal(59) => X_Logic0_port, zeroSignal(58) => 
                           X_Logic0_port, zeroSignal(57) => X_Logic0_port, 
                           zeroSignal(56) => X_Logic0_port, zeroSignal(55) => 
                           X_Logic0_port, zeroSignal(54) => X_Logic0_port, 
                           zeroSignal(53) => X_Logic0_port, zeroSignal(52) => 
                           X_Logic0_port, zeroSignal(51) => X_Logic0_port, 
                           zeroSignal(50) => X_Logic0_port, zeroSignal(49) => 
                           X_Logic0_port, zeroSignal(48) => X_Logic0_port, 
                           zeroSignal(47) => X_Logic0_port, zeroSignal(46) => 
                           X_Logic0_port, zeroSignal(45) => X_Logic0_port, 
                           zeroSignal(44) => X_Logic0_port, zeroSignal(43) => 
                           X_Logic0_port, zeroSignal(42) => X_Logic0_port, 
                           zeroSignal(41) => X_Logic0_port, zeroSignal(40) => 
                           X_Logic0_port, zeroSignal(39) => X_Logic0_port, 
                           zeroSignal(38) => X_Logic0_port, zeroSignal(37) => 
                           X_Logic0_port, zeroSignal(36) => X_Logic0_port, 
                           zeroSignal(35) => X_Logic0_port, zeroSignal(34) => 
                           X_Logic0_port, zeroSignal(33) => X_Logic0_port, 
                           zeroSignal(32) => X_Logic0_port, zeroSignal(31) => 
                           X_Logic0_port, zeroSignal(30) => X_Logic0_port, 
                           zeroSignal(29) => X_Logic0_port, zeroSignal(28) => 
                           X_Logic0_port, zeroSignal(27) => X_Logic0_port, 
                           zeroSignal(26) => X_Logic0_port, zeroSignal(25) => 
                           X_Logic0_port, zeroSignal(24) => X_Logic0_port, 
                           zeroSignal(23) => X_Logic0_port, zeroSignal(22) => 
                           X_Logic0_port, zeroSignal(21) => X_Logic0_port, 
                           zeroSignal(20) => X_Logic0_port, zeroSignal(19) => 
                           X_Logic0_port, zeroSignal(18) => X_Logic0_port, 
                           zeroSignal(17) => X_Logic0_port, zeroSignal(16) => 
                           X_Logic0_port, zeroSignal(15) => X_Logic0_port, 
                           zeroSignal(14) => X_Logic0_port, zeroSignal(13) => 
                           X_Logic0_port, zeroSignal(12) => X_Logic0_port, 
                           zeroSignal(11) => X_Logic0_port, zeroSignal(10) => 
                           X_Logic0_port, zeroSignal(9) => X_Logic0_port, 
                           zeroSignal(8) => X_Logic0_port, zeroSignal(7) => 
                           X_Logic0_port, zeroSignal(6) => X_Logic0_port, 
                           zeroSignal(5) => X_Logic0_port, zeroSignal(4) => 
                           X_Logic0_port, zeroSignal(3) => X_Logic0_port, 
                           zeroSignal(2) => X_Logic0_port, zeroSignal(1) => 
                           X_Logic0_port, zeroSignal(0) => X_Logic0_port, 
                           A_signal(63) => positive_inputs_10_63_port, 
                           A_signal(62) => positive_inputs_10_62_port, 
                           A_signal(61) => positive_inputs_10_61_port, 
                           A_signal(60) => positive_inputs_10_60_port, 
                           A_signal(59) => positive_inputs_10_59_port, 
                           A_signal(58) => positive_inputs_10_58_port, 
                           A_signal(57) => positive_inputs_10_57_port, 
                           A_signal(56) => positive_inputs_10_56_port, 
                           A_signal(55) => positive_inputs_10_55_port, 
                           A_signal(54) => positive_inputs_10_54_port, 
                           A_signal(53) => positive_inputs_10_53_port, 
                           A_signal(52) => positive_inputs_10_52_port, 
                           A_signal(51) => positive_inputs_10_51_port, 
                           A_signal(50) => positive_inputs_10_50_port, 
                           A_signal(49) => positive_inputs_10_49_port, 
                           A_signal(48) => n63, A_signal(47) => 
                           positive_inputs_10_47_port, A_signal(46) => 
                           positive_inputs_10_46_port, A_signal(45) => 
                           positive_inputs_10_45_port, A_signal(44) => 
                           positive_inputs_10_44_port, A_signal(43) => 
                           positive_inputs_10_43_port, A_signal(42) => 
                           positive_inputs_10_42_port, A_signal(41) => 
                           positive_inputs_10_41_port, A_signal(40) => 
                           positive_inputs_10_40_port, A_signal(39) => 
                           positive_inputs_10_39_port, A_signal(38) => 
                           positive_inputs_10_38_port, A_signal(37) => 
                           positive_inputs_10_37_port, A_signal(36) => 
                           positive_inputs_10_36_port, A_signal(35) => 
                           positive_inputs_10_35_port, A_signal(34) => 
                           positive_inputs_10_34_port, A_signal(33) => 
                           positive_inputs_10_33_port, A_signal(32) => 
                           positive_inputs_10_32_port, A_signal(31) => 
                           positive_inputs_10_31_port, A_signal(30) => 
                           positive_inputs_10_30_port, A_signal(29) => 
                           positive_inputs_10_29_port, A_signal(28) => 
                           positive_inputs_10_28_port, A_signal(27) => 
                           positive_inputs_10_27_port, A_signal(26) => 
                           positive_inputs_10_26_port, A_signal(25) => 
                           positive_inputs_10_25_port, A_signal(24) => 
                           positive_inputs_10_24_port, A_signal(23) => 
                           positive_inputs_10_23_port, A_signal(22) => 
                           positive_inputs_10_22_port, A_signal(21) => 
                           positive_inputs_10_21_port, A_signal(20) => 
                           positive_inputs_10_20_port, A_signal(19) => 
                           positive_inputs_10_19_port, A_signal(18) => 
                           positive_inputs_10_18_port, A_signal(17) => 
                           positive_inputs_10_17_port, A_signal(16) => 
                           positive_inputs_10_16_port, A_signal(15) => 
                           positive_inputs_10_15_port, A_signal(14) => 
                           positive_inputs_10_14_port, A_signal(13) => 
                           positive_inputs_10_13_port, A_signal(12) => 
                           positive_inputs_10_12_port, A_signal(11) => 
                           positive_inputs_10_11_port, A_signal(10) => 
                           positive_inputs_10_10_port, A_signal(9) => 
                           positive_inputs_10_9_port, A_signal(8) => 
                           positive_inputs_10_8_port, A_signal(7) => 
                           positive_inputs_10_7_port, A_signal(6) => 
                           positive_inputs_10_6_port, A_signal(5) => 
                           positive_inputs_10_5_port, A_signal(4) => 
                           positive_inputs_10_4_port, A_signal(3) => 
                           positive_inputs_10_3_port, A_signal(2) => 
                           positive_inputs_10_2_port, A_signal(1) => 
                           positive_inputs_10_1_port, A_signal(0) => n9, 
                           A_neg(63) => negative_inputs_10_63_port, A_neg(62) 
                           => negative_inputs_10_62_port, A_neg(61) => 
                           negative_inputs_10_61_port, A_neg(60) => 
                           negative_inputs_10_60_port, A_neg(59) => 
                           negative_inputs_10_59_port, A_neg(58) => 
                           negative_inputs_10_58_port, A_neg(57) => 
                           negative_inputs_10_57_port, A_neg(56) => 
                           negative_inputs_10_56_port, A_neg(55) => 
                           negative_inputs_10_55_port, A_neg(54) => 
                           negative_inputs_10_54_port, A_neg(53) => 
                           negative_inputs_10_53_port, A_neg(52) => 
                           negative_inputs_10_52_port, A_neg(51) => 
                           negative_inputs_10_51_port, A_neg(50) => 
                           negative_inputs_10_50_port, A_neg(49) => 
                           negative_inputs_10_49_port, A_neg(48) => n150, 
                           A_neg(47) => negative_inputs_10_47_port, A_neg(46) 
                           => negative_inputs_10_46_port, A_neg(45) => 
                           negative_inputs_10_45_port, A_neg(44) => 
                           negative_inputs_10_44_port, A_neg(43) => 
                           negative_inputs_10_43_port, A_neg(42) => 
                           negative_inputs_10_42_port, A_neg(41) => 
                           negative_inputs_10_41_port, A_neg(40) => 
                           negative_inputs_10_40_port, A_neg(39) => 
                           negative_inputs_10_39_port, A_neg(38) => 
                           negative_inputs_10_38_port, A_neg(37) => 
                           negative_inputs_10_37_port, A_neg(36) => 
                           negative_inputs_10_36_port, A_neg(35) => 
                           negative_inputs_10_35_port, A_neg(34) => 
                           negative_inputs_10_34_port, A_neg(33) => 
                           negative_inputs_10_33_port, A_neg(32) => 
                           negative_inputs_10_32_port, A_neg(31) => 
                           negative_inputs_10_31_port, A_neg(30) => 
                           negative_inputs_10_30_port, A_neg(29) => 
                           negative_inputs_10_29_port, A_neg(28) => 
                           negative_inputs_10_28_port, A_neg(27) => 
                           negative_inputs_10_27_port, A_neg(26) => 
                           negative_inputs_10_26_port, A_neg(25) => 
                           negative_inputs_10_25_port, A_neg(24) => 
                           negative_inputs_10_24_port, A_neg(23) => 
                           negative_inputs_10_23_port, A_neg(22) => 
                           negative_inputs_10_22_port, A_neg(21) => 
                           negative_inputs_10_21_port, A_neg(20) => 
                           negative_inputs_10_20_port, A_neg(19) => 
                           negative_inputs_10_19_port, A_neg(18) => 
                           negative_inputs_10_18_port, A_neg(17) => 
                           negative_inputs_10_17_port, A_neg(16) => 
                           negative_inputs_10_16_port, A_neg(15) => 
                           negative_inputs_10_15_port, A_neg(14) => 
                           negative_inputs_10_14_port, A_neg(13) => 
                           negative_inputs_10_13_port, A_neg(12) => 
                           negative_inputs_10_12_port, A_neg(11) => 
                           negative_inputs_10_11_port, A_neg(10) => 
                           negative_inputs_10_10_port, A_neg(9) => 
                           negative_inputs_10_9_port, A_neg(8) => 
                           negative_inputs_10_8_port, A_neg(7) => 
                           negative_inputs_10_7_port, A_neg(6) => 
                           negative_inputs_10_6_port, A_neg(5) => 
                           negative_inputs_10_5_port, A_neg(4) => 
                           negative_inputs_10_4_port, A_neg(3) => 
                           negative_inputs_10_3_port, A_neg(2) => 
                           negative_inputs_10_2_port, A_neg(1) => 
                           negative_inputs_10_1_port, A_neg(0) => n9, 
                           A_shifted(63) => positive_inputs_11_63_port, 
                           A_shifted(62) => positive_inputs_11_62_port, 
                           A_shifted(61) => positive_inputs_11_61_port, 
                           A_shifted(60) => positive_inputs_11_60_port, 
                           A_shifted(59) => positive_inputs_11_59_port, 
                           A_shifted(58) => positive_inputs_11_58_port, 
                           A_shifted(57) => positive_inputs_11_57_port, 
                           A_shifted(56) => positive_inputs_11_56_port, 
                           A_shifted(55) => positive_inputs_11_55_port, 
                           A_shifted(54) => positive_inputs_11_54_port, 
                           A_shifted(53) => positive_inputs_11_53_port, 
                           A_shifted(52) => positive_inputs_11_52_port, 
                           A_shifted(51) => positive_inputs_11_51_port, 
                           A_shifted(50) => positive_inputs_11_50_port, 
                           A_shifted(49) => positive_inputs_11_49_port, 
                           A_shifted(48) => n62, A_shifted(47) => 
                           positive_inputs_11_47_port, A_shifted(46) => 
                           positive_inputs_11_46_port, A_shifted(45) => 
                           positive_inputs_11_45_port, A_shifted(44) => 
                           positive_inputs_11_44_port, A_shifted(43) => 
                           positive_inputs_11_43_port, A_shifted(42) => 
                           positive_inputs_11_42_port, A_shifted(41) => 
                           positive_inputs_11_41_port, A_shifted(40) => 
                           positive_inputs_11_40_port, A_shifted(39) => 
                           positive_inputs_11_39_port, A_shifted(38) => 
                           positive_inputs_11_38_port, A_shifted(37) => 
                           positive_inputs_11_37_port, A_shifted(36) => 
                           positive_inputs_11_36_port, A_shifted(35) => 
                           positive_inputs_11_35_port, A_shifted(34) => 
                           positive_inputs_11_34_port, A_shifted(33) => 
                           positive_inputs_11_33_port, A_shifted(32) => 
                           positive_inputs_11_32_port, A_shifted(31) => 
                           positive_inputs_11_31_port, A_shifted(30) => 
                           positive_inputs_11_30_port, A_shifted(29) => 
                           positive_inputs_11_29_port, A_shifted(28) => 
                           positive_inputs_11_28_port, A_shifted(27) => 
                           positive_inputs_11_27_port, A_shifted(26) => 
                           positive_inputs_11_26_port, A_shifted(25) => 
                           positive_inputs_11_25_port, A_shifted(24) => 
                           positive_inputs_11_24_port, A_shifted(23) => 
                           positive_inputs_11_23_port, A_shifted(22) => 
                           positive_inputs_11_22_port, A_shifted(21) => 
                           positive_inputs_11_21_port, A_shifted(20) => 
                           positive_inputs_11_20_port, A_shifted(19) => 
                           positive_inputs_11_19_port, A_shifted(18) => 
                           positive_inputs_11_18_port, A_shifted(17) => 
                           positive_inputs_11_17_port, A_shifted(16) => 
                           positive_inputs_11_16_port, A_shifted(15) => 
                           positive_inputs_11_15_port, A_shifted(14) => 
                           positive_inputs_11_14_port, A_shifted(13) => 
                           positive_inputs_11_13_port, A_shifted(12) => 
                           positive_inputs_11_12_port, A_shifted(11) => 
                           positive_inputs_11_11_port, A_shifted(10) => 
                           positive_inputs_11_10_port, A_shifted(9) => 
                           positive_inputs_11_9_port, A_shifted(8) => 
                           positive_inputs_11_8_port, A_shifted(7) => 
                           positive_inputs_11_7_port, A_shifted(6) => 
                           positive_inputs_11_6_port, A_shifted(5) => 
                           positive_inputs_11_5_port, A_shifted(4) => 
                           positive_inputs_11_4_port, A_shifted(3) => 
                           positive_inputs_11_3_port, A_shifted(2) => 
                           positive_inputs_11_2_port, A_shifted(1) => 
                           positive_inputs_11_1_port, A_shifted(0) => n9, 
                           A_neg_shifted(63) => negative_inputs_11_63_port, 
                           A_neg_shifted(62) => negative_inputs_11_62_port, 
                           A_neg_shifted(61) => negative_inputs_11_61_port, 
                           A_neg_shifted(60) => negative_inputs_11_60_port, 
                           A_neg_shifted(59) => negative_inputs_11_59_port, 
                           A_neg_shifted(58) => negative_inputs_11_58_port, 
                           A_neg_shifted(57) => negative_inputs_11_57_port, 
                           A_neg_shifted(56) => negative_inputs_11_56_port, 
                           A_neg_shifted(55) => negative_inputs_11_55_port, 
                           A_neg_shifted(54) => negative_inputs_11_54_port, 
                           A_neg_shifted(53) => negative_inputs_11_53_port, 
                           A_neg_shifted(52) => negative_inputs_11_52_port, 
                           A_neg_shifted(51) => negative_inputs_11_51_port, 
                           A_neg_shifted(50) => negative_inputs_11_50_port, 
                           A_neg_shifted(49) => negative_inputs_11_49_port, 
                           A_neg_shifted(48) => n148, A_neg_shifted(47) => 
                           negative_inputs_11_47_port, A_neg_shifted(46) => 
                           negative_inputs_11_46_port, A_neg_shifted(45) => 
                           negative_inputs_11_45_port, A_neg_shifted(44) => 
                           negative_inputs_11_44_port, A_neg_shifted(43) => 
                           negative_inputs_11_43_port, A_neg_shifted(42) => 
                           negative_inputs_11_42_port, A_neg_shifted(41) => 
                           negative_inputs_11_41_port, A_neg_shifted(40) => 
                           negative_inputs_11_40_port, A_neg_shifted(39) => 
                           negative_inputs_11_39_port, A_neg_shifted(38) => 
                           negative_inputs_11_38_port, A_neg_shifted(37) => 
                           negative_inputs_11_37_port, A_neg_shifted(36) => 
                           negative_inputs_11_36_port, A_neg_shifted(35) => 
                           negative_inputs_11_35_port, A_neg_shifted(34) => 
                           negative_inputs_11_34_port, A_neg_shifted(33) => 
                           negative_inputs_11_33_port, A_neg_shifted(32) => 
                           negative_inputs_11_32_port, A_neg_shifted(31) => 
                           negative_inputs_11_31_port, A_neg_shifted(30) => 
                           negative_inputs_11_30_port, A_neg_shifted(29) => 
                           negative_inputs_11_29_port, A_neg_shifted(28) => 
                           negative_inputs_11_28_port, A_neg_shifted(27) => 
                           negative_inputs_11_27_port, A_neg_shifted(26) => 
                           negative_inputs_11_26_port, A_neg_shifted(25) => 
                           negative_inputs_11_25_port, A_neg_shifted(24) => 
                           negative_inputs_11_24_port, A_neg_shifted(23) => 
                           negative_inputs_11_23_port, A_neg_shifted(22) => 
                           negative_inputs_11_22_port, A_neg_shifted(21) => 
                           negative_inputs_11_21_port, A_neg_shifted(20) => 
                           negative_inputs_11_20_port, A_neg_shifted(19) => 
                           negative_inputs_11_19_port, A_neg_shifted(18) => 
                           negative_inputs_11_18_port, A_neg_shifted(17) => 
                           negative_inputs_11_17_port, A_neg_shifted(16) => 
                           negative_inputs_11_16_port, A_neg_shifted(15) => 
                           negative_inputs_11_15_port, A_neg_shifted(14) => 
                           negative_inputs_11_14_port, A_neg_shifted(13) => 
                           negative_inputs_11_13_port, A_neg_shifted(12) => 
                           negative_inputs_11_12_port, A_neg_shifted(11) => 
                           negative_inputs_11_11_port, A_neg_shifted(10) => 
                           negative_inputs_11_10_port, A_neg_shifted(9) => 
                           negative_inputs_11_9_port, A_neg_shifted(8) => 
                           negative_inputs_11_8_port, A_neg_shifted(7) => 
                           negative_inputs_11_7_port, A_neg_shifted(6) => 
                           negative_inputs_11_6_port, A_neg_shifted(5) => 
                           negative_inputs_11_5_port, A_neg_shifted(4) => 
                           negative_inputs_11_4_port, A_neg_shifted(3) => 
                           negative_inputs_11_3_port, A_neg_shifted(2) => 
                           negative_inputs_11_2_port, A_neg_shifted(1) => 
                           negative_inputs_11_1_port, A_neg_shifted(0) => n9, 
                           Sel(2) => sel_5_2_port, Sel(1) => sel_5_1_port, 
                           Sel(0) => sel_5_0_port, Y(63) => 
                           MuxOutputs_5_63_port, Y(62) => MuxOutputs_5_62_port,
                           Y(61) => MuxOutputs_5_61_port, Y(60) => 
                           MuxOutputs_5_60_port, Y(59) => MuxOutputs_5_59_port,
                           Y(58) => MuxOutputs_5_58_port, Y(57) => 
                           MuxOutputs_5_57_port, Y(56) => MuxOutputs_5_56_port,
                           Y(55) => MuxOutputs_5_55_port, Y(54) => 
                           MuxOutputs_5_54_port, Y(53) => MuxOutputs_5_53_port,
                           Y(52) => MuxOutputs_5_52_port, Y(51) => 
                           MuxOutputs_5_51_port, Y(50) => MuxOutputs_5_50_port,
                           Y(49) => MuxOutputs_5_49_port, Y(48) => 
                           MuxOutputs_5_48_port, Y(47) => MuxOutputs_5_47_port,
                           Y(46) => MuxOutputs_5_46_port, Y(45) => 
                           MuxOutputs_5_45_port, Y(44) => MuxOutputs_5_44_port,
                           Y(43) => MuxOutputs_5_43_port, Y(42) => 
                           MuxOutputs_5_42_port, Y(41) => MuxOutputs_5_41_port,
                           Y(40) => MuxOutputs_5_40_port, Y(39) => 
                           MuxOutputs_5_39_port, Y(38) => MuxOutputs_5_38_port,
                           Y(37) => MuxOutputs_5_37_port, Y(36) => 
                           MuxOutputs_5_36_port, Y(35) => MuxOutputs_5_35_port,
                           Y(34) => MuxOutputs_5_34_port, Y(33) => 
                           MuxOutputs_5_33_port, Y(32) => MuxOutputs_5_32_port,
                           Y(31) => MuxOutputs_5_31_port, Y(30) => 
                           MuxOutputs_5_30_port, Y(29) => MuxOutputs_5_29_port,
                           Y(28) => MuxOutputs_5_28_port, Y(27) => 
                           MuxOutputs_5_27_port, Y(26) => MuxOutputs_5_26_port,
                           Y(25) => MuxOutputs_5_25_port, Y(24) => 
                           MuxOutputs_5_24_port, Y(23) => MuxOutputs_5_23_port,
                           Y(22) => MuxOutputs_5_22_port, Y(21) => 
                           MuxOutputs_5_21_port, Y(20) => MuxOutputs_5_20_port,
                           Y(19) => MuxOutputs_5_19_port, Y(18) => 
                           MuxOutputs_5_18_port, Y(17) => MuxOutputs_5_17_port,
                           Y(16) => MuxOutputs_5_16_port, Y(15) => 
                           MuxOutputs_5_15_port, Y(14) => MuxOutputs_5_14_port,
                           Y(13) => MuxOutputs_5_13_port, Y(12) => 
                           MuxOutputs_5_12_port, Y(11) => MuxOutputs_5_11_port,
                           Y(10) => MuxOutputs_5_10_port, Y(9) => 
                           MuxOutputs_5_9_port, Y(8) => MuxOutputs_5_8_port, 
                           Y(7) => MuxOutputs_5_7_port, Y(6) => 
                           MuxOutputs_5_6_port, Y(5) => MuxOutputs_5_5_port, 
                           Y(4) => MuxOutputs_5_4_port, Y(3) => 
                           MuxOutputs_5_3_port, Y(2) => MuxOutputs_5_2_port, 
                           Y(1) => MuxOutputs_5_1_port, Y(0) => 
                           MuxOutputs_5_0_port);
   encoderI_6 : encoder_10 port map( pieceofB(2) => B(13), pieceofB(1) => B(12)
                           , pieceofB(0) => B(11), sel(2) => sel_6_2_port, 
                           sel(1) => sel_6_1_port, sel(0) => sel_6_0_port);
   MUXI_6 : MUX51_MuxNbit64_10 port map( zeroSignal(63) => X_Logic0_port, 
                           zeroSignal(62) => X_Logic0_port, zeroSignal(61) => 
                           X_Logic0_port, zeroSignal(60) => X_Logic0_port, 
                           zeroSignal(59) => X_Logic0_port, zeroSignal(58) => 
                           X_Logic0_port, zeroSignal(57) => X_Logic0_port, 
                           zeroSignal(56) => X_Logic0_port, zeroSignal(55) => 
                           X_Logic0_port, zeroSignal(54) => X_Logic0_port, 
                           zeroSignal(53) => X_Logic0_port, zeroSignal(52) => 
                           X_Logic0_port, zeroSignal(51) => X_Logic0_port, 
                           zeroSignal(50) => X_Logic0_port, zeroSignal(49) => 
                           X_Logic0_port, zeroSignal(48) => X_Logic0_port, 
                           zeroSignal(47) => X_Logic0_port, zeroSignal(46) => 
                           X_Logic0_port, zeroSignal(45) => X_Logic0_port, 
                           zeroSignal(44) => X_Logic0_port, zeroSignal(43) => 
                           X_Logic0_port, zeroSignal(42) => X_Logic0_port, 
                           zeroSignal(41) => X_Logic0_port, zeroSignal(40) => 
                           X_Logic0_port, zeroSignal(39) => X_Logic0_port, 
                           zeroSignal(38) => X_Logic0_port, zeroSignal(37) => 
                           X_Logic0_port, zeroSignal(36) => X_Logic0_port, 
                           zeroSignal(35) => X_Logic0_port, zeroSignal(34) => 
                           X_Logic0_port, zeroSignal(33) => X_Logic0_port, 
                           zeroSignal(32) => X_Logic0_port, zeroSignal(31) => 
                           X_Logic0_port, zeroSignal(30) => X_Logic0_port, 
                           zeroSignal(29) => X_Logic0_port, zeroSignal(28) => 
                           X_Logic0_port, zeroSignal(27) => X_Logic0_port, 
                           zeroSignal(26) => X_Logic0_port, zeroSignal(25) => 
                           X_Logic0_port, zeroSignal(24) => X_Logic0_port, 
                           zeroSignal(23) => X_Logic0_port, zeroSignal(22) => 
                           X_Logic0_port, zeroSignal(21) => X_Logic0_port, 
                           zeroSignal(20) => X_Logic0_port, zeroSignal(19) => 
                           X_Logic0_port, zeroSignal(18) => X_Logic0_port, 
                           zeroSignal(17) => X_Logic0_port, zeroSignal(16) => 
                           X_Logic0_port, zeroSignal(15) => X_Logic0_port, 
                           zeroSignal(14) => X_Logic0_port, zeroSignal(13) => 
                           X_Logic0_port, zeroSignal(12) => X_Logic0_port, 
                           zeroSignal(11) => X_Logic0_port, zeroSignal(10) => 
                           X_Logic0_port, zeroSignal(9) => X_Logic0_port, 
                           zeroSignal(8) => X_Logic0_port, zeroSignal(7) => 
                           X_Logic0_port, zeroSignal(6) => X_Logic0_port, 
                           zeroSignal(5) => X_Logic0_port, zeroSignal(4) => 
                           X_Logic0_port, zeroSignal(3) => X_Logic0_port, 
                           zeroSignal(2) => X_Logic0_port, zeroSignal(1) => 
                           X_Logic0_port, zeroSignal(0) => X_Logic0_port, 
                           A_signal(63) => positive_inputs_12_63_port, 
                           A_signal(62) => positive_inputs_12_62_port, 
                           A_signal(61) => positive_inputs_12_61_port, 
                           A_signal(60) => positive_inputs_12_60_port, 
                           A_signal(59) => positive_inputs_12_59_port, 
                           A_signal(58) => positive_inputs_12_58_port, 
                           A_signal(57) => positive_inputs_12_57_port, 
                           A_signal(56) => positive_inputs_12_56_port, 
                           A_signal(55) => positive_inputs_12_55_port, 
                           A_signal(54) => positive_inputs_12_54_port, 
                           A_signal(53) => positive_inputs_12_53_port, 
                           A_signal(52) => positive_inputs_12_52_port, 
                           A_signal(51) => positive_inputs_12_51_port, 
                           A_signal(50) => positive_inputs_12_50_port, 
                           A_signal(49) => positive_inputs_12_49_port, 
                           A_signal(48) => n61, A_signal(47) => 
                           positive_inputs_12_47_port, A_signal(46) => 
                           positive_inputs_12_46_port, A_signal(45) => 
                           positive_inputs_12_45_port, A_signal(44) => 
                           positive_inputs_12_44_port, A_signal(43) => 
                           positive_inputs_12_43_port, A_signal(42) => 
                           positive_inputs_12_42_port, A_signal(41) => 
                           positive_inputs_12_41_port, A_signal(40) => 
                           positive_inputs_12_40_port, A_signal(39) => 
                           positive_inputs_12_39_port, A_signal(38) => 
                           positive_inputs_12_38_port, A_signal(37) => 
                           positive_inputs_12_37_port, A_signal(36) => 
                           positive_inputs_12_36_port, A_signal(35) => 
                           positive_inputs_12_35_port, A_signal(34) => 
                           positive_inputs_12_34_port, A_signal(33) => 
                           positive_inputs_12_33_port, A_signal(32) => 
                           positive_inputs_12_32_port, A_signal(31) => 
                           positive_inputs_12_31_port, A_signal(30) => 
                           positive_inputs_12_30_port, A_signal(29) => 
                           positive_inputs_12_29_port, A_signal(28) => 
                           positive_inputs_12_28_port, A_signal(27) => 
                           positive_inputs_12_27_port, A_signal(26) => 
                           positive_inputs_12_26_port, A_signal(25) => 
                           positive_inputs_12_25_port, A_signal(24) => 
                           positive_inputs_12_24_port, A_signal(23) => 
                           positive_inputs_12_23_port, A_signal(22) => 
                           positive_inputs_12_22_port, A_signal(21) => 
                           positive_inputs_12_21_port, A_signal(20) => 
                           positive_inputs_12_20_port, A_signal(19) => 
                           positive_inputs_12_19_port, A_signal(18) => 
                           positive_inputs_12_18_port, A_signal(17) => 
                           positive_inputs_12_17_port, A_signal(16) => 
                           positive_inputs_12_16_port, A_signal(15) => 
                           positive_inputs_12_15_port, A_signal(14) => 
                           positive_inputs_12_14_port, A_signal(13) => 
                           positive_inputs_12_13_port, A_signal(12) => 
                           positive_inputs_12_12_port, A_signal(11) => 
                           positive_inputs_12_11_port, A_signal(10) => 
                           positive_inputs_12_10_port, A_signal(9) => 
                           positive_inputs_12_9_port, A_signal(8) => 
                           positive_inputs_12_8_port, A_signal(7) => 
                           positive_inputs_12_7_port, A_signal(6) => 
                           positive_inputs_12_6_port, A_signal(5) => 
                           positive_inputs_12_5_port, A_signal(4) => 
                           positive_inputs_12_4_port, A_signal(3) => 
                           positive_inputs_12_3_port, A_signal(2) => 
                           positive_inputs_12_2_port, A_signal(1) => 
                           positive_inputs_12_1_port, A_signal(0) => n9, 
                           A_neg(63) => negative_inputs_12_63_port, A_neg(62) 
                           => negative_inputs_12_62_port, A_neg(61) => 
                           negative_inputs_12_61_port, A_neg(60) => 
                           negative_inputs_12_60_port, A_neg(59) => 
                           negative_inputs_12_59_port, A_neg(58) => 
                           negative_inputs_12_58_port, A_neg(57) => 
                           negative_inputs_12_57_port, A_neg(56) => 
                           negative_inputs_12_56_port, A_neg(55) => 
                           negative_inputs_12_55_port, A_neg(54) => 
                           negative_inputs_12_54_port, A_neg(53) => 
                           negative_inputs_12_53_port, A_neg(52) => 
                           negative_inputs_12_52_port, A_neg(51) => 
                           negative_inputs_12_51_port, A_neg(50) => 
                           negative_inputs_12_50_port, A_neg(49) => 
                           negative_inputs_12_49_port, A_neg(48) => n146, 
                           A_neg(47) => negative_inputs_12_47_port, A_neg(46) 
                           => negative_inputs_12_46_port, A_neg(45) => 
                           negative_inputs_12_45_port, A_neg(44) => 
                           negative_inputs_12_44_port, A_neg(43) => 
                           negative_inputs_12_43_port, A_neg(42) => 
                           negative_inputs_12_42_port, A_neg(41) => 
                           negative_inputs_12_41_port, A_neg(40) => 
                           negative_inputs_12_40_port, A_neg(39) => 
                           negative_inputs_12_39_port, A_neg(38) => 
                           negative_inputs_12_38_port, A_neg(37) => 
                           negative_inputs_12_37_port, A_neg(36) => 
                           negative_inputs_12_36_port, A_neg(35) => 
                           negative_inputs_12_35_port, A_neg(34) => 
                           negative_inputs_12_34_port, A_neg(33) => 
                           negative_inputs_12_33_port, A_neg(32) => 
                           negative_inputs_12_32_port, A_neg(31) => 
                           negative_inputs_12_31_port, A_neg(30) => 
                           negative_inputs_12_30_port, A_neg(29) => 
                           negative_inputs_12_29_port, A_neg(28) => 
                           negative_inputs_12_28_port, A_neg(27) => 
                           negative_inputs_12_27_port, A_neg(26) => 
                           negative_inputs_12_26_port, A_neg(25) => 
                           negative_inputs_12_25_port, A_neg(24) => 
                           negative_inputs_12_24_port, A_neg(23) => 
                           negative_inputs_12_23_port, A_neg(22) => 
                           negative_inputs_12_22_port, A_neg(21) => 
                           negative_inputs_12_21_port, A_neg(20) => 
                           negative_inputs_12_20_port, A_neg(19) => 
                           negative_inputs_12_19_port, A_neg(18) => 
                           negative_inputs_12_18_port, A_neg(17) => 
                           negative_inputs_12_17_port, A_neg(16) => 
                           negative_inputs_12_16_port, A_neg(15) => 
                           negative_inputs_12_15_port, A_neg(14) => 
                           negative_inputs_12_14_port, A_neg(13) => 
                           negative_inputs_12_13_port, A_neg(12) => 
                           negative_inputs_12_12_port, A_neg(11) => 
                           negative_inputs_12_11_port, A_neg(10) => 
                           negative_inputs_12_10_port, A_neg(9) => 
                           negative_inputs_12_9_port, A_neg(8) => 
                           negative_inputs_12_8_port, A_neg(7) => 
                           negative_inputs_12_7_port, A_neg(6) => 
                           negative_inputs_12_6_port, A_neg(5) => 
                           negative_inputs_12_5_port, A_neg(4) => 
                           negative_inputs_12_4_port, A_neg(3) => 
                           negative_inputs_12_3_port, A_neg(2) => 
                           negative_inputs_12_2_port, A_neg(1) => 
                           negative_inputs_12_1_port, A_neg(0) => n9, 
                           A_shifted(63) => positive_inputs_13_63_port, 
                           A_shifted(62) => positive_inputs_13_62_port, 
                           A_shifted(61) => positive_inputs_13_61_port, 
                           A_shifted(60) => positive_inputs_13_60_port, 
                           A_shifted(59) => positive_inputs_13_59_port, 
                           A_shifted(58) => positive_inputs_13_58_port, 
                           A_shifted(57) => positive_inputs_13_57_port, 
                           A_shifted(56) => positive_inputs_13_56_port, 
                           A_shifted(55) => positive_inputs_13_55_port, 
                           A_shifted(54) => positive_inputs_13_54_port, 
                           A_shifted(53) => positive_inputs_13_53_port, 
                           A_shifted(52) => positive_inputs_13_52_port, 
                           A_shifted(51) => positive_inputs_13_51_port, 
                           A_shifted(50) => positive_inputs_13_50_port, 
                           A_shifted(49) => positive_inputs_13_49_port, 
                           A_shifted(48) => n60, A_shifted(47) => 
                           positive_inputs_13_47_port, A_shifted(46) => 
                           positive_inputs_13_46_port, A_shifted(45) => 
                           positive_inputs_13_45_port, A_shifted(44) => 
                           positive_inputs_13_44_port, A_shifted(43) => 
                           positive_inputs_13_43_port, A_shifted(42) => 
                           positive_inputs_13_42_port, A_shifted(41) => 
                           positive_inputs_13_41_port, A_shifted(40) => 
                           positive_inputs_13_40_port, A_shifted(39) => 
                           positive_inputs_13_39_port, A_shifted(38) => 
                           positive_inputs_13_38_port, A_shifted(37) => 
                           positive_inputs_13_37_port, A_shifted(36) => 
                           positive_inputs_13_36_port, A_shifted(35) => 
                           positive_inputs_13_35_port, A_shifted(34) => 
                           positive_inputs_13_34_port, A_shifted(33) => 
                           positive_inputs_13_33_port, A_shifted(32) => 
                           positive_inputs_13_32_port, A_shifted(31) => 
                           positive_inputs_13_31_port, A_shifted(30) => 
                           positive_inputs_13_30_port, A_shifted(29) => 
                           positive_inputs_13_29_port, A_shifted(28) => 
                           positive_inputs_13_28_port, A_shifted(27) => 
                           positive_inputs_13_27_port, A_shifted(26) => 
                           positive_inputs_13_26_port, A_shifted(25) => 
                           positive_inputs_13_25_port, A_shifted(24) => 
                           positive_inputs_13_24_port, A_shifted(23) => 
                           positive_inputs_13_23_port, A_shifted(22) => 
                           positive_inputs_13_22_port, A_shifted(21) => 
                           positive_inputs_13_21_port, A_shifted(20) => 
                           positive_inputs_13_20_port, A_shifted(19) => 
                           positive_inputs_13_19_port, A_shifted(18) => 
                           positive_inputs_13_18_port, A_shifted(17) => 
                           positive_inputs_13_17_port, A_shifted(16) => 
                           positive_inputs_13_16_port, A_shifted(15) => 
                           positive_inputs_13_15_port, A_shifted(14) => 
                           positive_inputs_13_14_port, A_shifted(13) => 
                           positive_inputs_13_13_port, A_shifted(12) => 
                           positive_inputs_13_12_port, A_shifted(11) => 
                           positive_inputs_13_11_port, A_shifted(10) => 
                           positive_inputs_13_10_port, A_shifted(9) => 
                           positive_inputs_13_9_port, A_shifted(8) => 
                           positive_inputs_13_8_port, A_shifted(7) => 
                           positive_inputs_13_7_port, A_shifted(6) => 
                           positive_inputs_13_6_port, A_shifted(5) => 
                           positive_inputs_13_5_port, A_shifted(4) => 
                           positive_inputs_13_4_port, A_shifted(3) => 
                           positive_inputs_13_3_port, A_shifted(2) => 
                           positive_inputs_13_2_port, A_shifted(1) => 
                           positive_inputs_13_1_port, A_shifted(0) => n9, 
                           A_neg_shifted(63) => negative_inputs_13_63_port, 
                           A_neg_shifted(62) => negative_inputs_13_62_port, 
                           A_neg_shifted(61) => negative_inputs_13_61_port, 
                           A_neg_shifted(60) => negative_inputs_13_60_port, 
                           A_neg_shifted(59) => negative_inputs_13_59_port, 
                           A_neg_shifted(58) => negative_inputs_13_58_port, 
                           A_neg_shifted(57) => negative_inputs_13_57_port, 
                           A_neg_shifted(56) => negative_inputs_13_56_port, 
                           A_neg_shifted(55) => negative_inputs_13_55_port, 
                           A_neg_shifted(54) => negative_inputs_13_54_port, 
                           A_neg_shifted(53) => negative_inputs_13_53_port, 
                           A_neg_shifted(52) => negative_inputs_13_52_port, 
                           A_neg_shifted(51) => negative_inputs_13_51_port, 
                           A_neg_shifted(50) => negative_inputs_13_50_port, 
                           A_neg_shifted(49) => negative_inputs_13_49_port, 
                           A_neg_shifted(48) => n144, A_neg_shifted(47) => 
                           negative_inputs_13_47_port, A_neg_shifted(46) => 
                           negative_inputs_13_46_port, A_neg_shifted(45) => 
                           negative_inputs_13_45_port, A_neg_shifted(44) => 
                           negative_inputs_13_44_port, A_neg_shifted(43) => 
                           negative_inputs_13_43_port, A_neg_shifted(42) => 
                           negative_inputs_13_42_port, A_neg_shifted(41) => 
                           negative_inputs_13_41_port, A_neg_shifted(40) => 
                           negative_inputs_13_40_port, A_neg_shifted(39) => 
                           negative_inputs_13_39_port, A_neg_shifted(38) => 
                           negative_inputs_13_38_port, A_neg_shifted(37) => 
                           negative_inputs_13_37_port, A_neg_shifted(36) => 
                           negative_inputs_13_36_port, A_neg_shifted(35) => 
                           negative_inputs_13_35_port, A_neg_shifted(34) => 
                           negative_inputs_13_34_port, A_neg_shifted(33) => 
                           negative_inputs_13_33_port, A_neg_shifted(32) => 
                           negative_inputs_13_32_port, A_neg_shifted(31) => 
                           negative_inputs_13_31_port, A_neg_shifted(30) => 
                           negative_inputs_13_30_port, A_neg_shifted(29) => 
                           negative_inputs_13_29_port, A_neg_shifted(28) => 
                           negative_inputs_13_28_port, A_neg_shifted(27) => 
                           negative_inputs_13_27_port, A_neg_shifted(26) => 
                           negative_inputs_13_26_port, A_neg_shifted(25) => 
                           negative_inputs_13_25_port, A_neg_shifted(24) => 
                           negative_inputs_13_24_port, A_neg_shifted(23) => 
                           negative_inputs_13_23_port, A_neg_shifted(22) => 
                           negative_inputs_13_22_port, A_neg_shifted(21) => 
                           negative_inputs_13_21_port, A_neg_shifted(20) => 
                           negative_inputs_13_20_port, A_neg_shifted(19) => 
                           negative_inputs_13_19_port, A_neg_shifted(18) => 
                           negative_inputs_13_18_port, A_neg_shifted(17) => 
                           negative_inputs_13_17_port, A_neg_shifted(16) => 
                           negative_inputs_13_16_port, A_neg_shifted(15) => 
                           negative_inputs_13_15_port, A_neg_shifted(14) => 
                           negative_inputs_13_14_port, A_neg_shifted(13) => 
                           negative_inputs_13_13_port, A_neg_shifted(12) => 
                           negative_inputs_13_12_port, A_neg_shifted(11) => 
                           negative_inputs_13_11_port, A_neg_shifted(10) => 
                           negative_inputs_13_10_port, A_neg_shifted(9) => 
                           negative_inputs_13_9_port, A_neg_shifted(8) => 
                           negative_inputs_13_8_port, A_neg_shifted(7) => 
                           negative_inputs_13_7_port, A_neg_shifted(6) => 
                           negative_inputs_13_6_port, A_neg_shifted(5) => 
                           negative_inputs_13_5_port, A_neg_shifted(4) => 
                           negative_inputs_13_4_port, A_neg_shifted(3) => 
                           negative_inputs_13_3_port, A_neg_shifted(2) => 
                           negative_inputs_13_2_port, A_neg_shifted(1) => 
                           negative_inputs_13_1_port, A_neg_shifted(0) => n9, 
                           Sel(2) => sel_6_2_port, Sel(1) => sel_6_1_port, 
                           Sel(0) => sel_6_0_port, Y(63) => 
                           MuxOutputs_6_63_port, Y(62) => MuxOutputs_6_62_port,
                           Y(61) => MuxOutputs_6_61_port, Y(60) => 
                           MuxOutputs_6_60_port, Y(59) => MuxOutputs_6_59_port,
                           Y(58) => MuxOutputs_6_58_port, Y(57) => 
                           MuxOutputs_6_57_port, Y(56) => MuxOutputs_6_56_port,
                           Y(55) => MuxOutputs_6_55_port, Y(54) => 
                           MuxOutputs_6_54_port, Y(53) => MuxOutputs_6_53_port,
                           Y(52) => MuxOutputs_6_52_port, Y(51) => 
                           MuxOutputs_6_51_port, Y(50) => MuxOutputs_6_50_port,
                           Y(49) => MuxOutputs_6_49_port, Y(48) => 
                           MuxOutputs_6_48_port, Y(47) => MuxOutputs_6_47_port,
                           Y(46) => MuxOutputs_6_46_port, Y(45) => 
                           MuxOutputs_6_45_port, Y(44) => MuxOutputs_6_44_port,
                           Y(43) => MuxOutputs_6_43_port, Y(42) => 
                           MuxOutputs_6_42_port, Y(41) => MuxOutputs_6_41_port,
                           Y(40) => MuxOutputs_6_40_port, Y(39) => 
                           MuxOutputs_6_39_port, Y(38) => MuxOutputs_6_38_port,
                           Y(37) => MuxOutputs_6_37_port, Y(36) => 
                           MuxOutputs_6_36_port, Y(35) => MuxOutputs_6_35_port,
                           Y(34) => MuxOutputs_6_34_port, Y(33) => 
                           MuxOutputs_6_33_port, Y(32) => MuxOutputs_6_32_port,
                           Y(31) => MuxOutputs_6_31_port, Y(30) => 
                           MuxOutputs_6_30_port, Y(29) => MuxOutputs_6_29_port,
                           Y(28) => MuxOutputs_6_28_port, Y(27) => 
                           MuxOutputs_6_27_port, Y(26) => MuxOutputs_6_26_port,
                           Y(25) => MuxOutputs_6_25_port, Y(24) => 
                           MuxOutputs_6_24_port, Y(23) => MuxOutputs_6_23_port,
                           Y(22) => MuxOutputs_6_22_port, Y(21) => 
                           MuxOutputs_6_21_port, Y(20) => MuxOutputs_6_20_port,
                           Y(19) => MuxOutputs_6_19_port, Y(18) => 
                           MuxOutputs_6_18_port, Y(17) => MuxOutputs_6_17_port,
                           Y(16) => MuxOutputs_6_16_port, Y(15) => 
                           MuxOutputs_6_15_port, Y(14) => MuxOutputs_6_14_port,
                           Y(13) => MuxOutputs_6_13_port, Y(12) => 
                           MuxOutputs_6_12_port, Y(11) => MuxOutputs_6_11_port,
                           Y(10) => MuxOutputs_6_10_port, Y(9) => 
                           MuxOutputs_6_9_port, Y(8) => MuxOutputs_6_8_port, 
                           Y(7) => MuxOutputs_6_7_port, Y(6) => 
                           MuxOutputs_6_6_port, Y(5) => MuxOutputs_6_5_port, 
                           Y(4) => MuxOutputs_6_4_port, Y(3) => 
                           MuxOutputs_6_3_port, Y(2) => MuxOutputs_6_2_port, 
                           Y(1) => MuxOutputs_6_1_port, Y(0) => 
                           MuxOutputs_6_0_port);
   encoderI_7 : encoder_9 port map( pieceofB(2) => B(15), pieceofB(1) => B(14),
                           pieceofB(0) => B(13), sel(2) => sel_7_2_port, sel(1)
                           => sel_7_1_port, sel(0) => sel_7_0_port);
   MUXI_7 : MUX51_MuxNbit64_9 port map( zeroSignal(63) => X_Logic0_port, 
                           zeroSignal(62) => X_Logic0_port, zeroSignal(61) => 
                           X_Logic0_port, zeroSignal(60) => X_Logic0_port, 
                           zeroSignal(59) => X_Logic0_port, zeroSignal(58) => 
                           X_Logic0_port, zeroSignal(57) => X_Logic0_port, 
                           zeroSignal(56) => X_Logic0_port, zeroSignal(55) => 
                           X_Logic0_port, zeroSignal(54) => X_Logic0_port, 
                           zeroSignal(53) => X_Logic0_port, zeroSignal(52) => 
                           X_Logic0_port, zeroSignal(51) => X_Logic0_port, 
                           zeroSignal(50) => X_Logic0_port, zeroSignal(49) => 
                           X_Logic0_port, zeroSignal(48) => X_Logic0_port, 
                           zeroSignal(47) => X_Logic0_port, zeroSignal(46) => 
                           X_Logic0_port, zeroSignal(45) => X_Logic0_port, 
                           zeroSignal(44) => X_Logic0_port, zeroSignal(43) => 
                           X_Logic0_port, zeroSignal(42) => X_Logic0_port, 
                           zeroSignal(41) => X_Logic0_port, zeroSignal(40) => 
                           X_Logic0_port, zeroSignal(39) => X_Logic0_port, 
                           zeroSignal(38) => X_Logic0_port, zeroSignal(37) => 
                           X_Logic0_port, zeroSignal(36) => X_Logic0_port, 
                           zeroSignal(35) => X_Logic0_port, zeroSignal(34) => 
                           X_Logic0_port, zeroSignal(33) => X_Logic0_port, 
                           zeroSignal(32) => X_Logic0_port, zeroSignal(31) => 
                           X_Logic0_port, zeroSignal(30) => X_Logic0_port, 
                           zeroSignal(29) => X_Logic0_port, zeroSignal(28) => 
                           X_Logic0_port, zeroSignal(27) => X_Logic0_port, 
                           zeroSignal(26) => X_Logic0_port, zeroSignal(25) => 
                           X_Logic0_port, zeroSignal(24) => X_Logic0_port, 
                           zeroSignal(23) => X_Logic0_port, zeroSignal(22) => 
                           X_Logic0_port, zeroSignal(21) => X_Logic0_port, 
                           zeroSignal(20) => X_Logic0_port, zeroSignal(19) => 
                           X_Logic0_port, zeroSignal(18) => X_Logic0_port, 
                           zeroSignal(17) => X_Logic0_port, zeroSignal(16) => 
                           X_Logic0_port, zeroSignal(15) => X_Logic0_port, 
                           zeroSignal(14) => X_Logic0_port, zeroSignal(13) => 
                           X_Logic0_port, zeroSignal(12) => X_Logic0_port, 
                           zeroSignal(11) => X_Logic0_port, zeroSignal(10) => 
                           X_Logic0_port, zeroSignal(9) => X_Logic0_port, 
                           zeroSignal(8) => X_Logic0_port, zeroSignal(7) => 
                           X_Logic0_port, zeroSignal(6) => X_Logic0_port, 
                           zeroSignal(5) => X_Logic0_port, zeroSignal(4) => 
                           X_Logic0_port, zeroSignal(3) => X_Logic0_port, 
                           zeroSignal(2) => X_Logic0_port, zeroSignal(1) => 
                           X_Logic0_port, zeroSignal(0) => X_Logic0_port, 
                           A_signal(63) => positive_inputs_14_63_port, 
                           A_signal(62) => positive_inputs_14_62_port, 
                           A_signal(61) => positive_inputs_14_61_port, 
                           A_signal(60) => positive_inputs_14_60_port, 
                           A_signal(59) => positive_inputs_14_59_port, 
                           A_signal(58) => positive_inputs_14_58_port, 
                           A_signal(57) => positive_inputs_14_57_port, 
                           A_signal(56) => positive_inputs_14_56_port, 
                           A_signal(55) => positive_inputs_14_55_port, 
                           A_signal(54) => positive_inputs_14_54_port, 
                           A_signal(53) => positive_inputs_14_53_port, 
                           A_signal(52) => positive_inputs_14_52_port, 
                           A_signal(51) => positive_inputs_14_51_port, 
                           A_signal(50) => positive_inputs_14_50_port, 
                           A_signal(49) => positive_inputs_14_49_port, 
                           A_signal(48) => n59, A_signal(47) => 
                           positive_inputs_14_47_port, A_signal(46) => 
                           positive_inputs_14_46_port, A_signal(45) => 
                           positive_inputs_14_45_port, A_signal(44) => 
                           positive_inputs_14_44_port, A_signal(43) => 
                           positive_inputs_14_43_port, A_signal(42) => 
                           positive_inputs_14_42_port, A_signal(41) => 
                           positive_inputs_14_41_port, A_signal(40) => 
                           positive_inputs_14_40_port, A_signal(39) => 
                           positive_inputs_14_39_port, A_signal(38) => 
                           positive_inputs_14_38_port, A_signal(37) => 
                           positive_inputs_14_37_port, A_signal(36) => 
                           positive_inputs_14_36_port, A_signal(35) => 
                           positive_inputs_14_35_port, A_signal(34) => 
                           positive_inputs_14_34_port, A_signal(33) => 
                           positive_inputs_14_33_port, A_signal(32) => 
                           positive_inputs_14_32_port, A_signal(31) => 
                           positive_inputs_14_31_port, A_signal(30) => 
                           positive_inputs_14_30_port, A_signal(29) => 
                           positive_inputs_14_29_port, A_signal(28) => 
                           positive_inputs_14_28_port, A_signal(27) => 
                           positive_inputs_14_27_port, A_signal(26) => 
                           positive_inputs_14_26_port, A_signal(25) => 
                           positive_inputs_14_25_port, A_signal(24) => 
                           positive_inputs_14_24_port, A_signal(23) => 
                           positive_inputs_14_23_port, A_signal(22) => 
                           positive_inputs_14_22_port, A_signal(21) => 
                           positive_inputs_14_21_port, A_signal(20) => 
                           positive_inputs_14_20_port, A_signal(19) => 
                           positive_inputs_14_19_port, A_signal(18) => 
                           positive_inputs_14_18_port, A_signal(17) => 
                           positive_inputs_14_17_port, A_signal(16) => 
                           positive_inputs_14_16_port, A_signal(15) => 
                           positive_inputs_14_15_port, A_signal(14) => 
                           positive_inputs_14_14_port, A_signal(13) => 
                           positive_inputs_14_13_port, A_signal(12) => 
                           positive_inputs_14_12_port, A_signal(11) => 
                           positive_inputs_14_11_port, A_signal(10) => 
                           positive_inputs_14_10_port, A_signal(9) => 
                           positive_inputs_14_9_port, A_signal(8) => 
                           positive_inputs_14_8_port, A_signal(7) => 
                           positive_inputs_14_7_port, A_signal(6) => 
                           positive_inputs_14_6_port, A_signal(5) => 
                           positive_inputs_14_5_port, A_signal(4) => 
                           positive_inputs_14_4_port, A_signal(3) => 
                           positive_inputs_14_3_port, A_signal(2) => 
                           positive_inputs_14_2_port, A_signal(1) => 
                           positive_inputs_14_1_port, A_signal(0) => n9, 
                           A_neg(63) => negative_inputs_14_63_port, A_neg(62) 
                           => negative_inputs_14_62_port, A_neg(61) => 
                           negative_inputs_14_61_port, A_neg(60) => 
                           negative_inputs_14_60_port, A_neg(59) => 
                           negative_inputs_14_59_port, A_neg(58) => 
                           negative_inputs_14_58_port, A_neg(57) => 
                           negative_inputs_14_57_port, A_neg(56) => 
                           negative_inputs_14_56_port, A_neg(55) => 
                           negative_inputs_14_55_port, A_neg(54) => 
                           negative_inputs_14_54_port, A_neg(53) => 
                           negative_inputs_14_53_port, A_neg(52) => 
                           negative_inputs_14_52_port, A_neg(51) => 
                           negative_inputs_14_51_port, A_neg(50) => 
                           negative_inputs_14_50_port, A_neg(49) => 
                           negative_inputs_14_49_port, A_neg(48) => n142, 
                           A_neg(47) => negative_inputs_14_47_port, A_neg(46) 
                           => negative_inputs_14_46_port, A_neg(45) => 
                           negative_inputs_14_45_port, A_neg(44) => 
                           negative_inputs_14_44_port, A_neg(43) => 
                           negative_inputs_14_43_port, A_neg(42) => 
                           negative_inputs_14_42_port, A_neg(41) => 
                           negative_inputs_14_41_port, A_neg(40) => 
                           negative_inputs_14_40_port, A_neg(39) => 
                           negative_inputs_14_39_port, A_neg(38) => 
                           negative_inputs_14_38_port, A_neg(37) => 
                           negative_inputs_14_37_port, A_neg(36) => 
                           negative_inputs_14_36_port, A_neg(35) => 
                           negative_inputs_14_35_port, A_neg(34) => 
                           negative_inputs_14_34_port, A_neg(33) => 
                           negative_inputs_14_33_port, A_neg(32) => 
                           negative_inputs_14_32_port, A_neg(31) => 
                           negative_inputs_14_31_port, A_neg(30) => 
                           negative_inputs_14_30_port, A_neg(29) => 
                           negative_inputs_14_29_port, A_neg(28) => 
                           negative_inputs_14_28_port, A_neg(27) => 
                           negative_inputs_14_27_port, A_neg(26) => 
                           negative_inputs_14_26_port, A_neg(25) => 
                           negative_inputs_14_25_port, A_neg(24) => 
                           negative_inputs_14_24_port, A_neg(23) => 
                           negative_inputs_14_23_port, A_neg(22) => 
                           negative_inputs_14_22_port, A_neg(21) => 
                           negative_inputs_14_21_port, A_neg(20) => 
                           negative_inputs_14_20_port, A_neg(19) => 
                           negative_inputs_14_19_port, A_neg(18) => 
                           negative_inputs_14_18_port, A_neg(17) => 
                           negative_inputs_14_17_port, A_neg(16) => 
                           negative_inputs_14_16_port, A_neg(15) => 
                           negative_inputs_14_15_port, A_neg(14) => 
                           negative_inputs_14_14_port, A_neg(13) => 
                           negative_inputs_14_13_port, A_neg(12) => 
                           negative_inputs_14_12_port, A_neg(11) => 
                           negative_inputs_14_11_port, A_neg(10) => 
                           negative_inputs_14_10_port, A_neg(9) => 
                           negative_inputs_14_9_port, A_neg(8) => 
                           negative_inputs_14_8_port, A_neg(7) => 
                           negative_inputs_14_7_port, A_neg(6) => 
                           negative_inputs_14_6_port, A_neg(5) => 
                           negative_inputs_14_5_port, A_neg(4) => 
                           negative_inputs_14_4_port, A_neg(3) => 
                           negative_inputs_14_3_port, A_neg(2) => 
                           negative_inputs_14_2_port, A_neg(1) => 
                           negative_inputs_14_1_port, A_neg(0) => n9, 
                           A_shifted(63) => positive_inputs_15_63_port, 
                           A_shifted(62) => positive_inputs_15_62_port, 
                           A_shifted(61) => positive_inputs_15_61_port, 
                           A_shifted(60) => positive_inputs_15_60_port, 
                           A_shifted(59) => positive_inputs_15_59_port, 
                           A_shifted(58) => positive_inputs_15_58_port, 
                           A_shifted(57) => positive_inputs_15_57_port, 
                           A_shifted(56) => positive_inputs_15_56_port, 
                           A_shifted(55) => positive_inputs_15_55_port, 
                           A_shifted(54) => positive_inputs_15_54_port, 
                           A_shifted(53) => positive_inputs_15_53_port, 
                           A_shifted(52) => positive_inputs_15_52_port, 
                           A_shifted(51) => positive_inputs_15_51_port, 
                           A_shifted(50) => positive_inputs_15_50_port, 
                           A_shifted(49) => positive_inputs_15_49_port, 
                           A_shifted(48) => n58, A_shifted(47) => 
                           positive_inputs_15_47_port, A_shifted(46) => 
                           positive_inputs_15_46_port, A_shifted(45) => 
                           positive_inputs_15_45_port, A_shifted(44) => 
                           positive_inputs_15_44_port, A_shifted(43) => 
                           positive_inputs_15_43_port, A_shifted(42) => 
                           positive_inputs_15_42_port, A_shifted(41) => 
                           positive_inputs_15_41_port, A_shifted(40) => 
                           positive_inputs_15_40_port, A_shifted(39) => 
                           positive_inputs_15_39_port, A_shifted(38) => 
                           positive_inputs_15_38_port, A_shifted(37) => 
                           positive_inputs_15_37_port, A_shifted(36) => 
                           positive_inputs_15_36_port, A_shifted(35) => 
                           positive_inputs_15_35_port, A_shifted(34) => 
                           positive_inputs_15_34_port, A_shifted(33) => 
                           positive_inputs_15_33_port, A_shifted(32) => 
                           positive_inputs_15_32_port, A_shifted(31) => 
                           positive_inputs_15_31_port, A_shifted(30) => 
                           positive_inputs_15_30_port, A_shifted(29) => 
                           positive_inputs_15_29_port, A_shifted(28) => 
                           positive_inputs_15_28_port, A_shifted(27) => 
                           positive_inputs_15_27_port, A_shifted(26) => 
                           positive_inputs_15_26_port, A_shifted(25) => 
                           positive_inputs_15_25_port, A_shifted(24) => 
                           positive_inputs_15_24_port, A_shifted(23) => 
                           positive_inputs_15_23_port, A_shifted(22) => 
                           positive_inputs_15_22_port, A_shifted(21) => 
                           positive_inputs_15_21_port, A_shifted(20) => 
                           positive_inputs_15_20_port, A_shifted(19) => 
                           positive_inputs_15_19_port, A_shifted(18) => 
                           positive_inputs_15_18_port, A_shifted(17) => 
                           positive_inputs_15_17_port, A_shifted(16) => 
                           positive_inputs_15_16_port, A_shifted(15) => 
                           positive_inputs_15_15_port, A_shifted(14) => 
                           positive_inputs_15_14_port, A_shifted(13) => 
                           positive_inputs_15_13_port, A_shifted(12) => 
                           positive_inputs_15_12_port, A_shifted(11) => 
                           positive_inputs_15_11_port, A_shifted(10) => 
                           positive_inputs_15_10_port, A_shifted(9) => 
                           positive_inputs_15_9_port, A_shifted(8) => 
                           positive_inputs_15_8_port, A_shifted(7) => 
                           positive_inputs_15_7_port, A_shifted(6) => 
                           positive_inputs_15_6_port, A_shifted(5) => 
                           positive_inputs_15_5_port, A_shifted(4) => 
                           positive_inputs_15_4_port, A_shifted(3) => 
                           positive_inputs_15_3_port, A_shifted(2) => 
                           positive_inputs_15_2_port, A_shifted(1) => 
                           positive_inputs_15_1_port, A_shifted(0) => n9, 
                           A_neg_shifted(63) => negative_inputs_15_63_port, 
                           A_neg_shifted(62) => negative_inputs_15_62_port, 
                           A_neg_shifted(61) => negative_inputs_15_61_port, 
                           A_neg_shifted(60) => negative_inputs_15_60_port, 
                           A_neg_shifted(59) => negative_inputs_15_59_port, 
                           A_neg_shifted(58) => negative_inputs_15_58_port, 
                           A_neg_shifted(57) => negative_inputs_15_57_port, 
                           A_neg_shifted(56) => negative_inputs_15_56_port, 
                           A_neg_shifted(55) => negative_inputs_15_55_port, 
                           A_neg_shifted(54) => negative_inputs_15_54_port, 
                           A_neg_shifted(53) => negative_inputs_15_53_port, 
                           A_neg_shifted(52) => negative_inputs_15_52_port, 
                           A_neg_shifted(51) => negative_inputs_15_51_port, 
                           A_neg_shifted(50) => negative_inputs_15_50_port, 
                           A_neg_shifted(49) => negative_inputs_15_49_port, 
                           A_neg_shifted(48) => n140, A_neg_shifted(47) => 
                           negative_inputs_15_47_port, A_neg_shifted(46) => 
                           negative_inputs_15_46_port, A_neg_shifted(45) => 
                           negative_inputs_15_45_port, A_neg_shifted(44) => 
                           negative_inputs_15_44_port, A_neg_shifted(43) => 
                           negative_inputs_15_43_port, A_neg_shifted(42) => 
                           negative_inputs_15_42_port, A_neg_shifted(41) => 
                           negative_inputs_15_41_port, A_neg_shifted(40) => 
                           negative_inputs_15_40_port, A_neg_shifted(39) => 
                           negative_inputs_15_39_port, A_neg_shifted(38) => 
                           negative_inputs_15_38_port, A_neg_shifted(37) => 
                           negative_inputs_15_37_port, A_neg_shifted(36) => 
                           negative_inputs_15_36_port, A_neg_shifted(35) => 
                           negative_inputs_15_35_port, A_neg_shifted(34) => 
                           negative_inputs_15_34_port, A_neg_shifted(33) => 
                           negative_inputs_15_33_port, A_neg_shifted(32) => 
                           negative_inputs_15_32_port, A_neg_shifted(31) => 
                           negative_inputs_15_31_port, A_neg_shifted(30) => 
                           negative_inputs_15_30_port, A_neg_shifted(29) => 
                           negative_inputs_15_29_port, A_neg_shifted(28) => 
                           negative_inputs_15_28_port, A_neg_shifted(27) => 
                           negative_inputs_15_27_port, A_neg_shifted(26) => 
                           negative_inputs_15_26_port, A_neg_shifted(25) => 
                           negative_inputs_15_25_port, A_neg_shifted(24) => 
                           negative_inputs_15_24_port, A_neg_shifted(23) => 
                           negative_inputs_15_23_port, A_neg_shifted(22) => 
                           negative_inputs_15_22_port, A_neg_shifted(21) => 
                           negative_inputs_15_21_port, A_neg_shifted(20) => 
                           negative_inputs_15_20_port, A_neg_shifted(19) => 
                           negative_inputs_15_19_port, A_neg_shifted(18) => 
                           negative_inputs_15_18_port, A_neg_shifted(17) => 
                           negative_inputs_15_17_port, A_neg_shifted(16) => 
                           negative_inputs_15_16_port, A_neg_shifted(15) => 
                           negative_inputs_15_15_port, A_neg_shifted(14) => 
                           negative_inputs_15_14_port, A_neg_shifted(13) => 
                           negative_inputs_15_13_port, A_neg_shifted(12) => 
                           negative_inputs_15_12_port, A_neg_shifted(11) => 
                           negative_inputs_15_11_port, A_neg_shifted(10) => 
                           negative_inputs_15_10_port, A_neg_shifted(9) => 
                           negative_inputs_15_9_port, A_neg_shifted(8) => 
                           negative_inputs_15_8_port, A_neg_shifted(7) => 
                           negative_inputs_15_7_port, A_neg_shifted(6) => 
                           negative_inputs_15_6_port, A_neg_shifted(5) => 
                           negative_inputs_15_5_port, A_neg_shifted(4) => 
                           negative_inputs_15_4_port, A_neg_shifted(3) => 
                           negative_inputs_15_3_port, A_neg_shifted(2) => 
                           negative_inputs_15_2_port, A_neg_shifted(1) => 
                           negative_inputs_15_1_port, A_neg_shifted(0) => n9, 
                           Sel(2) => sel_7_2_port, Sel(1) => sel_7_1_port, 
                           Sel(0) => sel_7_0_port, Y(63) => 
                           MuxOutputs_7_63_port, Y(62) => MuxOutputs_7_62_port,
                           Y(61) => MuxOutputs_7_61_port, Y(60) => 
                           MuxOutputs_7_60_port, Y(59) => MuxOutputs_7_59_port,
                           Y(58) => MuxOutputs_7_58_port, Y(57) => 
                           MuxOutputs_7_57_port, Y(56) => MuxOutputs_7_56_port,
                           Y(55) => MuxOutputs_7_55_port, Y(54) => 
                           MuxOutputs_7_54_port, Y(53) => MuxOutputs_7_53_port,
                           Y(52) => MuxOutputs_7_52_port, Y(51) => 
                           MuxOutputs_7_51_port, Y(50) => MuxOutputs_7_50_port,
                           Y(49) => MuxOutputs_7_49_port, Y(48) => 
                           MuxOutputs_7_48_port, Y(47) => MuxOutputs_7_47_port,
                           Y(46) => MuxOutputs_7_46_port, Y(45) => 
                           MuxOutputs_7_45_port, Y(44) => MuxOutputs_7_44_port,
                           Y(43) => MuxOutputs_7_43_port, Y(42) => 
                           MuxOutputs_7_42_port, Y(41) => MuxOutputs_7_41_port,
                           Y(40) => MuxOutputs_7_40_port, Y(39) => 
                           MuxOutputs_7_39_port, Y(38) => MuxOutputs_7_38_port,
                           Y(37) => MuxOutputs_7_37_port, Y(36) => 
                           MuxOutputs_7_36_port, Y(35) => MuxOutputs_7_35_port,
                           Y(34) => MuxOutputs_7_34_port, Y(33) => 
                           MuxOutputs_7_33_port, Y(32) => MuxOutputs_7_32_port,
                           Y(31) => MuxOutputs_7_31_port, Y(30) => 
                           MuxOutputs_7_30_port, Y(29) => MuxOutputs_7_29_port,
                           Y(28) => MuxOutputs_7_28_port, Y(27) => 
                           MuxOutputs_7_27_port, Y(26) => MuxOutputs_7_26_port,
                           Y(25) => MuxOutputs_7_25_port, Y(24) => 
                           MuxOutputs_7_24_port, Y(23) => MuxOutputs_7_23_port,
                           Y(22) => MuxOutputs_7_22_port, Y(21) => 
                           MuxOutputs_7_21_port, Y(20) => MuxOutputs_7_20_port,
                           Y(19) => MuxOutputs_7_19_port, Y(18) => 
                           MuxOutputs_7_18_port, Y(17) => MuxOutputs_7_17_port,
                           Y(16) => MuxOutputs_7_16_port, Y(15) => 
                           MuxOutputs_7_15_port, Y(14) => MuxOutputs_7_14_port,
                           Y(13) => MuxOutputs_7_13_port, Y(12) => 
                           MuxOutputs_7_12_port, Y(11) => MuxOutputs_7_11_port,
                           Y(10) => MuxOutputs_7_10_port, Y(9) => 
                           MuxOutputs_7_9_port, Y(8) => MuxOutputs_7_8_port, 
                           Y(7) => MuxOutputs_7_7_port, Y(6) => 
                           MuxOutputs_7_6_port, Y(5) => MuxOutputs_7_5_port, 
                           Y(4) => MuxOutputs_7_4_port, Y(3) => 
                           MuxOutputs_7_3_port, Y(2) => MuxOutputs_7_2_port, 
                           Y(1) => MuxOutputs_7_1_port, Y(0) => 
                           MuxOutputs_7_0_port);
   encoderI_8 : encoder_8 port map( pieceofB(2) => B(17), pieceofB(1) => B(16),
                           pieceofB(0) => B(15), sel(2) => sel_8_2_port, sel(1)
                           => sel_8_1_port, sel(0) => sel_8_0_port);
   MUXI_8 : MUX51_MuxNbit64_8 port map( zeroSignal(63) => X_Logic0_port, 
                           zeroSignal(62) => X_Logic0_port, zeroSignal(61) => 
                           X_Logic0_port, zeroSignal(60) => X_Logic0_port, 
                           zeroSignal(59) => X_Logic0_port, zeroSignal(58) => 
                           X_Logic0_port, zeroSignal(57) => X_Logic0_port, 
                           zeroSignal(56) => X_Logic0_port, zeroSignal(55) => 
                           X_Logic0_port, zeroSignal(54) => X_Logic0_port, 
                           zeroSignal(53) => X_Logic0_port, zeroSignal(52) => 
                           X_Logic0_port, zeroSignal(51) => X_Logic0_port, 
                           zeroSignal(50) => X_Logic0_port, zeroSignal(49) => 
                           X_Logic0_port, zeroSignal(48) => X_Logic0_port, 
                           zeroSignal(47) => X_Logic0_port, zeroSignal(46) => 
                           X_Logic0_port, zeroSignal(45) => X_Logic0_port, 
                           zeroSignal(44) => X_Logic0_port, zeroSignal(43) => 
                           X_Logic0_port, zeroSignal(42) => X_Logic0_port, 
                           zeroSignal(41) => X_Logic0_port, zeroSignal(40) => 
                           X_Logic0_port, zeroSignal(39) => X_Logic0_port, 
                           zeroSignal(38) => X_Logic0_port, zeroSignal(37) => 
                           X_Logic0_port, zeroSignal(36) => X_Logic0_port, 
                           zeroSignal(35) => X_Logic0_port, zeroSignal(34) => 
                           X_Logic0_port, zeroSignal(33) => X_Logic0_port, 
                           zeroSignal(32) => X_Logic0_port, zeroSignal(31) => 
                           X_Logic0_port, zeroSignal(30) => X_Logic0_port, 
                           zeroSignal(29) => X_Logic0_port, zeroSignal(28) => 
                           X_Logic0_port, zeroSignal(27) => X_Logic0_port, 
                           zeroSignal(26) => X_Logic0_port, zeroSignal(25) => 
                           X_Logic0_port, zeroSignal(24) => X_Logic0_port, 
                           zeroSignal(23) => X_Logic0_port, zeroSignal(22) => 
                           X_Logic0_port, zeroSignal(21) => X_Logic0_port, 
                           zeroSignal(20) => X_Logic0_port, zeroSignal(19) => 
                           X_Logic0_port, zeroSignal(18) => X_Logic0_port, 
                           zeroSignal(17) => X_Logic0_port, zeroSignal(16) => 
                           X_Logic0_port, zeroSignal(15) => X_Logic0_port, 
                           zeroSignal(14) => X_Logic0_port, zeroSignal(13) => 
                           X_Logic0_port, zeroSignal(12) => X_Logic0_port, 
                           zeroSignal(11) => X_Logic0_port, zeroSignal(10) => 
                           X_Logic0_port, zeroSignal(9) => X_Logic0_port, 
                           zeroSignal(8) => X_Logic0_port, zeroSignal(7) => 
                           X_Logic0_port, zeroSignal(6) => X_Logic0_port, 
                           zeroSignal(5) => X_Logic0_port, zeroSignal(4) => 
                           X_Logic0_port, zeroSignal(3) => X_Logic0_port, 
                           zeroSignal(2) => X_Logic0_port, zeroSignal(1) => 
                           X_Logic0_port, zeroSignal(0) => X_Logic0_port, 
                           A_signal(63) => positive_inputs_16_63_port, 
                           A_signal(62) => positive_inputs_16_62_port, 
                           A_signal(61) => positive_inputs_16_61_port, 
                           A_signal(60) => positive_inputs_16_60_port, 
                           A_signal(59) => positive_inputs_16_59_port, 
                           A_signal(58) => positive_inputs_16_58_port, 
                           A_signal(57) => positive_inputs_16_57_port, 
                           A_signal(56) => positive_inputs_16_56_port, 
                           A_signal(55) => positive_inputs_16_55_port, 
                           A_signal(54) => positive_inputs_16_54_port, 
                           A_signal(53) => positive_inputs_16_53_port, 
                           A_signal(52) => positive_inputs_16_52_port, 
                           A_signal(51) => positive_inputs_16_51_port, 
                           A_signal(50) => positive_inputs_16_50_port, 
                           A_signal(49) => positive_inputs_16_49_port, 
                           A_signal(48) => n57, A_signal(47) => n56, 
                           A_signal(46) => n215, A_signal(45) => n213, 
                           A_signal(44) => n211, A_signal(43) => n209, 
                           A_signal(42) => n207, A_signal(41) => n205, 
                           A_signal(40) => n203, A_signal(39) => n201, 
                           A_signal(38) => n199, A_signal(37) => n197, 
                           A_signal(36) => n195, A_signal(35) => n193, 
                           A_signal(34) => n191, A_signal(33) => n189, 
                           A_signal(32) => n187, A_signal(31) => n185, 
                           A_signal(30) => n183, A_signal(29) => n181, 
                           A_signal(28) => n179, A_signal(27) => n177, 
                           A_signal(26) => n175, A_signal(25) => n173, 
                           A_signal(24) => n171, A_signal(23) => n169, 
                           A_signal(22) => n167, A_signal(21) => n165, 
                           A_signal(20) => n163, A_signal(19) => n161, 
                           A_signal(18) => n159, A_signal(17) => n157, 
                           A_signal(16) => n155, A_signal(15) => 
                           positive_inputs_16_15_port, A_signal(14) => 
                           positive_inputs_16_14_port, A_signal(13) => 
                           positive_inputs_16_13_port, A_signal(12) => 
                           positive_inputs_16_12_port, A_signal(11) => 
                           positive_inputs_16_11_port, A_signal(10) => 
                           positive_inputs_16_10_port, A_signal(9) => 
                           positive_inputs_16_9_port, A_signal(8) => 
                           positive_inputs_16_8_port, A_signal(7) => 
                           positive_inputs_16_7_port, A_signal(6) => 
                           positive_inputs_16_6_port, A_signal(5) => 
                           positive_inputs_16_5_port, A_signal(4) => 
                           positive_inputs_16_4_port, A_signal(3) => 
                           positive_inputs_16_3_port, A_signal(2) => 
                           positive_inputs_16_2_port, A_signal(1) => 
                           positive_inputs_16_1_port, A_signal(0) => n9, 
                           A_neg(63) => negative_inputs_16_63_port, A_neg(62) 
                           => negative_inputs_16_62_port, A_neg(61) => 
                           negative_inputs_16_61_port, A_neg(60) => 
                           negative_inputs_16_60_port, A_neg(59) => 
                           negative_inputs_16_59_port, A_neg(58) => 
                           negative_inputs_16_58_port, A_neg(57) => 
                           negative_inputs_16_57_port, A_neg(56) => 
                           negative_inputs_16_56_port, A_neg(55) => 
                           negative_inputs_16_55_port, A_neg(54) => 
                           negative_inputs_16_54_port, A_neg(53) => 
                           negative_inputs_16_53_port, A_neg(52) => 
                           negative_inputs_16_52_port, A_neg(51) => 
                           negative_inputs_16_51_port, A_neg(50) => 
                           negative_inputs_16_50_port, A_neg(49) => 
                           negative_inputs_16_49_port, A_neg(48) => n138, 
                           A_neg(47) => n136, A_neg(46) => n134, A_neg(45) => 
                           n132, A_neg(44) => n130, A_neg(43) => n128, 
                           A_neg(42) => n126, A_neg(41) => n124, A_neg(40) => 
                           n122, A_neg(39) => n120, A_neg(38) => n118, 
                           A_neg(37) => n116, A_neg(36) => n114, A_neg(35) => 
                           n112, A_neg(34) => n110, A_neg(33) => n108, 
                           A_neg(32) => n106, A_neg(31) => n104, A_neg(30) => 
                           n102, A_neg(29) => n100, A_neg(28) => n98, A_neg(27)
                           => n96, A_neg(26) => n94, A_neg(25) => n92, 
                           A_neg(24) => n90, A_neg(23) => n88, A_neg(22) => n86
                           , A_neg(21) => n84, A_neg(20) => n82, A_neg(19) => 
                           n80, A_neg(18) => n78, A_neg(17) => n76, A_neg(16) 
                           => n74, A_neg(15) => negative_inputs_16_15_port, 
                           A_neg(14) => negative_inputs_16_14_port, A_neg(13) 
                           => negative_inputs_16_13_port, A_neg(12) => 
                           negative_inputs_16_12_port, A_neg(11) => 
                           negative_inputs_16_11_port, A_neg(10) => 
                           negative_inputs_16_10_port, A_neg(9) => 
                           negative_inputs_16_9_port, A_neg(8) => 
                           negative_inputs_16_8_port, A_neg(7) => 
                           negative_inputs_16_7_port, A_neg(6) => 
                           negative_inputs_16_6_port, A_neg(5) => 
                           negative_inputs_16_5_port, A_neg(4) => 
                           negative_inputs_16_4_port, A_neg(3) => 
                           negative_inputs_16_3_port, A_neg(2) => 
                           negative_inputs_16_2_port, A_neg(1) => 
                           negative_inputs_16_1_port, A_neg(0) => n9, 
                           A_shifted(63) => positive_inputs_17_63_port, 
                           A_shifted(62) => positive_inputs_17_62_port, 
                           A_shifted(61) => positive_inputs_17_61_port, 
                           A_shifted(60) => positive_inputs_17_60_port, 
                           A_shifted(59) => positive_inputs_17_59_port, 
                           A_shifted(58) => positive_inputs_17_58_port, 
                           A_shifted(57) => positive_inputs_17_57_port, 
                           A_shifted(56) => positive_inputs_17_56_port, 
                           A_shifted(55) => positive_inputs_17_55_port, 
                           A_shifted(54) => positive_inputs_17_54_port, 
                           A_shifted(53) => positive_inputs_17_53_port, 
                           A_shifted(52) => positive_inputs_17_52_port, 
                           A_shifted(51) => positive_inputs_17_51_port, 
                           A_shifted(50) => positive_inputs_17_50_port, 
                           A_shifted(49) => positive_inputs_17_49_port, 
                           A_shifted(48) => positive_inputs_17_48_port, 
                           A_shifted(47) => positive_inputs_17_47_port, 
                           A_shifted(46) => positive_inputs_17_46_port, 
                           A_shifted(45) => positive_inputs_17_45_port, 
                           A_shifted(44) => positive_inputs_17_44_port, 
                           A_shifted(43) => positive_inputs_17_43_port, 
                           A_shifted(42) => positive_inputs_17_42_port, 
                           A_shifted(41) => positive_inputs_17_41_port, 
                           A_shifted(40) => positive_inputs_17_40_port, 
                           A_shifted(39) => positive_inputs_17_39_port, 
                           A_shifted(38) => positive_inputs_17_38_port, 
                           A_shifted(37) => positive_inputs_17_37_port, 
                           A_shifted(36) => positive_inputs_17_36_port, 
                           A_shifted(35) => positive_inputs_17_35_port, 
                           A_shifted(34) => positive_inputs_17_34_port, 
                           A_shifted(33) => positive_inputs_17_33_port, 
                           A_shifted(32) => positive_inputs_17_32_port, 
                           A_shifted(31) => positive_inputs_17_31_port, 
                           A_shifted(30) => positive_inputs_17_30_port, 
                           A_shifted(29) => positive_inputs_17_29_port, 
                           A_shifted(28) => positive_inputs_17_28_port, 
                           A_shifted(27) => positive_inputs_17_27_port, 
                           A_shifted(26) => positive_inputs_17_26_port, 
                           A_shifted(25) => positive_inputs_17_25_port, 
                           A_shifted(24) => positive_inputs_17_24_port, 
                           A_shifted(23) => positive_inputs_17_23_port, 
                           A_shifted(22) => positive_inputs_17_22_port, 
                           A_shifted(21) => positive_inputs_17_21_port, 
                           A_shifted(20) => positive_inputs_17_20_port, 
                           A_shifted(19) => positive_inputs_17_19_port, 
                           A_shifted(18) => positive_inputs_17_18_port, 
                           A_shifted(17) => positive_inputs_17_17_port, 
                           A_shifted(16) => positive_inputs_17_16_port, 
                           A_shifted(15) => positive_inputs_17_15_port, 
                           A_shifted(14) => positive_inputs_17_14_port, 
                           A_shifted(13) => positive_inputs_17_13_port, 
                           A_shifted(12) => positive_inputs_17_12_port, 
                           A_shifted(11) => positive_inputs_17_11_port, 
                           A_shifted(10) => positive_inputs_17_10_port, 
                           A_shifted(9) => positive_inputs_17_9_port, 
                           A_shifted(8) => positive_inputs_17_8_port, 
                           A_shifted(7) => positive_inputs_17_7_port, 
                           A_shifted(6) => positive_inputs_17_6_port, 
                           A_shifted(5) => positive_inputs_17_5_port, 
                           A_shifted(4) => positive_inputs_17_4_port, 
                           A_shifted(3) => positive_inputs_17_3_port, 
                           A_shifted(2) => positive_inputs_17_2_port, 
                           A_shifted(1) => positive_inputs_17_1_port, 
                           A_shifted(0) => n9, A_neg_shifted(63) => 
                           negative_inputs_17_63_port, A_neg_shifted(62) => 
                           negative_inputs_17_62_port, A_neg_shifted(61) => 
                           negative_inputs_17_61_port, A_neg_shifted(60) => 
                           negative_inputs_17_60_port, A_neg_shifted(59) => 
                           negative_inputs_17_59_port, A_neg_shifted(58) => 
                           negative_inputs_17_58_port, A_neg_shifted(57) => 
                           negative_inputs_17_57_port, A_neg_shifted(56) => 
                           negative_inputs_17_56_port, A_neg_shifted(55) => 
                           negative_inputs_17_55_port, A_neg_shifted(54) => 
                           negative_inputs_17_54_port, A_neg_shifted(53) => 
                           negative_inputs_17_53_port, A_neg_shifted(52) => 
                           negative_inputs_17_52_port, A_neg_shifted(51) => 
                           negative_inputs_17_51_port, A_neg_shifted(50) => 
                           negative_inputs_17_50_port, A_neg_shifted(49) => 
                           negative_inputs_17_49_port, A_neg_shifted(48) => 
                           negative_inputs_17_48_port, A_neg_shifted(47) => 
                           negative_inputs_17_47_port, A_neg_shifted(46) => 
                           negative_inputs_17_46_port, A_neg_shifted(45) => 
                           negative_inputs_17_45_port, A_neg_shifted(44) => 
                           negative_inputs_17_44_port, A_neg_shifted(43) => 
                           negative_inputs_17_43_port, A_neg_shifted(42) => 
                           negative_inputs_17_42_port, A_neg_shifted(41) => 
                           negative_inputs_17_41_port, A_neg_shifted(40) => 
                           negative_inputs_17_40_port, A_neg_shifted(39) => 
                           negative_inputs_17_39_port, A_neg_shifted(38) => 
                           negative_inputs_17_38_port, A_neg_shifted(37) => 
                           negative_inputs_17_37_port, A_neg_shifted(36) => 
                           negative_inputs_17_36_port, A_neg_shifted(35) => 
                           negative_inputs_17_35_port, A_neg_shifted(34) => 
                           negative_inputs_17_34_port, A_neg_shifted(33) => 
                           negative_inputs_17_33_port, A_neg_shifted(32) => 
                           negative_inputs_17_32_port, A_neg_shifted(31) => 
                           negative_inputs_17_31_port, A_neg_shifted(30) => 
                           negative_inputs_17_30_port, A_neg_shifted(29) => 
                           negative_inputs_17_29_port, A_neg_shifted(28) => 
                           negative_inputs_17_28_port, A_neg_shifted(27) => 
                           negative_inputs_17_27_port, A_neg_shifted(26) => 
                           negative_inputs_17_26_port, A_neg_shifted(25) => 
                           negative_inputs_17_25_port, A_neg_shifted(24) => 
                           negative_inputs_17_24_port, A_neg_shifted(23) => 
                           negative_inputs_17_23_port, A_neg_shifted(22) => 
                           negative_inputs_17_22_port, A_neg_shifted(21) => 
                           negative_inputs_17_21_port, A_neg_shifted(20) => 
                           negative_inputs_17_20_port, A_neg_shifted(19) => 
                           negative_inputs_17_19_port, A_neg_shifted(18) => 
                           negative_inputs_17_18_port, A_neg_shifted(17) => 
                           negative_inputs_17_17_port, A_neg_shifted(16) => 
                           negative_inputs_17_16_port, A_neg_shifted(15) => 
                           negative_inputs_17_15_port, A_neg_shifted(14) => 
                           negative_inputs_17_14_port, A_neg_shifted(13) => 
                           negative_inputs_17_13_port, A_neg_shifted(12) => 
                           negative_inputs_17_12_port, A_neg_shifted(11) => 
                           negative_inputs_17_11_port, A_neg_shifted(10) => 
                           negative_inputs_17_10_port, A_neg_shifted(9) => 
                           negative_inputs_17_9_port, A_neg_shifted(8) => 
                           negative_inputs_17_8_port, A_neg_shifted(7) => 
                           negative_inputs_17_7_port, A_neg_shifted(6) => 
                           negative_inputs_17_6_port, A_neg_shifted(5) => 
                           negative_inputs_17_5_port, A_neg_shifted(4) => 
                           negative_inputs_17_4_port, A_neg_shifted(3) => 
                           negative_inputs_17_3_port, A_neg_shifted(2) => 
                           negative_inputs_17_2_port, A_neg_shifted(1) => 
                           negative_inputs_17_1_port, A_neg_shifted(0) => n9, 
                           Sel(2) => sel_8_2_port, Sel(1) => sel_8_1_port, 
                           Sel(0) => sel_8_0_port, Y(63) => 
                           MuxOutputs_8_63_port, Y(62) => MuxOutputs_8_62_port,
                           Y(61) => MuxOutputs_8_61_port, Y(60) => 
                           MuxOutputs_8_60_port, Y(59) => MuxOutputs_8_59_port,
                           Y(58) => MuxOutputs_8_58_port, Y(57) => 
                           MuxOutputs_8_57_port, Y(56) => MuxOutputs_8_56_port,
                           Y(55) => MuxOutputs_8_55_port, Y(54) => 
                           MuxOutputs_8_54_port, Y(53) => MuxOutputs_8_53_port,
                           Y(52) => MuxOutputs_8_52_port, Y(51) => 
                           MuxOutputs_8_51_port, Y(50) => MuxOutputs_8_50_port,
                           Y(49) => MuxOutputs_8_49_port, Y(48) => 
                           MuxOutputs_8_48_port, Y(47) => MuxOutputs_8_47_port,
                           Y(46) => MuxOutputs_8_46_port, Y(45) => 
                           MuxOutputs_8_45_port, Y(44) => MuxOutputs_8_44_port,
                           Y(43) => MuxOutputs_8_43_port, Y(42) => 
                           MuxOutputs_8_42_port, Y(41) => MuxOutputs_8_41_port,
                           Y(40) => MuxOutputs_8_40_port, Y(39) => 
                           MuxOutputs_8_39_port, Y(38) => MuxOutputs_8_38_port,
                           Y(37) => MuxOutputs_8_37_port, Y(36) => 
                           MuxOutputs_8_36_port, Y(35) => MuxOutputs_8_35_port,
                           Y(34) => MuxOutputs_8_34_port, Y(33) => 
                           MuxOutputs_8_33_port, Y(32) => MuxOutputs_8_32_port,
                           Y(31) => MuxOutputs_8_31_port, Y(30) => 
                           MuxOutputs_8_30_port, Y(29) => MuxOutputs_8_29_port,
                           Y(28) => MuxOutputs_8_28_port, Y(27) => 
                           MuxOutputs_8_27_port, Y(26) => MuxOutputs_8_26_port,
                           Y(25) => MuxOutputs_8_25_port, Y(24) => 
                           MuxOutputs_8_24_port, Y(23) => MuxOutputs_8_23_port,
                           Y(22) => MuxOutputs_8_22_port, Y(21) => 
                           MuxOutputs_8_21_port, Y(20) => MuxOutputs_8_20_port,
                           Y(19) => MuxOutputs_8_19_port, Y(18) => 
                           MuxOutputs_8_18_port, Y(17) => MuxOutputs_8_17_port,
                           Y(16) => MuxOutputs_8_16_port, Y(15) => 
                           MuxOutputs_8_15_port, Y(14) => MuxOutputs_8_14_port,
                           Y(13) => MuxOutputs_8_13_port, Y(12) => 
                           MuxOutputs_8_12_port, Y(11) => MuxOutputs_8_11_port,
                           Y(10) => MuxOutputs_8_10_port, Y(9) => 
                           MuxOutputs_8_9_port, Y(8) => MuxOutputs_8_8_port, 
                           Y(7) => MuxOutputs_8_7_port, Y(6) => 
                           MuxOutputs_8_6_port, Y(5) => MuxOutputs_8_5_port, 
                           Y(4) => MuxOutputs_8_4_port, Y(3) => 
                           MuxOutputs_8_3_port, Y(2) => MuxOutputs_8_2_port, 
                           Y(1) => MuxOutputs_8_1_port, Y(0) => 
                           MuxOutputs_8_0_port);
   encoderI_9 : encoder_7 port map( pieceofB(2) => B(19), pieceofB(1) => B(18),
                           pieceofB(0) => B(17), sel(2) => sel_9_2_port, sel(1)
                           => sel_9_1_port, sel(0) => sel_9_0_port);
   MUXI_9 : MUX51_MuxNbit64_7 port map( zeroSignal(63) => X_Logic0_port, 
                           zeroSignal(62) => X_Logic0_port, zeroSignal(61) => 
                           X_Logic0_port, zeroSignal(60) => X_Logic0_port, 
                           zeroSignal(59) => X_Logic0_port, zeroSignal(58) => 
                           X_Logic0_port, zeroSignal(57) => X_Logic0_port, 
                           zeroSignal(56) => X_Logic0_port, zeroSignal(55) => 
                           X_Logic0_port, zeroSignal(54) => X_Logic0_port, 
                           zeroSignal(53) => X_Logic0_port, zeroSignal(52) => 
                           X_Logic0_port, zeroSignal(51) => X_Logic0_port, 
                           zeroSignal(50) => X_Logic0_port, zeroSignal(49) => 
                           X_Logic0_port, zeroSignal(48) => X_Logic0_port, 
                           zeroSignal(47) => X_Logic0_port, zeroSignal(46) => 
                           X_Logic0_port, zeroSignal(45) => X_Logic0_port, 
                           zeroSignal(44) => X_Logic0_port, zeroSignal(43) => 
                           X_Logic0_port, zeroSignal(42) => X_Logic0_port, 
                           zeroSignal(41) => X_Logic0_port, zeroSignal(40) => 
                           X_Logic0_port, zeroSignal(39) => X_Logic0_port, 
                           zeroSignal(38) => X_Logic0_port, zeroSignal(37) => 
                           X_Logic0_port, zeroSignal(36) => X_Logic0_port, 
                           zeroSignal(35) => X_Logic0_port, zeroSignal(34) => 
                           X_Logic0_port, zeroSignal(33) => X_Logic0_port, 
                           zeroSignal(32) => X_Logic0_port, zeroSignal(31) => 
                           X_Logic0_port, zeroSignal(30) => X_Logic0_port, 
                           zeroSignal(29) => X_Logic0_port, zeroSignal(28) => 
                           X_Logic0_port, zeroSignal(27) => X_Logic0_port, 
                           zeroSignal(26) => X_Logic0_port, zeroSignal(25) => 
                           X_Logic0_port, zeroSignal(24) => X_Logic0_port, 
                           zeroSignal(23) => X_Logic0_port, zeroSignal(22) => 
                           X_Logic0_port, zeroSignal(21) => X_Logic0_port, 
                           zeroSignal(20) => X_Logic0_port, zeroSignal(19) => 
                           X_Logic0_port, zeroSignal(18) => X_Logic0_port, 
                           zeroSignal(17) => X_Logic0_port, zeroSignal(16) => 
                           X_Logic0_port, zeroSignal(15) => X_Logic0_port, 
                           zeroSignal(14) => X_Logic0_port, zeroSignal(13) => 
                           X_Logic0_port, zeroSignal(12) => X_Logic0_port, 
                           zeroSignal(11) => X_Logic0_port, zeroSignal(10) => 
                           X_Logic0_port, zeroSignal(9) => X_Logic0_port, 
                           zeroSignal(8) => X_Logic0_port, zeroSignal(7) => 
                           X_Logic0_port, zeroSignal(6) => X_Logic0_port, 
                           zeroSignal(5) => X_Logic0_port, zeroSignal(4) => 
                           X_Logic0_port, zeroSignal(3) => X_Logic0_port, 
                           zeroSignal(2) => X_Logic0_port, zeroSignal(1) => 
                           X_Logic0_port, zeroSignal(0) => X_Logic0_port, 
                           A_signal(63) => positive_inputs_18_63_port, 
                           A_signal(62) => positive_inputs_18_62_port, 
                           A_signal(61) => positive_inputs_18_61_port, 
                           A_signal(60) => positive_inputs_18_60_port, 
                           A_signal(59) => positive_inputs_18_59_port, 
                           A_signal(58) => positive_inputs_18_58_port, 
                           A_signal(57) => positive_inputs_18_57_port, 
                           A_signal(56) => positive_inputs_18_56_port, 
                           A_signal(55) => positive_inputs_18_55_port, 
                           A_signal(54) => positive_inputs_18_54_port, 
                           A_signal(53) => positive_inputs_18_53_port, 
                           A_signal(52) => positive_inputs_18_52_port, 
                           A_signal(51) => positive_inputs_18_51_port, 
                           A_signal(50) => positive_inputs_18_50_port, 
                           A_signal(49) => positive_inputs_18_49_port, 
                           A_signal(48) => positive_inputs_18_48_port, 
                           A_signal(47) => positive_inputs_18_47_port, 
                           A_signal(46) => positive_inputs_18_46_port, 
                           A_signal(45) => positive_inputs_18_45_port, 
                           A_signal(44) => positive_inputs_18_44_port, 
                           A_signal(43) => positive_inputs_18_43_port, 
                           A_signal(42) => positive_inputs_18_42_port, 
                           A_signal(41) => positive_inputs_18_41_port, 
                           A_signal(40) => positive_inputs_18_40_port, 
                           A_signal(39) => positive_inputs_18_39_port, 
                           A_signal(38) => positive_inputs_18_38_port, 
                           A_signal(37) => positive_inputs_18_37_port, 
                           A_signal(36) => positive_inputs_18_36_port, 
                           A_signal(35) => positive_inputs_18_35_port, 
                           A_signal(34) => positive_inputs_18_34_port, 
                           A_signal(33) => positive_inputs_18_33_port, 
                           A_signal(32) => positive_inputs_18_32_port, 
                           A_signal(31) => positive_inputs_18_31_port, 
                           A_signal(30) => positive_inputs_18_30_port, 
                           A_signal(29) => positive_inputs_18_29_port, 
                           A_signal(28) => positive_inputs_18_28_port, 
                           A_signal(27) => positive_inputs_18_27_port, 
                           A_signal(26) => positive_inputs_18_26_port, 
                           A_signal(25) => positive_inputs_18_25_port, 
                           A_signal(24) => positive_inputs_18_24_port, 
                           A_signal(23) => positive_inputs_18_23_port, 
                           A_signal(22) => positive_inputs_18_22_port, 
                           A_signal(21) => positive_inputs_18_21_port, 
                           A_signal(20) => positive_inputs_18_20_port, 
                           A_signal(19) => positive_inputs_18_19_port, 
                           A_signal(18) => positive_inputs_18_18_port, 
                           A_signal(17) => positive_inputs_18_17_port, 
                           A_signal(16) => positive_inputs_18_16_port, 
                           A_signal(15) => positive_inputs_18_15_port, 
                           A_signal(14) => positive_inputs_18_14_port, 
                           A_signal(13) => positive_inputs_18_13_port, 
                           A_signal(12) => positive_inputs_18_12_port, 
                           A_signal(11) => positive_inputs_18_11_port, 
                           A_signal(10) => positive_inputs_18_10_port, 
                           A_signal(9) => positive_inputs_18_9_port, 
                           A_signal(8) => positive_inputs_18_8_port, 
                           A_signal(7) => positive_inputs_18_7_port, 
                           A_signal(6) => positive_inputs_18_6_port, 
                           A_signal(5) => positive_inputs_18_5_port, 
                           A_signal(4) => positive_inputs_18_4_port, 
                           A_signal(3) => positive_inputs_18_3_port, 
                           A_signal(2) => positive_inputs_18_2_port, 
                           A_signal(1) => positive_inputs_18_1_port, 
                           A_signal(0) => n9, A_neg(63) => 
                           negative_inputs_18_63_port, A_neg(62) => 
                           negative_inputs_18_62_port, A_neg(61) => 
                           negative_inputs_18_61_port, A_neg(60) => 
                           negative_inputs_18_60_port, A_neg(59) => 
                           negative_inputs_18_59_port, A_neg(58) => 
                           negative_inputs_18_58_port, A_neg(57) => 
                           negative_inputs_18_57_port, A_neg(56) => 
                           negative_inputs_18_56_port, A_neg(55) => 
                           negative_inputs_18_55_port, A_neg(54) => 
                           negative_inputs_18_54_port, A_neg(53) => 
                           negative_inputs_18_53_port, A_neg(52) => 
                           negative_inputs_18_52_port, A_neg(51) => 
                           negative_inputs_18_51_port, A_neg(50) => 
                           negative_inputs_18_50_port, A_neg(49) => 
                           negative_inputs_18_49_port, A_neg(48) => 
                           negative_inputs_18_48_port, A_neg(47) => 
                           negative_inputs_18_47_port, A_neg(46) => 
                           negative_inputs_18_46_port, A_neg(45) => 
                           negative_inputs_18_45_port, A_neg(44) => 
                           negative_inputs_18_44_port, A_neg(43) => 
                           negative_inputs_18_43_port, A_neg(42) => 
                           negative_inputs_18_42_port, A_neg(41) => 
                           negative_inputs_18_41_port, A_neg(40) => 
                           negative_inputs_18_40_port, A_neg(39) => 
                           negative_inputs_18_39_port, A_neg(38) => 
                           negative_inputs_18_38_port, A_neg(37) => 
                           negative_inputs_18_37_port, A_neg(36) => 
                           negative_inputs_18_36_port, A_neg(35) => 
                           negative_inputs_18_35_port, A_neg(34) => 
                           negative_inputs_18_34_port, A_neg(33) => 
                           negative_inputs_18_33_port, A_neg(32) => 
                           negative_inputs_18_32_port, A_neg(31) => 
                           negative_inputs_18_31_port, A_neg(30) => 
                           negative_inputs_18_30_port, A_neg(29) => 
                           negative_inputs_18_29_port, A_neg(28) => 
                           negative_inputs_18_28_port, A_neg(27) => 
                           negative_inputs_18_27_port, A_neg(26) => 
                           negative_inputs_18_26_port, A_neg(25) => 
                           negative_inputs_18_25_port, A_neg(24) => 
                           negative_inputs_18_24_port, A_neg(23) => 
                           negative_inputs_18_23_port, A_neg(22) => 
                           negative_inputs_18_22_port, A_neg(21) => 
                           negative_inputs_18_21_port, A_neg(20) => 
                           negative_inputs_18_20_port, A_neg(19) => 
                           negative_inputs_18_19_port, A_neg(18) => 
                           negative_inputs_18_18_port, A_neg(17) => 
                           negative_inputs_18_17_port, A_neg(16) => 
                           negative_inputs_18_16_port, A_neg(15) => 
                           negative_inputs_18_15_port, A_neg(14) => 
                           negative_inputs_18_14_port, A_neg(13) => 
                           negative_inputs_18_13_port, A_neg(12) => 
                           negative_inputs_18_12_port, A_neg(11) => 
                           negative_inputs_18_11_port, A_neg(10) => 
                           negative_inputs_18_10_port, A_neg(9) => 
                           negative_inputs_18_9_port, A_neg(8) => 
                           negative_inputs_18_8_port, A_neg(7) => 
                           negative_inputs_18_7_port, A_neg(6) => 
                           negative_inputs_18_6_port, A_neg(5) => 
                           negative_inputs_18_5_port, A_neg(4) => 
                           negative_inputs_18_4_port, A_neg(3) => 
                           negative_inputs_18_3_port, A_neg(2) => 
                           negative_inputs_18_2_port, A_neg(1) => 
                           negative_inputs_18_1_port, A_neg(0) => n9, 
                           A_shifted(63) => positive_inputs_19_63_port, 
                           A_shifted(62) => positive_inputs_19_62_port, 
                           A_shifted(61) => positive_inputs_19_61_port, 
                           A_shifted(60) => positive_inputs_19_60_port, 
                           A_shifted(59) => positive_inputs_19_59_port, 
                           A_shifted(58) => positive_inputs_19_58_port, 
                           A_shifted(57) => positive_inputs_19_57_port, 
                           A_shifted(56) => positive_inputs_19_56_port, 
                           A_shifted(55) => positive_inputs_19_55_port, 
                           A_shifted(54) => positive_inputs_19_54_port, 
                           A_shifted(53) => positive_inputs_19_53_port, 
                           A_shifted(52) => positive_inputs_19_52_port, 
                           A_shifted(51) => positive_inputs_19_51_port, 
                           A_shifted(50) => positive_inputs_19_50_port, 
                           A_shifted(49) => positive_inputs_19_49_port, 
                           A_shifted(48) => positive_inputs_19_48_port, 
                           A_shifted(47) => positive_inputs_19_47_port, 
                           A_shifted(46) => positive_inputs_19_46_port, 
                           A_shifted(45) => positive_inputs_19_45_port, 
                           A_shifted(44) => positive_inputs_19_44_port, 
                           A_shifted(43) => positive_inputs_19_43_port, 
                           A_shifted(42) => positive_inputs_19_42_port, 
                           A_shifted(41) => positive_inputs_19_41_port, 
                           A_shifted(40) => positive_inputs_19_40_port, 
                           A_shifted(39) => positive_inputs_19_39_port, 
                           A_shifted(38) => positive_inputs_19_38_port, 
                           A_shifted(37) => positive_inputs_19_37_port, 
                           A_shifted(36) => positive_inputs_19_36_port, 
                           A_shifted(35) => positive_inputs_19_35_port, 
                           A_shifted(34) => positive_inputs_19_34_port, 
                           A_shifted(33) => positive_inputs_19_33_port, 
                           A_shifted(32) => positive_inputs_19_32_port, 
                           A_shifted(31) => positive_inputs_19_31_port, 
                           A_shifted(30) => positive_inputs_19_30_port, 
                           A_shifted(29) => positive_inputs_19_29_port, 
                           A_shifted(28) => positive_inputs_19_28_port, 
                           A_shifted(27) => positive_inputs_19_27_port, 
                           A_shifted(26) => positive_inputs_19_26_port, 
                           A_shifted(25) => positive_inputs_19_25_port, 
                           A_shifted(24) => positive_inputs_19_24_port, 
                           A_shifted(23) => positive_inputs_19_23_port, 
                           A_shifted(22) => positive_inputs_19_22_port, 
                           A_shifted(21) => positive_inputs_19_21_port, 
                           A_shifted(20) => positive_inputs_19_20_port, 
                           A_shifted(19) => positive_inputs_19_19_port, 
                           A_shifted(18) => positive_inputs_19_18_port, 
                           A_shifted(17) => positive_inputs_19_17_port, 
                           A_shifted(16) => positive_inputs_19_16_port, 
                           A_shifted(15) => positive_inputs_19_15_port, 
                           A_shifted(14) => positive_inputs_19_14_port, 
                           A_shifted(13) => positive_inputs_19_13_port, 
                           A_shifted(12) => positive_inputs_19_12_port, 
                           A_shifted(11) => positive_inputs_19_11_port, 
                           A_shifted(10) => positive_inputs_19_10_port, 
                           A_shifted(9) => positive_inputs_19_9_port, 
                           A_shifted(8) => positive_inputs_19_8_port, 
                           A_shifted(7) => positive_inputs_19_7_port, 
                           A_shifted(6) => positive_inputs_19_6_port, 
                           A_shifted(5) => positive_inputs_19_5_port, 
                           A_shifted(4) => positive_inputs_19_4_port, 
                           A_shifted(3) => positive_inputs_19_3_port, 
                           A_shifted(2) => positive_inputs_19_2_port, 
                           A_shifted(1) => positive_inputs_19_1_port, 
                           A_shifted(0) => n9, A_neg_shifted(63) => 
                           negative_inputs_19_63_port, A_neg_shifted(62) => 
                           negative_inputs_19_62_port, A_neg_shifted(61) => 
                           negative_inputs_19_61_port, A_neg_shifted(60) => 
                           negative_inputs_19_60_port, A_neg_shifted(59) => 
                           negative_inputs_19_59_port, A_neg_shifted(58) => 
                           negative_inputs_19_58_port, A_neg_shifted(57) => 
                           negative_inputs_19_57_port, A_neg_shifted(56) => 
                           negative_inputs_19_56_port, A_neg_shifted(55) => 
                           negative_inputs_19_55_port, A_neg_shifted(54) => 
                           negative_inputs_19_54_port, A_neg_shifted(53) => 
                           negative_inputs_19_53_port, A_neg_shifted(52) => 
                           negative_inputs_19_52_port, A_neg_shifted(51) => 
                           negative_inputs_19_51_port, A_neg_shifted(50) => 
                           negative_inputs_19_50_port, A_neg_shifted(49) => 
                           negative_inputs_19_49_port, A_neg_shifted(48) => 
                           negative_inputs_19_48_port, A_neg_shifted(47) => 
                           negative_inputs_19_47_port, A_neg_shifted(46) => 
                           negative_inputs_19_46_port, A_neg_shifted(45) => 
                           negative_inputs_19_45_port, A_neg_shifted(44) => 
                           negative_inputs_19_44_port, A_neg_shifted(43) => 
                           negative_inputs_19_43_port, A_neg_shifted(42) => 
                           negative_inputs_19_42_port, A_neg_shifted(41) => 
                           negative_inputs_19_41_port, A_neg_shifted(40) => 
                           negative_inputs_19_40_port, A_neg_shifted(39) => 
                           negative_inputs_19_39_port, A_neg_shifted(38) => 
                           negative_inputs_19_38_port, A_neg_shifted(37) => 
                           negative_inputs_19_37_port, A_neg_shifted(36) => 
                           negative_inputs_19_36_port, A_neg_shifted(35) => 
                           negative_inputs_19_35_port, A_neg_shifted(34) => 
                           negative_inputs_19_34_port, A_neg_shifted(33) => 
                           negative_inputs_19_33_port, A_neg_shifted(32) => 
                           negative_inputs_19_32_port, A_neg_shifted(31) => 
                           negative_inputs_19_31_port, A_neg_shifted(30) => 
                           negative_inputs_19_30_port, A_neg_shifted(29) => 
                           negative_inputs_19_29_port, A_neg_shifted(28) => 
                           negative_inputs_19_28_port, A_neg_shifted(27) => 
                           negative_inputs_19_27_port, A_neg_shifted(26) => 
                           negative_inputs_19_26_port, A_neg_shifted(25) => 
                           negative_inputs_19_25_port, A_neg_shifted(24) => 
                           negative_inputs_19_24_port, A_neg_shifted(23) => 
                           negative_inputs_19_23_port, A_neg_shifted(22) => 
                           negative_inputs_19_22_port, A_neg_shifted(21) => 
                           negative_inputs_19_21_port, A_neg_shifted(20) => 
                           negative_inputs_19_20_port, A_neg_shifted(19) => 
                           negative_inputs_19_19_port, A_neg_shifted(18) => 
                           negative_inputs_19_18_port, A_neg_shifted(17) => 
                           negative_inputs_19_17_port, A_neg_shifted(16) => 
                           negative_inputs_19_16_port, A_neg_shifted(15) => 
                           negative_inputs_19_15_port, A_neg_shifted(14) => 
                           negative_inputs_19_14_port, A_neg_shifted(13) => 
                           negative_inputs_19_13_port, A_neg_shifted(12) => 
                           negative_inputs_19_12_port, A_neg_shifted(11) => 
                           negative_inputs_19_11_port, A_neg_shifted(10) => 
                           negative_inputs_19_10_port, A_neg_shifted(9) => 
                           negative_inputs_19_9_port, A_neg_shifted(8) => 
                           negative_inputs_19_8_port, A_neg_shifted(7) => 
                           negative_inputs_19_7_port, A_neg_shifted(6) => 
                           negative_inputs_19_6_port, A_neg_shifted(5) => 
                           negative_inputs_19_5_port, A_neg_shifted(4) => 
                           negative_inputs_19_4_port, A_neg_shifted(3) => 
                           negative_inputs_19_3_port, A_neg_shifted(2) => 
                           negative_inputs_19_2_port, A_neg_shifted(1) => 
                           negative_inputs_19_1_port, A_neg_shifted(0) => n9, 
                           Sel(2) => sel_9_2_port, Sel(1) => sel_9_1_port, 
                           Sel(0) => sel_9_0_port, Y(63) => 
                           MuxOutputs_9_63_port, Y(62) => MuxOutputs_9_62_port,
                           Y(61) => MuxOutputs_9_61_port, Y(60) => 
                           MuxOutputs_9_60_port, Y(59) => MuxOutputs_9_59_port,
                           Y(58) => MuxOutputs_9_58_port, Y(57) => 
                           MuxOutputs_9_57_port, Y(56) => MuxOutputs_9_56_port,
                           Y(55) => MuxOutputs_9_55_port, Y(54) => 
                           MuxOutputs_9_54_port, Y(53) => MuxOutputs_9_53_port,
                           Y(52) => MuxOutputs_9_52_port, Y(51) => 
                           MuxOutputs_9_51_port, Y(50) => MuxOutputs_9_50_port,
                           Y(49) => MuxOutputs_9_49_port, Y(48) => 
                           MuxOutputs_9_48_port, Y(47) => MuxOutputs_9_47_port,
                           Y(46) => MuxOutputs_9_46_port, Y(45) => 
                           MuxOutputs_9_45_port, Y(44) => MuxOutputs_9_44_port,
                           Y(43) => MuxOutputs_9_43_port, Y(42) => 
                           MuxOutputs_9_42_port, Y(41) => MuxOutputs_9_41_port,
                           Y(40) => MuxOutputs_9_40_port, Y(39) => 
                           MuxOutputs_9_39_port, Y(38) => MuxOutputs_9_38_port,
                           Y(37) => MuxOutputs_9_37_port, Y(36) => 
                           MuxOutputs_9_36_port, Y(35) => MuxOutputs_9_35_port,
                           Y(34) => MuxOutputs_9_34_port, Y(33) => 
                           MuxOutputs_9_33_port, Y(32) => MuxOutputs_9_32_port,
                           Y(31) => MuxOutputs_9_31_port, Y(30) => 
                           MuxOutputs_9_30_port, Y(29) => MuxOutputs_9_29_port,
                           Y(28) => MuxOutputs_9_28_port, Y(27) => 
                           MuxOutputs_9_27_port, Y(26) => MuxOutputs_9_26_port,
                           Y(25) => MuxOutputs_9_25_port, Y(24) => 
                           MuxOutputs_9_24_port, Y(23) => MuxOutputs_9_23_port,
                           Y(22) => MuxOutputs_9_22_port, Y(21) => 
                           MuxOutputs_9_21_port, Y(20) => MuxOutputs_9_20_port,
                           Y(19) => MuxOutputs_9_19_port, Y(18) => 
                           MuxOutputs_9_18_port, Y(17) => MuxOutputs_9_17_port,
                           Y(16) => MuxOutputs_9_16_port, Y(15) => 
                           MuxOutputs_9_15_port, Y(14) => MuxOutputs_9_14_port,
                           Y(13) => MuxOutputs_9_13_port, Y(12) => 
                           MuxOutputs_9_12_port, Y(11) => MuxOutputs_9_11_port,
                           Y(10) => MuxOutputs_9_10_port, Y(9) => 
                           MuxOutputs_9_9_port, Y(8) => MuxOutputs_9_8_port, 
                           Y(7) => MuxOutputs_9_7_port, Y(6) => 
                           MuxOutputs_9_6_port, Y(5) => MuxOutputs_9_5_port, 
                           Y(4) => MuxOutputs_9_4_port, Y(3) => 
                           MuxOutputs_9_3_port, Y(2) => MuxOutputs_9_2_port, 
                           Y(1) => MuxOutputs_9_1_port, Y(0) => 
                           MuxOutputs_9_0_port);
   encoderI_10 : encoder_6 port map( pieceofB(2) => B(21), pieceofB(1) => B(20)
                           , pieceofB(0) => B(19), sel(2) => sel_10_2_port, 
                           sel(1) => sel_10_1_port, sel(0) => sel_10_0_port);
   MUXI_10 : MUX51_MuxNbit64_6 port map( zeroSignal(63) => X_Logic0_port, 
                           zeroSignal(62) => X_Logic0_port, zeroSignal(61) => 
                           X_Logic0_port, zeroSignal(60) => X_Logic0_port, 
                           zeroSignal(59) => X_Logic0_port, zeroSignal(58) => 
                           X_Logic0_port, zeroSignal(57) => X_Logic0_port, 
                           zeroSignal(56) => X_Logic0_port, zeroSignal(55) => 
                           X_Logic0_port, zeroSignal(54) => X_Logic0_port, 
                           zeroSignal(53) => X_Logic0_port, zeroSignal(52) => 
                           X_Logic0_port, zeroSignal(51) => X_Logic0_port, 
                           zeroSignal(50) => X_Logic0_port, zeroSignal(49) => 
                           X_Logic0_port, zeroSignal(48) => X_Logic0_port, 
                           zeroSignal(47) => X_Logic0_port, zeroSignal(46) => 
                           X_Logic0_port, zeroSignal(45) => X_Logic0_port, 
                           zeroSignal(44) => X_Logic0_port, zeroSignal(43) => 
                           X_Logic0_port, zeroSignal(42) => X_Logic0_port, 
                           zeroSignal(41) => X_Logic0_port, zeroSignal(40) => 
                           X_Logic0_port, zeroSignal(39) => X_Logic0_port, 
                           zeroSignal(38) => X_Logic0_port, zeroSignal(37) => 
                           X_Logic0_port, zeroSignal(36) => X_Logic0_port, 
                           zeroSignal(35) => X_Logic0_port, zeroSignal(34) => 
                           X_Logic0_port, zeroSignal(33) => X_Logic0_port, 
                           zeroSignal(32) => X_Logic0_port, zeroSignal(31) => 
                           X_Logic0_port, zeroSignal(30) => X_Logic0_port, 
                           zeroSignal(29) => X_Logic0_port, zeroSignal(28) => 
                           X_Logic0_port, zeroSignal(27) => X_Logic0_port, 
                           zeroSignal(26) => X_Logic0_port, zeroSignal(25) => 
                           X_Logic0_port, zeroSignal(24) => X_Logic0_port, 
                           zeroSignal(23) => X_Logic0_port, zeroSignal(22) => 
                           X_Logic0_port, zeroSignal(21) => X_Logic0_port, 
                           zeroSignal(20) => X_Logic0_port, zeroSignal(19) => 
                           X_Logic0_port, zeroSignal(18) => X_Logic0_port, 
                           zeroSignal(17) => X_Logic0_port, zeroSignal(16) => 
                           X_Logic0_port, zeroSignal(15) => X_Logic0_port, 
                           zeroSignal(14) => X_Logic0_port, zeroSignal(13) => 
                           X_Logic0_port, zeroSignal(12) => X_Logic0_port, 
                           zeroSignal(11) => X_Logic0_port, zeroSignal(10) => 
                           X_Logic0_port, zeroSignal(9) => X_Logic0_port, 
                           zeroSignal(8) => X_Logic0_port, zeroSignal(7) => 
                           X_Logic0_port, zeroSignal(6) => X_Logic0_port, 
                           zeroSignal(5) => X_Logic0_port, zeroSignal(4) => 
                           X_Logic0_port, zeroSignal(3) => X_Logic0_port, 
                           zeroSignal(2) => X_Logic0_port, zeroSignal(1) => 
                           X_Logic0_port, zeroSignal(0) => X_Logic0_port, 
                           A_signal(63) => positive_inputs_20_63_port, 
                           A_signal(62) => positive_inputs_20_62_port, 
                           A_signal(61) => positive_inputs_20_61_port, 
                           A_signal(60) => positive_inputs_20_60_port, 
                           A_signal(59) => positive_inputs_20_59_port, 
                           A_signal(58) => positive_inputs_20_58_port, 
                           A_signal(57) => positive_inputs_20_57_port, 
                           A_signal(56) => positive_inputs_20_56_port, 
                           A_signal(55) => positive_inputs_20_55_port, 
                           A_signal(54) => positive_inputs_20_54_port, 
                           A_signal(53) => positive_inputs_20_53_port, 
                           A_signal(52) => positive_inputs_20_52_port, 
                           A_signal(51) => positive_inputs_20_51_port, 
                           A_signal(50) => positive_inputs_20_50_port, 
                           A_signal(49) => positive_inputs_20_49_port, 
                           A_signal(48) => positive_inputs_20_48_port, 
                           A_signal(47) => positive_inputs_20_47_port, 
                           A_signal(46) => positive_inputs_20_46_port, 
                           A_signal(45) => positive_inputs_20_45_port, 
                           A_signal(44) => positive_inputs_20_44_port, 
                           A_signal(43) => positive_inputs_20_43_port, 
                           A_signal(42) => positive_inputs_20_42_port, 
                           A_signal(41) => positive_inputs_20_41_port, 
                           A_signal(40) => positive_inputs_20_40_port, 
                           A_signal(39) => positive_inputs_20_39_port, 
                           A_signal(38) => positive_inputs_20_38_port, 
                           A_signal(37) => positive_inputs_20_37_port, 
                           A_signal(36) => positive_inputs_20_36_port, 
                           A_signal(35) => positive_inputs_20_35_port, 
                           A_signal(34) => positive_inputs_20_34_port, 
                           A_signal(33) => positive_inputs_20_33_port, 
                           A_signal(32) => positive_inputs_20_32_port, 
                           A_signal(31) => positive_inputs_20_31_port, 
                           A_signal(30) => positive_inputs_20_30_port, 
                           A_signal(29) => positive_inputs_20_29_port, 
                           A_signal(28) => positive_inputs_20_28_port, 
                           A_signal(27) => positive_inputs_20_27_port, 
                           A_signal(26) => positive_inputs_20_26_port, 
                           A_signal(25) => positive_inputs_20_25_port, 
                           A_signal(24) => positive_inputs_20_24_port, 
                           A_signal(23) => positive_inputs_20_23_port, 
                           A_signal(22) => positive_inputs_20_22_port, 
                           A_signal(21) => positive_inputs_20_21_port, 
                           A_signal(20) => positive_inputs_20_20_port, 
                           A_signal(19) => positive_inputs_20_19_port, 
                           A_signal(18) => positive_inputs_20_18_port, 
                           A_signal(17) => positive_inputs_20_17_port, 
                           A_signal(16) => positive_inputs_20_16_port, 
                           A_signal(15) => positive_inputs_20_15_port, 
                           A_signal(14) => positive_inputs_20_14_port, 
                           A_signal(13) => positive_inputs_20_13_port, 
                           A_signal(12) => positive_inputs_20_12_port, 
                           A_signal(11) => positive_inputs_20_11_port, 
                           A_signal(10) => positive_inputs_20_10_port, 
                           A_signal(9) => positive_inputs_20_9_port, 
                           A_signal(8) => positive_inputs_20_8_port, 
                           A_signal(7) => positive_inputs_20_7_port, 
                           A_signal(6) => positive_inputs_20_6_port, 
                           A_signal(5) => positive_inputs_20_5_port, 
                           A_signal(4) => positive_inputs_20_4_port, 
                           A_signal(3) => positive_inputs_20_3_port, 
                           A_signal(2) => positive_inputs_20_2_port, 
                           A_signal(1) => positive_inputs_20_1_port, 
                           A_signal(0) => n9, A_neg(63) => 
                           negative_inputs_20_63_port, A_neg(62) => 
                           negative_inputs_20_62_port, A_neg(61) => 
                           negative_inputs_20_61_port, A_neg(60) => 
                           negative_inputs_20_60_port, A_neg(59) => 
                           negative_inputs_20_59_port, A_neg(58) => 
                           negative_inputs_20_58_port, A_neg(57) => 
                           negative_inputs_20_57_port, A_neg(56) => 
                           negative_inputs_20_56_port, A_neg(55) => 
                           negative_inputs_20_55_port, A_neg(54) => 
                           negative_inputs_20_54_port, A_neg(53) => 
                           negative_inputs_20_53_port, A_neg(52) => 
                           negative_inputs_20_52_port, A_neg(51) => 
                           negative_inputs_20_51_port, A_neg(50) => 
                           negative_inputs_20_50_port, A_neg(49) => 
                           negative_inputs_20_49_port, A_neg(48) => 
                           negative_inputs_20_48_port, A_neg(47) => 
                           negative_inputs_20_47_port, A_neg(46) => 
                           negative_inputs_20_46_port, A_neg(45) => 
                           negative_inputs_20_45_port, A_neg(44) => 
                           negative_inputs_20_44_port, A_neg(43) => 
                           negative_inputs_20_43_port, A_neg(42) => 
                           negative_inputs_20_42_port, A_neg(41) => 
                           negative_inputs_20_41_port, A_neg(40) => 
                           negative_inputs_20_40_port, A_neg(39) => 
                           negative_inputs_20_39_port, A_neg(38) => 
                           negative_inputs_20_38_port, A_neg(37) => 
                           negative_inputs_20_37_port, A_neg(36) => 
                           negative_inputs_20_36_port, A_neg(35) => 
                           negative_inputs_20_35_port, A_neg(34) => 
                           negative_inputs_20_34_port, A_neg(33) => 
                           negative_inputs_20_33_port, A_neg(32) => 
                           negative_inputs_20_32_port, A_neg(31) => 
                           negative_inputs_20_31_port, A_neg(30) => 
                           negative_inputs_20_30_port, A_neg(29) => 
                           negative_inputs_20_29_port, A_neg(28) => 
                           negative_inputs_20_28_port, A_neg(27) => 
                           negative_inputs_20_27_port, A_neg(26) => 
                           negative_inputs_20_26_port, A_neg(25) => 
                           negative_inputs_20_25_port, A_neg(24) => 
                           negative_inputs_20_24_port, A_neg(23) => 
                           negative_inputs_20_23_port, A_neg(22) => 
                           negative_inputs_20_22_port, A_neg(21) => 
                           negative_inputs_20_21_port, A_neg(20) => 
                           negative_inputs_20_20_port, A_neg(19) => 
                           negative_inputs_20_19_port, A_neg(18) => 
                           negative_inputs_20_18_port, A_neg(17) => 
                           negative_inputs_20_17_port, A_neg(16) => 
                           negative_inputs_20_16_port, A_neg(15) => 
                           negative_inputs_20_15_port, A_neg(14) => 
                           negative_inputs_20_14_port, A_neg(13) => 
                           negative_inputs_20_13_port, A_neg(12) => 
                           negative_inputs_20_12_port, A_neg(11) => 
                           negative_inputs_20_11_port, A_neg(10) => 
                           negative_inputs_20_10_port, A_neg(9) => 
                           negative_inputs_20_9_port, A_neg(8) => 
                           negative_inputs_20_8_port, A_neg(7) => 
                           negative_inputs_20_7_port, A_neg(6) => 
                           negative_inputs_20_6_port, A_neg(5) => 
                           negative_inputs_20_5_port, A_neg(4) => 
                           negative_inputs_20_4_port, A_neg(3) => 
                           negative_inputs_20_3_port, A_neg(2) => 
                           negative_inputs_20_2_port, A_neg(1) => 
                           negative_inputs_20_1_port, A_neg(0) => n9, 
                           A_shifted(63) => positive_inputs_21_63_port, 
                           A_shifted(62) => positive_inputs_21_62_port, 
                           A_shifted(61) => positive_inputs_21_61_port, 
                           A_shifted(60) => positive_inputs_21_60_port, 
                           A_shifted(59) => positive_inputs_21_59_port, 
                           A_shifted(58) => positive_inputs_21_58_port, 
                           A_shifted(57) => positive_inputs_21_57_port, 
                           A_shifted(56) => positive_inputs_21_56_port, 
                           A_shifted(55) => positive_inputs_21_55_port, 
                           A_shifted(54) => positive_inputs_21_54_port, 
                           A_shifted(53) => positive_inputs_21_53_port, 
                           A_shifted(52) => positive_inputs_21_52_port, 
                           A_shifted(51) => positive_inputs_21_51_port, 
                           A_shifted(50) => positive_inputs_21_50_port, 
                           A_shifted(49) => positive_inputs_21_49_port, 
                           A_shifted(48) => positive_inputs_21_48_port, 
                           A_shifted(47) => positive_inputs_21_47_port, 
                           A_shifted(46) => positive_inputs_21_46_port, 
                           A_shifted(45) => positive_inputs_21_45_port, 
                           A_shifted(44) => positive_inputs_21_44_port, 
                           A_shifted(43) => positive_inputs_21_43_port, 
                           A_shifted(42) => positive_inputs_21_42_port, 
                           A_shifted(41) => positive_inputs_21_41_port, 
                           A_shifted(40) => positive_inputs_21_40_port, 
                           A_shifted(39) => positive_inputs_21_39_port, 
                           A_shifted(38) => positive_inputs_21_38_port, 
                           A_shifted(37) => positive_inputs_21_37_port, 
                           A_shifted(36) => positive_inputs_21_36_port, 
                           A_shifted(35) => positive_inputs_21_35_port, 
                           A_shifted(34) => positive_inputs_21_34_port, 
                           A_shifted(33) => positive_inputs_21_33_port, 
                           A_shifted(32) => positive_inputs_21_32_port, 
                           A_shifted(31) => positive_inputs_21_31_port, 
                           A_shifted(30) => positive_inputs_21_30_port, 
                           A_shifted(29) => positive_inputs_21_29_port, 
                           A_shifted(28) => positive_inputs_21_28_port, 
                           A_shifted(27) => positive_inputs_21_27_port, 
                           A_shifted(26) => positive_inputs_21_26_port, 
                           A_shifted(25) => positive_inputs_21_25_port, 
                           A_shifted(24) => positive_inputs_21_24_port, 
                           A_shifted(23) => positive_inputs_21_23_port, 
                           A_shifted(22) => positive_inputs_21_22_port, 
                           A_shifted(21) => positive_inputs_21_21_port, 
                           A_shifted(20) => positive_inputs_21_20_port, 
                           A_shifted(19) => positive_inputs_21_19_port, 
                           A_shifted(18) => positive_inputs_21_18_port, 
                           A_shifted(17) => positive_inputs_21_17_port, 
                           A_shifted(16) => positive_inputs_21_16_port, 
                           A_shifted(15) => positive_inputs_21_15_port, 
                           A_shifted(14) => positive_inputs_21_14_port, 
                           A_shifted(13) => positive_inputs_21_13_port, 
                           A_shifted(12) => positive_inputs_21_12_port, 
                           A_shifted(11) => positive_inputs_21_11_port, 
                           A_shifted(10) => positive_inputs_21_10_port, 
                           A_shifted(9) => positive_inputs_21_9_port, 
                           A_shifted(8) => positive_inputs_21_8_port, 
                           A_shifted(7) => positive_inputs_21_7_port, 
                           A_shifted(6) => positive_inputs_21_6_port, 
                           A_shifted(5) => positive_inputs_21_5_port, 
                           A_shifted(4) => positive_inputs_21_4_port, 
                           A_shifted(3) => positive_inputs_21_3_port, 
                           A_shifted(2) => positive_inputs_21_2_port, 
                           A_shifted(1) => positive_inputs_21_1_port, 
                           A_shifted(0) => n9, A_neg_shifted(63) => 
                           negative_inputs_21_63_port, A_neg_shifted(62) => 
                           negative_inputs_21_62_port, A_neg_shifted(61) => 
                           negative_inputs_21_61_port, A_neg_shifted(60) => 
                           negative_inputs_21_60_port, A_neg_shifted(59) => 
                           negative_inputs_21_59_port, A_neg_shifted(58) => 
                           negative_inputs_21_58_port, A_neg_shifted(57) => 
                           negative_inputs_21_57_port, A_neg_shifted(56) => 
                           negative_inputs_21_56_port, A_neg_shifted(55) => 
                           negative_inputs_21_55_port, A_neg_shifted(54) => 
                           negative_inputs_21_54_port, A_neg_shifted(53) => 
                           negative_inputs_21_53_port, A_neg_shifted(52) => 
                           negative_inputs_21_52_port, A_neg_shifted(51) => 
                           negative_inputs_21_51_port, A_neg_shifted(50) => 
                           negative_inputs_21_50_port, A_neg_shifted(49) => 
                           negative_inputs_21_49_port, A_neg_shifted(48) => 
                           negative_inputs_21_48_port, A_neg_shifted(47) => 
                           negative_inputs_21_47_port, A_neg_shifted(46) => 
                           negative_inputs_21_46_port, A_neg_shifted(45) => 
                           negative_inputs_21_45_port, A_neg_shifted(44) => 
                           negative_inputs_21_44_port, A_neg_shifted(43) => 
                           negative_inputs_21_43_port, A_neg_shifted(42) => 
                           negative_inputs_21_42_port, A_neg_shifted(41) => 
                           negative_inputs_21_41_port, A_neg_shifted(40) => 
                           negative_inputs_21_40_port, A_neg_shifted(39) => 
                           negative_inputs_21_39_port, A_neg_shifted(38) => 
                           negative_inputs_21_38_port, A_neg_shifted(37) => 
                           negative_inputs_21_37_port, A_neg_shifted(36) => 
                           negative_inputs_21_36_port, A_neg_shifted(35) => 
                           negative_inputs_21_35_port, A_neg_shifted(34) => 
                           negative_inputs_21_34_port, A_neg_shifted(33) => 
                           negative_inputs_21_33_port, A_neg_shifted(32) => 
                           negative_inputs_21_32_port, A_neg_shifted(31) => 
                           negative_inputs_21_31_port, A_neg_shifted(30) => 
                           negative_inputs_21_30_port, A_neg_shifted(29) => 
                           negative_inputs_21_29_port, A_neg_shifted(28) => 
                           negative_inputs_21_28_port, A_neg_shifted(27) => 
                           negative_inputs_21_27_port, A_neg_shifted(26) => 
                           negative_inputs_21_26_port, A_neg_shifted(25) => 
                           negative_inputs_21_25_port, A_neg_shifted(24) => 
                           negative_inputs_21_24_port, A_neg_shifted(23) => 
                           negative_inputs_21_23_port, A_neg_shifted(22) => 
                           negative_inputs_21_22_port, A_neg_shifted(21) => 
                           negative_inputs_21_21_port, A_neg_shifted(20) => 
                           negative_inputs_21_20_port, A_neg_shifted(19) => 
                           negative_inputs_21_19_port, A_neg_shifted(18) => 
                           negative_inputs_21_18_port, A_neg_shifted(17) => 
                           negative_inputs_21_17_port, A_neg_shifted(16) => 
                           negative_inputs_21_16_port, A_neg_shifted(15) => 
                           negative_inputs_21_15_port, A_neg_shifted(14) => 
                           negative_inputs_21_14_port, A_neg_shifted(13) => 
                           negative_inputs_21_13_port, A_neg_shifted(12) => 
                           negative_inputs_21_12_port, A_neg_shifted(11) => 
                           negative_inputs_21_11_port, A_neg_shifted(10) => 
                           negative_inputs_21_10_port, A_neg_shifted(9) => 
                           negative_inputs_21_9_port, A_neg_shifted(8) => 
                           negative_inputs_21_8_port, A_neg_shifted(7) => 
                           negative_inputs_21_7_port, A_neg_shifted(6) => 
                           negative_inputs_21_6_port, A_neg_shifted(5) => 
                           negative_inputs_21_5_port, A_neg_shifted(4) => 
                           negative_inputs_21_4_port, A_neg_shifted(3) => 
                           negative_inputs_21_3_port, A_neg_shifted(2) => 
                           negative_inputs_21_2_port, A_neg_shifted(1) => 
                           negative_inputs_21_1_port, A_neg_shifted(0) => n9, 
                           Sel(2) => sel_10_2_port, Sel(1) => sel_10_1_port, 
                           Sel(0) => sel_10_0_port, Y(63) => 
                           MuxOutputs_10_63_port, Y(62) => 
                           MuxOutputs_10_62_port, Y(61) => 
                           MuxOutputs_10_61_port, Y(60) => 
                           MuxOutputs_10_60_port, Y(59) => 
                           MuxOutputs_10_59_port, Y(58) => 
                           MuxOutputs_10_58_port, Y(57) => 
                           MuxOutputs_10_57_port, Y(56) => 
                           MuxOutputs_10_56_port, Y(55) => 
                           MuxOutputs_10_55_port, Y(54) => 
                           MuxOutputs_10_54_port, Y(53) => 
                           MuxOutputs_10_53_port, Y(52) => 
                           MuxOutputs_10_52_port, Y(51) => 
                           MuxOutputs_10_51_port, Y(50) => 
                           MuxOutputs_10_50_port, Y(49) => 
                           MuxOutputs_10_49_port, Y(48) => 
                           MuxOutputs_10_48_port, Y(47) => 
                           MuxOutputs_10_47_port, Y(46) => 
                           MuxOutputs_10_46_port, Y(45) => 
                           MuxOutputs_10_45_port, Y(44) => 
                           MuxOutputs_10_44_port, Y(43) => 
                           MuxOutputs_10_43_port, Y(42) => 
                           MuxOutputs_10_42_port, Y(41) => 
                           MuxOutputs_10_41_port, Y(40) => 
                           MuxOutputs_10_40_port, Y(39) => 
                           MuxOutputs_10_39_port, Y(38) => 
                           MuxOutputs_10_38_port, Y(37) => 
                           MuxOutputs_10_37_port, Y(36) => 
                           MuxOutputs_10_36_port, Y(35) => 
                           MuxOutputs_10_35_port, Y(34) => 
                           MuxOutputs_10_34_port, Y(33) => 
                           MuxOutputs_10_33_port, Y(32) => 
                           MuxOutputs_10_32_port, Y(31) => 
                           MuxOutputs_10_31_port, Y(30) => 
                           MuxOutputs_10_30_port, Y(29) => 
                           MuxOutputs_10_29_port, Y(28) => 
                           MuxOutputs_10_28_port, Y(27) => 
                           MuxOutputs_10_27_port, Y(26) => 
                           MuxOutputs_10_26_port, Y(25) => 
                           MuxOutputs_10_25_port, Y(24) => 
                           MuxOutputs_10_24_port, Y(23) => 
                           MuxOutputs_10_23_port, Y(22) => 
                           MuxOutputs_10_22_port, Y(21) => 
                           MuxOutputs_10_21_port, Y(20) => 
                           MuxOutputs_10_20_port, Y(19) => 
                           MuxOutputs_10_19_port, Y(18) => 
                           MuxOutputs_10_18_port, Y(17) => 
                           MuxOutputs_10_17_port, Y(16) => 
                           MuxOutputs_10_16_port, Y(15) => 
                           MuxOutputs_10_15_port, Y(14) => 
                           MuxOutputs_10_14_port, Y(13) => 
                           MuxOutputs_10_13_port, Y(12) => 
                           MuxOutputs_10_12_port, Y(11) => 
                           MuxOutputs_10_11_port, Y(10) => 
                           MuxOutputs_10_10_port, Y(9) => MuxOutputs_10_9_port,
                           Y(8) => MuxOutputs_10_8_port, Y(7) => 
                           MuxOutputs_10_7_port, Y(6) => MuxOutputs_10_6_port, 
                           Y(5) => MuxOutputs_10_5_port, Y(4) => 
                           MuxOutputs_10_4_port, Y(3) => MuxOutputs_10_3_port, 
                           Y(2) => MuxOutputs_10_2_port, Y(1) => 
                           MuxOutputs_10_1_port, Y(0) => MuxOutputs_10_0_port);
   encoderI_11 : encoder_5 port map( pieceofB(2) => B(23), pieceofB(1) => B(22)
                           , pieceofB(0) => B(21), sel(2) => sel_11_2_port, 
                           sel(1) => sel_11_1_port, sel(0) => sel_11_0_port);
   MUXI_11 : MUX51_MuxNbit64_5 port map( zeroSignal(63) => X_Logic0_port, 
                           zeroSignal(62) => X_Logic0_port, zeroSignal(61) => 
                           X_Logic0_port, zeroSignal(60) => X_Logic0_port, 
                           zeroSignal(59) => X_Logic0_port, zeroSignal(58) => 
                           X_Logic0_port, zeroSignal(57) => X_Logic0_port, 
                           zeroSignal(56) => X_Logic0_port, zeroSignal(55) => 
                           X_Logic0_port, zeroSignal(54) => X_Logic0_port, 
                           zeroSignal(53) => X_Logic0_port, zeroSignal(52) => 
                           X_Logic0_port, zeroSignal(51) => X_Logic0_port, 
                           zeroSignal(50) => X_Logic0_port, zeroSignal(49) => 
                           X_Logic0_port, zeroSignal(48) => X_Logic0_port, 
                           zeroSignal(47) => X_Logic0_port, zeroSignal(46) => 
                           X_Logic0_port, zeroSignal(45) => X_Logic0_port, 
                           zeroSignal(44) => X_Logic0_port, zeroSignal(43) => 
                           X_Logic0_port, zeroSignal(42) => X_Logic0_port, 
                           zeroSignal(41) => X_Logic0_port, zeroSignal(40) => 
                           X_Logic0_port, zeroSignal(39) => X_Logic0_port, 
                           zeroSignal(38) => X_Logic0_port, zeroSignal(37) => 
                           X_Logic0_port, zeroSignal(36) => X_Logic0_port, 
                           zeroSignal(35) => X_Logic0_port, zeroSignal(34) => 
                           X_Logic0_port, zeroSignal(33) => X_Logic0_port, 
                           zeroSignal(32) => X_Logic0_port, zeroSignal(31) => 
                           X_Logic0_port, zeroSignal(30) => X_Logic0_port, 
                           zeroSignal(29) => X_Logic0_port, zeroSignal(28) => 
                           X_Logic0_port, zeroSignal(27) => X_Logic0_port, 
                           zeroSignal(26) => X_Logic0_port, zeroSignal(25) => 
                           X_Logic0_port, zeroSignal(24) => X_Logic0_port, 
                           zeroSignal(23) => X_Logic0_port, zeroSignal(22) => 
                           X_Logic0_port, zeroSignal(21) => X_Logic0_port, 
                           zeroSignal(20) => X_Logic0_port, zeroSignal(19) => 
                           X_Logic0_port, zeroSignal(18) => X_Logic0_port, 
                           zeroSignal(17) => X_Logic0_port, zeroSignal(16) => 
                           X_Logic0_port, zeroSignal(15) => X_Logic0_port, 
                           zeroSignal(14) => X_Logic0_port, zeroSignal(13) => 
                           X_Logic0_port, zeroSignal(12) => X_Logic0_port, 
                           zeroSignal(11) => X_Logic0_port, zeroSignal(10) => 
                           X_Logic0_port, zeroSignal(9) => X_Logic0_port, 
                           zeroSignal(8) => X_Logic0_port, zeroSignal(7) => 
                           X_Logic0_port, zeroSignal(6) => X_Logic0_port, 
                           zeroSignal(5) => X_Logic0_port, zeroSignal(4) => 
                           X_Logic0_port, zeroSignal(3) => X_Logic0_port, 
                           zeroSignal(2) => X_Logic0_port, zeroSignal(1) => 
                           X_Logic0_port, zeroSignal(0) => X_Logic0_port, 
                           A_signal(63) => positive_inputs_22_63_port, 
                           A_signal(62) => positive_inputs_22_62_port, 
                           A_signal(61) => positive_inputs_22_61_port, 
                           A_signal(60) => positive_inputs_22_60_port, 
                           A_signal(59) => positive_inputs_22_59_port, 
                           A_signal(58) => positive_inputs_22_58_port, 
                           A_signal(57) => positive_inputs_22_57_port, 
                           A_signal(56) => positive_inputs_22_56_port, 
                           A_signal(55) => positive_inputs_22_55_port, 
                           A_signal(54) => positive_inputs_22_54_port, 
                           A_signal(53) => positive_inputs_22_53_port, 
                           A_signal(52) => positive_inputs_22_52_port, 
                           A_signal(51) => positive_inputs_22_51_port, 
                           A_signal(50) => positive_inputs_22_50_port, 
                           A_signal(49) => positive_inputs_22_49_port, 
                           A_signal(48) => positive_inputs_22_48_port, 
                           A_signal(47) => positive_inputs_22_47_port, 
                           A_signal(46) => positive_inputs_22_46_port, 
                           A_signal(45) => positive_inputs_22_45_port, 
                           A_signal(44) => positive_inputs_22_44_port, 
                           A_signal(43) => positive_inputs_22_43_port, 
                           A_signal(42) => positive_inputs_22_42_port, 
                           A_signal(41) => positive_inputs_22_41_port, 
                           A_signal(40) => positive_inputs_22_40_port, 
                           A_signal(39) => positive_inputs_22_39_port, 
                           A_signal(38) => positive_inputs_22_38_port, 
                           A_signal(37) => positive_inputs_22_37_port, 
                           A_signal(36) => positive_inputs_22_36_port, 
                           A_signal(35) => positive_inputs_22_35_port, 
                           A_signal(34) => positive_inputs_22_34_port, 
                           A_signal(33) => positive_inputs_22_33_port, 
                           A_signal(32) => positive_inputs_22_32_port, 
                           A_signal(31) => positive_inputs_22_31_port, 
                           A_signal(30) => positive_inputs_22_30_port, 
                           A_signal(29) => positive_inputs_22_29_port, 
                           A_signal(28) => positive_inputs_22_28_port, 
                           A_signal(27) => positive_inputs_22_27_port, 
                           A_signal(26) => positive_inputs_22_26_port, 
                           A_signal(25) => positive_inputs_22_25_port, 
                           A_signal(24) => positive_inputs_22_24_port, 
                           A_signal(23) => positive_inputs_22_23_port, 
                           A_signal(22) => positive_inputs_22_22_port, 
                           A_signal(21) => positive_inputs_22_21_port, 
                           A_signal(20) => positive_inputs_22_20_port, 
                           A_signal(19) => positive_inputs_22_19_port, 
                           A_signal(18) => positive_inputs_22_18_port, 
                           A_signal(17) => positive_inputs_22_17_port, 
                           A_signal(16) => positive_inputs_22_16_port, 
                           A_signal(15) => positive_inputs_22_15_port, 
                           A_signal(14) => positive_inputs_22_14_port, 
                           A_signal(13) => positive_inputs_22_13_port, 
                           A_signal(12) => positive_inputs_22_12_port, 
                           A_signal(11) => positive_inputs_22_11_port, 
                           A_signal(10) => positive_inputs_22_10_port, 
                           A_signal(9) => positive_inputs_22_9_port, 
                           A_signal(8) => positive_inputs_22_8_port, 
                           A_signal(7) => positive_inputs_22_7_port, 
                           A_signal(6) => positive_inputs_22_6_port, 
                           A_signal(5) => positive_inputs_22_5_port, 
                           A_signal(4) => positive_inputs_22_4_port, 
                           A_signal(3) => positive_inputs_22_3_port, 
                           A_signal(2) => positive_inputs_22_2_port, 
                           A_signal(1) => positive_inputs_22_1_port, 
                           A_signal(0) => n9, A_neg(63) => 
                           negative_inputs_22_63_port, A_neg(62) => 
                           negative_inputs_22_62_port, A_neg(61) => 
                           negative_inputs_22_61_port, A_neg(60) => 
                           negative_inputs_22_60_port, A_neg(59) => 
                           negative_inputs_22_59_port, A_neg(58) => 
                           negative_inputs_22_58_port, A_neg(57) => 
                           negative_inputs_22_57_port, A_neg(56) => 
                           negative_inputs_22_56_port, A_neg(55) => 
                           negative_inputs_22_55_port, A_neg(54) => 
                           negative_inputs_22_54_port, A_neg(53) => 
                           negative_inputs_22_53_port, A_neg(52) => 
                           negative_inputs_22_52_port, A_neg(51) => 
                           negative_inputs_22_51_port, A_neg(50) => 
                           negative_inputs_22_50_port, A_neg(49) => 
                           negative_inputs_22_49_port, A_neg(48) => 
                           negative_inputs_22_48_port, A_neg(47) => 
                           negative_inputs_22_47_port, A_neg(46) => 
                           negative_inputs_22_46_port, A_neg(45) => 
                           negative_inputs_22_45_port, A_neg(44) => 
                           negative_inputs_22_44_port, A_neg(43) => 
                           negative_inputs_22_43_port, A_neg(42) => 
                           negative_inputs_22_42_port, A_neg(41) => 
                           negative_inputs_22_41_port, A_neg(40) => 
                           negative_inputs_22_40_port, A_neg(39) => 
                           negative_inputs_22_39_port, A_neg(38) => 
                           negative_inputs_22_38_port, A_neg(37) => 
                           negative_inputs_22_37_port, A_neg(36) => 
                           negative_inputs_22_36_port, A_neg(35) => 
                           negative_inputs_22_35_port, A_neg(34) => 
                           negative_inputs_22_34_port, A_neg(33) => 
                           negative_inputs_22_33_port, A_neg(32) => 
                           negative_inputs_22_32_port, A_neg(31) => 
                           negative_inputs_22_31_port, A_neg(30) => 
                           negative_inputs_22_30_port, A_neg(29) => 
                           negative_inputs_22_29_port, A_neg(28) => 
                           negative_inputs_22_28_port, A_neg(27) => 
                           negative_inputs_22_27_port, A_neg(26) => 
                           negative_inputs_22_26_port, A_neg(25) => 
                           negative_inputs_22_25_port, A_neg(24) => 
                           negative_inputs_22_24_port, A_neg(23) => 
                           negative_inputs_22_23_port, A_neg(22) => 
                           negative_inputs_22_22_port, A_neg(21) => 
                           negative_inputs_22_21_port, A_neg(20) => 
                           negative_inputs_22_20_port, A_neg(19) => 
                           negative_inputs_22_19_port, A_neg(18) => 
                           negative_inputs_22_18_port, A_neg(17) => 
                           negative_inputs_22_17_port, A_neg(16) => 
                           negative_inputs_22_16_port, A_neg(15) => 
                           negative_inputs_22_15_port, A_neg(14) => 
                           negative_inputs_22_14_port, A_neg(13) => 
                           negative_inputs_22_13_port, A_neg(12) => 
                           negative_inputs_22_12_port, A_neg(11) => 
                           negative_inputs_22_11_port, A_neg(10) => 
                           negative_inputs_22_10_port, A_neg(9) => 
                           negative_inputs_22_9_port, A_neg(8) => 
                           negative_inputs_22_8_port, A_neg(7) => 
                           negative_inputs_22_7_port, A_neg(6) => 
                           negative_inputs_22_6_port, A_neg(5) => 
                           negative_inputs_22_5_port, A_neg(4) => 
                           negative_inputs_22_4_port, A_neg(3) => 
                           negative_inputs_22_3_port, A_neg(2) => 
                           negative_inputs_22_2_port, A_neg(1) => 
                           negative_inputs_22_1_port, A_neg(0) => n9, 
                           A_shifted(63) => positive_inputs_23_63_port, 
                           A_shifted(62) => positive_inputs_23_62_port, 
                           A_shifted(61) => positive_inputs_23_61_port, 
                           A_shifted(60) => positive_inputs_23_60_port, 
                           A_shifted(59) => positive_inputs_23_59_port, 
                           A_shifted(58) => positive_inputs_23_58_port, 
                           A_shifted(57) => positive_inputs_23_57_port, 
                           A_shifted(56) => positive_inputs_23_56_port, 
                           A_shifted(55) => positive_inputs_23_55_port, 
                           A_shifted(54) => positive_inputs_23_54_port, 
                           A_shifted(53) => positive_inputs_23_53_port, 
                           A_shifted(52) => positive_inputs_23_52_port, 
                           A_shifted(51) => positive_inputs_23_51_port, 
                           A_shifted(50) => positive_inputs_23_50_port, 
                           A_shifted(49) => positive_inputs_23_49_port, 
                           A_shifted(48) => positive_inputs_23_48_port, 
                           A_shifted(47) => positive_inputs_23_47_port, 
                           A_shifted(46) => positive_inputs_23_46_port, 
                           A_shifted(45) => positive_inputs_23_45_port, 
                           A_shifted(44) => positive_inputs_23_44_port, 
                           A_shifted(43) => positive_inputs_23_43_port, 
                           A_shifted(42) => positive_inputs_23_42_port, 
                           A_shifted(41) => positive_inputs_23_41_port, 
                           A_shifted(40) => positive_inputs_23_40_port, 
                           A_shifted(39) => positive_inputs_23_39_port, 
                           A_shifted(38) => positive_inputs_23_38_port, 
                           A_shifted(37) => positive_inputs_23_37_port, 
                           A_shifted(36) => positive_inputs_23_36_port, 
                           A_shifted(35) => positive_inputs_23_35_port, 
                           A_shifted(34) => positive_inputs_23_34_port, 
                           A_shifted(33) => positive_inputs_23_33_port, 
                           A_shifted(32) => positive_inputs_23_32_port, 
                           A_shifted(31) => positive_inputs_23_31_port, 
                           A_shifted(30) => positive_inputs_23_30_port, 
                           A_shifted(29) => positive_inputs_23_29_port, 
                           A_shifted(28) => positive_inputs_23_28_port, 
                           A_shifted(27) => positive_inputs_23_27_port, 
                           A_shifted(26) => positive_inputs_23_26_port, 
                           A_shifted(25) => positive_inputs_23_25_port, 
                           A_shifted(24) => positive_inputs_23_24_port, 
                           A_shifted(23) => positive_inputs_23_23_port, 
                           A_shifted(22) => positive_inputs_23_22_port, 
                           A_shifted(21) => positive_inputs_23_21_port, 
                           A_shifted(20) => positive_inputs_23_20_port, 
                           A_shifted(19) => positive_inputs_23_19_port, 
                           A_shifted(18) => positive_inputs_23_18_port, 
                           A_shifted(17) => positive_inputs_23_17_port, 
                           A_shifted(16) => positive_inputs_23_16_port, 
                           A_shifted(15) => positive_inputs_23_15_port, 
                           A_shifted(14) => positive_inputs_23_14_port, 
                           A_shifted(13) => positive_inputs_23_13_port, 
                           A_shifted(12) => positive_inputs_23_12_port, 
                           A_shifted(11) => positive_inputs_23_11_port, 
                           A_shifted(10) => positive_inputs_23_10_port, 
                           A_shifted(9) => positive_inputs_23_9_port, 
                           A_shifted(8) => positive_inputs_23_8_port, 
                           A_shifted(7) => positive_inputs_23_7_port, 
                           A_shifted(6) => positive_inputs_23_6_port, 
                           A_shifted(5) => positive_inputs_23_5_port, 
                           A_shifted(4) => positive_inputs_23_4_port, 
                           A_shifted(3) => positive_inputs_23_3_port, 
                           A_shifted(2) => positive_inputs_23_2_port, 
                           A_shifted(1) => positive_inputs_23_1_port, 
                           A_shifted(0) => n9, A_neg_shifted(63) => 
                           negative_inputs_23_63_port, A_neg_shifted(62) => 
                           negative_inputs_23_62_port, A_neg_shifted(61) => 
                           negative_inputs_23_61_port, A_neg_shifted(60) => 
                           negative_inputs_23_60_port, A_neg_shifted(59) => 
                           negative_inputs_23_59_port, A_neg_shifted(58) => 
                           negative_inputs_23_58_port, A_neg_shifted(57) => 
                           negative_inputs_23_57_port, A_neg_shifted(56) => 
                           negative_inputs_23_56_port, A_neg_shifted(55) => 
                           negative_inputs_23_55_port, A_neg_shifted(54) => 
                           negative_inputs_23_54_port, A_neg_shifted(53) => 
                           negative_inputs_23_53_port, A_neg_shifted(52) => 
                           negative_inputs_23_52_port, A_neg_shifted(51) => 
                           negative_inputs_23_51_port, A_neg_shifted(50) => 
                           negative_inputs_23_50_port, A_neg_shifted(49) => 
                           negative_inputs_23_49_port, A_neg_shifted(48) => 
                           negative_inputs_23_48_port, A_neg_shifted(47) => 
                           negative_inputs_23_47_port, A_neg_shifted(46) => 
                           negative_inputs_23_46_port, A_neg_shifted(45) => 
                           negative_inputs_23_45_port, A_neg_shifted(44) => 
                           negative_inputs_23_44_port, A_neg_shifted(43) => 
                           negative_inputs_23_43_port, A_neg_shifted(42) => 
                           negative_inputs_23_42_port, A_neg_shifted(41) => 
                           negative_inputs_23_41_port, A_neg_shifted(40) => 
                           negative_inputs_23_40_port, A_neg_shifted(39) => 
                           negative_inputs_23_39_port, A_neg_shifted(38) => 
                           negative_inputs_23_38_port, A_neg_shifted(37) => 
                           negative_inputs_23_37_port, A_neg_shifted(36) => 
                           negative_inputs_23_36_port, A_neg_shifted(35) => 
                           negative_inputs_23_35_port, A_neg_shifted(34) => 
                           negative_inputs_23_34_port, A_neg_shifted(33) => 
                           negative_inputs_23_33_port, A_neg_shifted(32) => 
                           negative_inputs_23_32_port, A_neg_shifted(31) => 
                           negative_inputs_23_31_port, A_neg_shifted(30) => 
                           negative_inputs_23_30_port, A_neg_shifted(29) => 
                           negative_inputs_23_29_port, A_neg_shifted(28) => 
                           negative_inputs_23_28_port, A_neg_shifted(27) => 
                           negative_inputs_23_27_port, A_neg_shifted(26) => 
                           negative_inputs_23_26_port, A_neg_shifted(25) => 
                           negative_inputs_23_25_port, A_neg_shifted(24) => 
                           negative_inputs_23_24_port, A_neg_shifted(23) => 
                           negative_inputs_23_23_port, A_neg_shifted(22) => 
                           negative_inputs_23_22_port, A_neg_shifted(21) => 
                           negative_inputs_23_21_port, A_neg_shifted(20) => 
                           negative_inputs_23_20_port, A_neg_shifted(19) => 
                           negative_inputs_23_19_port, A_neg_shifted(18) => 
                           negative_inputs_23_18_port, A_neg_shifted(17) => 
                           negative_inputs_23_17_port, A_neg_shifted(16) => 
                           negative_inputs_23_16_port, A_neg_shifted(15) => 
                           negative_inputs_23_15_port, A_neg_shifted(14) => 
                           negative_inputs_23_14_port, A_neg_shifted(13) => 
                           negative_inputs_23_13_port, A_neg_shifted(12) => 
                           negative_inputs_23_12_port, A_neg_shifted(11) => 
                           negative_inputs_23_11_port, A_neg_shifted(10) => 
                           negative_inputs_23_10_port, A_neg_shifted(9) => 
                           negative_inputs_23_9_port, A_neg_shifted(8) => 
                           negative_inputs_23_8_port, A_neg_shifted(7) => 
                           negative_inputs_23_7_port, A_neg_shifted(6) => 
                           negative_inputs_23_6_port, A_neg_shifted(5) => 
                           negative_inputs_23_5_port, A_neg_shifted(4) => 
                           negative_inputs_23_4_port, A_neg_shifted(3) => 
                           negative_inputs_23_3_port, A_neg_shifted(2) => 
                           negative_inputs_23_2_port, A_neg_shifted(1) => 
                           negative_inputs_23_1_port, A_neg_shifted(0) => n9, 
                           Sel(2) => sel_11_2_port, Sel(1) => sel_11_1_port, 
                           Sel(0) => sel_11_0_port, Y(63) => 
                           MuxOutputs_11_63_port, Y(62) => 
                           MuxOutputs_11_62_port, Y(61) => 
                           MuxOutputs_11_61_port, Y(60) => 
                           MuxOutputs_11_60_port, Y(59) => 
                           MuxOutputs_11_59_port, Y(58) => 
                           MuxOutputs_11_58_port, Y(57) => 
                           MuxOutputs_11_57_port, Y(56) => 
                           MuxOutputs_11_56_port, Y(55) => 
                           MuxOutputs_11_55_port, Y(54) => 
                           MuxOutputs_11_54_port, Y(53) => 
                           MuxOutputs_11_53_port, Y(52) => 
                           MuxOutputs_11_52_port, Y(51) => 
                           MuxOutputs_11_51_port, Y(50) => 
                           MuxOutputs_11_50_port, Y(49) => 
                           MuxOutputs_11_49_port, Y(48) => 
                           MuxOutputs_11_48_port, Y(47) => 
                           MuxOutputs_11_47_port, Y(46) => 
                           MuxOutputs_11_46_port, Y(45) => 
                           MuxOutputs_11_45_port, Y(44) => 
                           MuxOutputs_11_44_port, Y(43) => 
                           MuxOutputs_11_43_port, Y(42) => 
                           MuxOutputs_11_42_port, Y(41) => 
                           MuxOutputs_11_41_port, Y(40) => 
                           MuxOutputs_11_40_port, Y(39) => 
                           MuxOutputs_11_39_port, Y(38) => 
                           MuxOutputs_11_38_port, Y(37) => 
                           MuxOutputs_11_37_port, Y(36) => 
                           MuxOutputs_11_36_port, Y(35) => 
                           MuxOutputs_11_35_port, Y(34) => 
                           MuxOutputs_11_34_port, Y(33) => 
                           MuxOutputs_11_33_port, Y(32) => 
                           MuxOutputs_11_32_port, Y(31) => 
                           MuxOutputs_11_31_port, Y(30) => 
                           MuxOutputs_11_30_port, Y(29) => 
                           MuxOutputs_11_29_port, Y(28) => 
                           MuxOutputs_11_28_port, Y(27) => 
                           MuxOutputs_11_27_port, Y(26) => 
                           MuxOutputs_11_26_port, Y(25) => 
                           MuxOutputs_11_25_port, Y(24) => 
                           MuxOutputs_11_24_port, Y(23) => 
                           MuxOutputs_11_23_port, Y(22) => 
                           MuxOutputs_11_22_port, Y(21) => 
                           MuxOutputs_11_21_port, Y(20) => 
                           MuxOutputs_11_20_port, Y(19) => 
                           MuxOutputs_11_19_port, Y(18) => 
                           MuxOutputs_11_18_port, Y(17) => 
                           MuxOutputs_11_17_port, Y(16) => 
                           MuxOutputs_11_16_port, Y(15) => 
                           MuxOutputs_11_15_port, Y(14) => 
                           MuxOutputs_11_14_port, Y(13) => 
                           MuxOutputs_11_13_port, Y(12) => 
                           MuxOutputs_11_12_port, Y(11) => 
                           MuxOutputs_11_11_port, Y(10) => 
                           MuxOutputs_11_10_port, Y(9) => MuxOutputs_11_9_port,
                           Y(8) => MuxOutputs_11_8_port, Y(7) => 
                           MuxOutputs_11_7_port, Y(6) => MuxOutputs_11_6_port, 
                           Y(5) => MuxOutputs_11_5_port, Y(4) => 
                           MuxOutputs_11_4_port, Y(3) => MuxOutputs_11_3_port, 
                           Y(2) => MuxOutputs_11_2_port, Y(1) => 
                           MuxOutputs_11_1_port, Y(0) => MuxOutputs_11_0_port);
   encoderI_12 : encoder_4 port map( pieceofB(2) => B(25), pieceofB(1) => B(24)
                           , pieceofB(0) => B(23), sel(2) => sel_12_2_port, 
                           sel(1) => sel_12_1_port, sel(0) => sel_12_0_port);
   MUXI_12 : MUX51_MuxNbit64_4 port map( zeroSignal(63) => X_Logic0_port, 
                           zeroSignal(62) => X_Logic0_port, zeroSignal(61) => 
                           X_Logic0_port, zeroSignal(60) => X_Logic0_port, 
                           zeroSignal(59) => X_Logic0_port, zeroSignal(58) => 
                           X_Logic0_port, zeroSignal(57) => X_Logic0_port, 
                           zeroSignal(56) => X_Logic0_port, zeroSignal(55) => 
                           X_Logic0_port, zeroSignal(54) => X_Logic0_port, 
                           zeroSignal(53) => X_Logic0_port, zeroSignal(52) => 
                           X_Logic0_port, zeroSignal(51) => X_Logic0_port, 
                           zeroSignal(50) => X_Logic0_port, zeroSignal(49) => 
                           X_Logic0_port, zeroSignal(48) => X_Logic0_port, 
                           zeroSignal(47) => X_Logic0_port, zeroSignal(46) => 
                           X_Logic0_port, zeroSignal(45) => X_Logic0_port, 
                           zeroSignal(44) => X_Logic0_port, zeroSignal(43) => 
                           X_Logic0_port, zeroSignal(42) => X_Logic0_port, 
                           zeroSignal(41) => X_Logic0_port, zeroSignal(40) => 
                           X_Logic0_port, zeroSignal(39) => X_Logic0_port, 
                           zeroSignal(38) => X_Logic0_port, zeroSignal(37) => 
                           X_Logic0_port, zeroSignal(36) => X_Logic0_port, 
                           zeroSignal(35) => X_Logic0_port, zeroSignal(34) => 
                           X_Logic0_port, zeroSignal(33) => X_Logic0_port, 
                           zeroSignal(32) => X_Logic0_port, zeroSignal(31) => 
                           X_Logic0_port, zeroSignal(30) => X_Logic0_port, 
                           zeroSignal(29) => X_Logic0_port, zeroSignal(28) => 
                           X_Logic0_port, zeroSignal(27) => X_Logic0_port, 
                           zeroSignal(26) => X_Logic0_port, zeroSignal(25) => 
                           X_Logic0_port, zeroSignal(24) => X_Logic0_port, 
                           zeroSignal(23) => X_Logic0_port, zeroSignal(22) => 
                           X_Logic0_port, zeroSignal(21) => X_Logic0_port, 
                           zeroSignal(20) => X_Logic0_port, zeroSignal(19) => 
                           X_Logic0_port, zeroSignal(18) => X_Logic0_port, 
                           zeroSignal(17) => X_Logic0_port, zeroSignal(16) => 
                           X_Logic0_port, zeroSignal(15) => X_Logic0_port, 
                           zeroSignal(14) => X_Logic0_port, zeroSignal(13) => 
                           X_Logic0_port, zeroSignal(12) => X_Logic0_port, 
                           zeroSignal(11) => X_Logic0_port, zeroSignal(10) => 
                           X_Logic0_port, zeroSignal(9) => X_Logic0_port, 
                           zeroSignal(8) => X_Logic0_port, zeroSignal(7) => 
                           X_Logic0_port, zeroSignal(6) => X_Logic0_port, 
                           zeroSignal(5) => X_Logic0_port, zeroSignal(4) => 
                           X_Logic0_port, zeroSignal(3) => X_Logic0_port, 
                           zeroSignal(2) => X_Logic0_port, zeroSignal(1) => 
                           X_Logic0_port, zeroSignal(0) => X_Logic0_port, 
                           A_signal(63) => positive_inputs_24_63_port, 
                           A_signal(62) => positive_inputs_24_62_port, 
                           A_signal(61) => positive_inputs_24_61_port, 
                           A_signal(60) => positive_inputs_24_60_port, 
                           A_signal(59) => positive_inputs_24_59_port, 
                           A_signal(58) => positive_inputs_24_58_port, 
                           A_signal(57) => positive_inputs_24_57_port, 
                           A_signal(56) => positive_inputs_24_56_port, 
                           A_signal(55) => positive_inputs_24_55_port, 
                           A_signal(54) => positive_inputs_24_54_port, 
                           A_signal(53) => positive_inputs_24_53_port, 
                           A_signal(52) => positive_inputs_24_52_port, 
                           A_signal(51) => positive_inputs_24_51_port, 
                           A_signal(50) => positive_inputs_24_50_port, 
                           A_signal(49) => positive_inputs_24_49_port, 
                           A_signal(48) => positive_inputs_24_48_port, 
                           A_signal(47) => positive_inputs_24_47_port, 
                           A_signal(46) => positive_inputs_24_46_port, 
                           A_signal(45) => positive_inputs_24_45_port, 
                           A_signal(44) => positive_inputs_24_44_port, 
                           A_signal(43) => positive_inputs_24_43_port, 
                           A_signal(42) => positive_inputs_24_42_port, 
                           A_signal(41) => positive_inputs_24_41_port, 
                           A_signal(40) => positive_inputs_24_40_port, 
                           A_signal(39) => positive_inputs_24_39_port, 
                           A_signal(38) => positive_inputs_24_38_port, 
                           A_signal(37) => positive_inputs_24_37_port, 
                           A_signal(36) => positive_inputs_24_36_port, 
                           A_signal(35) => positive_inputs_24_35_port, 
                           A_signal(34) => positive_inputs_24_34_port, 
                           A_signal(33) => positive_inputs_24_33_port, 
                           A_signal(32) => positive_inputs_24_32_port, 
                           A_signal(31) => positive_inputs_24_31_port, 
                           A_signal(30) => positive_inputs_24_30_port, 
                           A_signal(29) => positive_inputs_24_29_port, 
                           A_signal(28) => positive_inputs_24_28_port, 
                           A_signal(27) => positive_inputs_24_27_port, 
                           A_signal(26) => positive_inputs_24_26_port, 
                           A_signal(25) => positive_inputs_24_25_port, 
                           A_signal(24) => positive_inputs_24_24_port, 
                           A_signal(23) => positive_inputs_24_23_port, 
                           A_signal(22) => positive_inputs_24_22_port, 
                           A_signal(21) => positive_inputs_24_21_port, 
                           A_signal(20) => positive_inputs_24_20_port, 
                           A_signal(19) => positive_inputs_24_19_port, 
                           A_signal(18) => positive_inputs_24_18_port, 
                           A_signal(17) => positive_inputs_24_17_port, 
                           A_signal(16) => positive_inputs_24_16_port, 
                           A_signal(15) => positive_inputs_24_15_port, 
                           A_signal(14) => positive_inputs_24_14_port, 
                           A_signal(13) => positive_inputs_24_13_port, 
                           A_signal(12) => positive_inputs_24_12_port, 
                           A_signal(11) => positive_inputs_24_11_port, 
                           A_signal(10) => positive_inputs_24_10_port, 
                           A_signal(9) => positive_inputs_24_9_port, 
                           A_signal(8) => positive_inputs_24_8_port, 
                           A_signal(7) => positive_inputs_24_7_port, 
                           A_signal(6) => positive_inputs_24_6_port, 
                           A_signal(5) => positive_inputs_24_5_port, 
                           A_signal(4) => positive_inputs_24_4_port, 
                           A_signal(3) => positive_inputs_24_3_port, 
                           A_signal(2) => positive_inputs_24_2_port, 
                           A_signal(1) => positive_inputs_24_1_port, 
                           A_signal(0) => n9, A_neg(63) => 
                           negative_inputs_24_63_port, A_neg(62) => 
                           negative_inputs_24_62_port, A_neg(61) => 
                           negative_inputs_24_61_port, A_neg(60) => 
                           negative_inputs_24_60_port, A_neg(59) => 
                           negative_inputs_24_59_port, A_neg(58) => 
                           negative_inputs_24_58_port, A_neg(57) => 
                           negative_inputs_24_57_port, A_neg(56) => 
                           negative_inputs_24_56_port, A_neg(55) => 
                           negative_inputs_24_55_port, A_neg(54) => 
                           negative_inputs_24_54_port, A_neg(53) => 
                           negative_inputs_24_53_port, A_neg(52) => 
                           negative_inputs_24_52_port, A_neg(51) => 
                           negative_inputs_24_51_port, A_neg(50) => 
                           negative_inputs_24_50_port, A_neg(49) => 
                           negative_inputs_24_49_port, A_neg(48) => 
                           negative_inputs_24_48_port, A_neg(47) => 
                           negative_inputs_24_47_port, A_neg(46) => 
                           negative_inputs_24_46_port, A_neg(45) => 
                           negative_inputs_24_45_port, A_neg(44) => 
                           negative_inputs_24_44_port, A_neg(43) => 
                           negative_inputs_24_43_port, A_neg(42) => 
                           negative_inputs_24_42_port, A_neg(41) => 
                           negative_inputs_24_41_port, A_neg(40) => 
                           negative_inputs_24_40_port, A_neg(39) => 
                           negative_inputs_24_39_port, A_neg(38) => 
                           negative_inputs_24_38_port, A_neg(37) => 
                           negative_inputs_24_37_port, A_neg(36) => 
                           negative_inputs_24_36_port, A_neg(35) => 
                           negative_inputs_24_35_port, A_neg(34) => 
                           negative_inputs_24_34_port, A_neg(33) => 
                           negative_inputs_24_33_port, A_neg(32) => 
                           negative_inputs_24_32_port, A_neg(31) => 
                           negative_inputs_24_31_port, A_neg(30) => 
                           negative_inputs_24_30_port, A_neg(29) => 
                           negative_inputs_24_29_port, A_neg(28) => 
                           negative_inputs_24_28_port, A_neg(27) => 
                           negative_inputs_24_27_port, A_neg(26) => 
                           negative_inputs_24_26_port, A_neg(25) => 
                           negative_inputs_24_25_port, A_neg(24) => 
                           negative_inputs_24_24_port, A_neg(23) => 
                           negative_inputs_24_23_port, A_neg(22) => 
                           negative_inputs_24_22_port, A_neg(21) => 
                           negative_inputs_24_21_port, A_neg(20) => 
                           negative_inputs_24_20_port, A_neg(19) => 
                           negative_inputs_24_19_port, A_neg(18) => 
                           negative_inputs_24_18_port, A_neg(17) => 
                           negative_inputs_24_17_port, A_neg(16) => 
                           negative_inputs_24_16_port, A_neg(15) => 
                           negative_inputs_24_15_port, A_neg(14) => 
                           negative_inputs_24_14_port, A_neg(13) => 
                           negative_inputs_24_13_port, A_neg(12) => 
                           negative_inputs_24_12_port, A_neg(11) => 
                           negative_inputs_24_11_port, A_neg(10) => 
                           negative_inputs_24_10_port, A_neg(9) => 
                           negative_inputs_24_9_port, A_neg(8) => 
                           negative_inputs_24_8_port, A_neg(7) => 
                           negative_inputs_24_7_port, A_neg(6) => 
                           negative_inputs_24_6_port, A_neg(5) => 
                           negative_inputs_24_5_port, A_neg(4) => 
                           negative_inputs_24_4_port, A_neg(3) => 
                           negative_inputs_24_3_port, A_neg(2) => 
                           negative_inputs_24_2_port, A_neg(1) => 
                           negative_inputs_24_1_port, A_neg(0) => n9, 
                           A_shifted(63) => positive_inputs_25_63_port, 
                           A_shifted(62) => positive_inputs_25_62_port, 
                           A_shifted(61) => positive_inputs_25_61_port, 
                           A_shifted(60) => positive_inputs_25_60_port, 
                           A_shifted(59) => positive_inputs_25_59_port, 
                           A_shifted(58) => positive_inputs_25_58_port, 
                           A_shifted(57) => positive_inputs_25_57_port, 
                           A_shifted(56) => positive_inputs_25_56_port, 
                           A_shifted(55) => positive_inputs_25_55_port, 
                           A_shifted(54) => positive_inputs_25_54_port, 
                           A_shifted(53) => positive_inputs_25_53_port, 
                           A_shifted(52) => positive_inputs_25_52_port, 
                           A_shifted(51) => positive_inputs_25_51_port, 
                           A_shifted(50) => positive_inputs_25_50_port, 
                           A_shifted(49) => positive_inputs_25_49_port, 
                           A_shifted(48) => positive_inputs_25_48_port, 
                           A_shifted(47) => positive_inputs_25_47_port, 
                           A_shifted(46) => positive_inputs_25_46_port, 
                           A_shifted(45) => positive_inputs_25_45_port, 
                           A_shifted(44) => positive_inputs_25_44_port, 
                           A_shifted(43) => positive_inputs_25_43_port, 
                           A_shifted(42) => positive_inputs_25_42_port, 
                           A_shifted(41) => positive_inputs_25_41_port, 
                           A_shifted(40) => positive_inputs_25_40_port, 
                           A_shifted(39) => positive_inputs_25_39_port, 
                           A_shifted(38) => positive_inputs_25_38_port, 
                           A_shifted(37) => positive_inputs_25_37_port, 
                           A_shifted(36) => positive_inputs_25_36_port, 
                           A_shifted(35) => positive_inputs_25_35_port, 
                           A_shifted(34) => positive_inputs_25_34_port, 
                           A_shifted(33) => positive_inputs_25_33_port, 
                           A_shifted(32) => positive_inputs_25_32_port, 
                           A_shifted(31) => positive_inputs_25_31_port, 
                           A_shifted(30) => positive_inputs_25_30_port, 
                           A_shifted(29) => positive_inputs_25_29_port, 
                           A_shifted(28) => positive_inputs_25_28_port, 
                           A_shifted(27) => positive_inputs_25_27_port, 
                           A_shifted(26) => positive_inputs_25_26_port, 
                           A_shifted(25) => positive_inputs_25_25_port, 
                           A_shifted(24) => positive_inputs_25_24_port, 
                           A_shifted(23) => positive_inputs_25_23_port, 
                           A_shifted(22) => positive_inputs_25_22_port, 
                           A_shifted(21) => positive_inputs_25_21_port, 
                           A_shifted(20) => positive_inputs_25_20_port, 
                           A_shifted(19) => positive_inputs_25_19_port, 
                           A_shifted(18) => positive_inputs_25_18_port, 
                           A_shifted(17) => positive_inputs_25_17_port, 
                           A_shifted(16) => positive_inputs_25_16_port, 
                           A_shifted(15) => positive_inputs_25_15_port, 
                           A_shifted(14) => positive_inputs_25_14_port, 
                           A_shifted(13) => positive_inputs_25_13_port, 
                           A_shifted(12) => positive_inputs_25_12_port, 
                           A_shifted(11) => positive_inputs_25_11_port, 
                           A_shifted(10) => positive_inputs_25_10_port, 
                           A_shifted(9) => positive_inputs_25_9_port, 
                           A_shifted(8) => positive_inputs_25_8_port, 
                           A_shifted(7) => positive_inputs_25_7_port, 
                           A_shifted(6) => positive_inputs_25_6_port, 
                           A_shifted(5) => positive_inputs_25_5_port, 
                           A_shifted(4) => positive_inputs_25_4_port, 
                           A_shifted(3) => positive_inputs_25_3_port, 
                           A_shifted(2) => positive_inputs_25_2_port, 
                           A_shifted(1) => positive_inputs_25_1_port, 
                           A_shifted(0) => n9, A_neg_shifted(63) => 
                           negative_inputs_25_63_port, A_neg_shifted(62) => 
                           negative_inputs_25_62_port, A_neg_shifted(61) => 
                           negative_inputs_25_61_port, A_neg_shifted(60) => 
                           negative_inputs_25_60_port, A_neg_shifted(59) => 
                           negative_inputs_25_59_port, A_neg_shifted(58) => 
                           negative_inputs_25_58_port, A_neg_shifted(57) => 
                           negative_inputs_25_57_port, A_neg_shifted(56) => 
                           negative_inputs_25_56_port, A_neg_shifted(55) => 
                           negative_inputs_25_55_port, A_neg_shifted(54) => 
                           negative_inputs_25_54_port, A_neg_shifted(53) => 
                           negative_inputs_25_53_port, A_neg_shifted(52) => 
                           negative_inputs_25_52_port, A_neg_shifted(51) => 
                           negative_inputs_25_51_port, A_neg_shifted(50) => 
                           negative_inputs_25_50_port, A_neg_shifted(49) => 
                           negative_inputs_25_49_port, A_neg_shifted(48) => 
                           negative_inputs_25_48_port, A_neg_shifted(47) => 
                           negative_inputs_25_47_port, A_neg_shifted(46) => 
                           negative_inputs_25_46_port, A_neg_shifted(45) => 
                           negative_inputs_25_45_port, A_neg_shifted(44) => 
                           negative_inputs_25_44_port, A_neg_shifted(43) => 
                           negative_inputs_25_43_port, A_neg_shifted(42) => 
                           negative_inputs_25_42_port, A_neg_shifted(41) => 
                           negative_inputs_25_41_port, A_neg_shifted(40) => 
                           negative_inputs_25_40_port, A_neg_shifted(39) => 
                           negative_inputs_25_39_port, A_neg_shifted(38) => 
                           negative_inputs_25_38_port, A_neg_shifted(37) => 
                           negative_inputs_25_37_port, A_neg_shifted(36) => 
                           negative_inputs_25_36_port, A_neg_shifted(35) => 
                           negative_inputs_25_35_port, A_neg_shifted(34) => 
                           negative_inputs_25_34_port, A_neg_shifted(33) => 
                           negative_inputs_25_33_port, A_neg_shifted(32) => 
                           negative_inputs_25_32_port, A_neg_shifted(31) => 
                           negative_inputs_25_31_port, A_neg_shifted(30) => 
                           negative_inputs_25_30_port, A_neg_shifted(29) => 
                           negative_inputs_25_29_port, A_neg_shifted(28) => 
                           negative_inputs_25_28_port, A_neg_shifted(27) => 
                           negative_inputs_25_27_port, A_neg_shifted(26) => 
                           negative_inputs_25_26_port, A_neg_shifted(25) => 
                           negative_inputs_25_25_port, A_neg_shifted(24) => 
                           negative_inputs_25_24_port, A_neg_shifted(23) => 
                           negative_inputs_25_23_port, A_neg_shifted(22) => 
                           negative_inputs_25_22_port, A_neg_shifted(21) => 
                           negative_inputs_25_21_port, A_neg_shifted(20) => 
                           negative_inputs_25_20_port, A_neg_shifted(19) => 
                           negative_inputs_25_19_port, A_neg_shifted(18) => 
                           negative_inputs_25_18_port, A_neg_shifted(17) => 
                           negative_inputs_25_17_port, A_neg_shifted(16) => 
                           negative_inputs_25_16_port, A_neg_shifted(15) => 
                           negative_inputs_25_15_port, A_neg_shifted(14) => 
                           negative_inputs_25_14_port, A_neg_shifted(13) => 
                           negative_inputs_25_13_port, A_neg_shifted(12) => 
                           negative_inputs_25_12_port, A_neg_shifted(11) => 
                           negative_inputs_25_11_port, A_neg_shifted(10) => 
                           negative_inputs_25_10_port, A_neg_shifted(9) => 
                           negative_inputs_25_9_port, A_neg_shifted(8) => 
                           negative_inputs_25_8_port, A_neg_shifted(7) => 
                           negative_inputs_25_7_port, A_neg_shifted(6) => 
                           negative_inputs_25_6_port, A_neg_shifted(5) => 
                           negative_inputs_25_5_port, A_neg_shifted(4) => 
                           negative_inputs_25_4_port, A_neg_shifted(3) => 
                           negative_inputs_25_3_port, A_neg_shifted(2) => 
                           negative_inputs_25_2_port, A_neg_shifted(1) => 
                           negative_inputs_25_1_port, A_neg_shifted(0) => n9, 
                           Sel(2) => sel_12_2_port, Sel(1) => sel_12_1_port, 
                           Sel(0) => sel_12_0_port, Y(63) => 
                           MuxOutputs_12_63_port, Y(62) => 
                           MuxOutputs_12_62_port, Y(61) => 
                           MuxOutputs_12_61_port, Y(60) => 
                           MuxOutputs_12_60_port, Y(59) => 
                           MuxOutputs_12_59_port, Y(58) => 
                           MuxOutputs_12_58_port, Y(57) => 
                           MuxOutputs_12_57_port, Y(56) => 
                           MuxOutputs_12_56_port, Y(55) => 
                           MuxOutputs_12_55_port, Y(54) => 
                           MuxOutputs_12_54_port, Y(53) => 
                           MuxOutputs_12_53_port, Y(52) => 
                           MuxOutputs_12_52_port, Y(51) => 
                           MuxOutputs_12_51_port, Y(50) => 
                           MuxOutputs_12_50_port, Y(49) => 
                           MuxOutputs_12_49_port, Y(48) => 
                           MuxOutputs_12_48_port, Y(47) => 
                           MuxOutputs_12_47_port, Y(46) => 
                           MuxOutputs_12_46_port, Y(45) => 
                           MuxOutputs_12_45_port, Y(44) => 
                           MuxOutputs_12_44_port, Y(43) => 
                           MuxOutputs_12_43_port, Y(42) => 
                           MuxOutputs_12_42_port, Y(41) => 
                           MuxOutputs_12_41_port, Y(40) => 
                           MuxOutputs_12_40_port, Y(39) => 
                           MuxOutputs_12_39_port, Y(38) => 
                           MuxOutputs_12_38_port, Y(37) => 
                           MuxOutputs_12_37_port, Y(36) => 
                           MuxOutputs_12_36_port, Y(35) => 
                           MuxOutputs_12_35_port, Y(34) => 
                           MuxOutputs_12_34_port, Y(33) => 
                           MuxOutputs_12_33_port, Y(32) => 
                           MuxOutputs_12_32_port, Y(31) => 
                           MuxOutputs_12_31_port, Y(30) => 
                           MuxOutputs_12_30_port, Y(29) => 
                           MuxOutputs_12_29_port, Y(28) => 
                           MuxOutputs_12_28_port, Y(27) => 
                           MuxOutputs_12_27_port, Y(26) => 
                           MuxOutputs_12_26_port, Y(25) => 
                           MuxOutputs_12_25_port, Y(24) => 
                           MuxOutputs_12_24_port, Y(23) => 
                           MuxOutputs_12_23_port, Y(22) => 
                           MuxOutputs_12_22_port, Y(21) => 
                           MuxOutputs_12_21_port, Y(20) => 
                           MuxOutputs_12_20_port, Y(19) => 
                           MuxOutputs_12_19_port, Y(18) => 
                           MuxOutputs_12_18_port, Y(17) => 
                           MuxOutputs_12_17_port, Y(16) => 
                           MuxOutputs_12_16_port, Y(15) => 
                           MuxOutputs_12_15_port, Y(14) => 
                           MuxOutputs_12_14_port, Y(13) => 
                           MuxOutputs_12_13_port, Y(12) => 
                           MuxOutputs_12_12_port, Y(11) => 
                           MuxOutputs_12_11_port, Y(10) => 
                           MuxOutputs_12_10_port, Y(9) => MuxOutputs_12_9_port,
                           Y(8) => MuxOutputs_12_8_port, Y(7) => 
                           MuxOutputs_12_7_port, Y(6) => MuxOutputs_12_6_port, 
                           Y(5) => MuxOutputs_12_5_port, Y(4) => 
                           MuxOutputs_12_4_port, Y(3) => MuxOutputs_12_3_port, 
                           Y(2) => MuxOutputs_12_2_port, Y(1) => 
                           MuxOutputs_12_1_port, Y(0) => MuxOutputs_12_0_port);
   encoderI_13 : encoder_3 port map( pieceofB(2) => B(27), pieceofB(1) => B(26)
                           , pieceofB(0) => B(25), sel(2) => sel_13_2_port, 
                           sel(1) => sel_13_1_port, sel(0) => sel_13_0_port);
   MUXI_13 : MUX51_MuxNbit64_3 port map( zeroSignal(63) => X_Logic0_port, 
                           zeroSignal(62) => X_Logic0_port, zeroSignal(61) => 
                           X_Logic0_port, zeroSignal(60) => X_Logic0_port, 
                           zeroSignal(59) => X_Logic0_port, zeroSignal(58) => 
                           X_Logic0_port, zeroSignal(57) => X_Logic0_port, 
                           zeroSignal(56) => X_Logic0_port, zeroSignal(55) => 
                           X_Logic0_port, zeroSignal(54) => X_Logic0_port, 
                           zeroSignal(53) => X_Logic0_port, zeroSignal(52) => 
                           X_Logic0_port, zeroSignal(51) => X_Logic0_port, 
                           zeroSignal(50) => X_Logic0_port, zeroSignal(49) => 
                           X_Logic0_port, zeroSignal(48) => X_Logic0_port, 
                           zeroSignal(47) => X_Logic0_port, zeroSignal(46) => 
                           X_Logic0_port, zeroSignal(45) => X_Logic0_port, 
                           zeroSignal(44) => X_Logic0_port, zeroSignal(43) => 
                           X_Logic0_port, zeroSignal(42) => X_Logic0_port, 
                           zeroSignal(41) => X_Logic0_port, zeroSignal(40) => 
                           X_Logic0_port, zeroSignal(39) => X_Logic0_port, 
                           zeroSignal(38) => X_Logic0_port, zeroSignal(37) => 
                           X_Logic0_port, zeroSignal(36) => X_Logic0_port, 
                           zeroSignal(35) => X_Logic0_port, zeroSignal(34) => 
                           X_Logic0_port, zeroSignal(33) => X_Logic0_port, 
                           zeroSignal(32) => X_Logic0_port, zeroSignal(31) => 
                           X_Logic0_port, zeroSignal(30) => X_Logic0_port, 
                           zeroSignal(29) => X_Logic0_port, zeroSignal(28) => 
                           X_Logic0_port, zeroSignal(27) => X_Logic0_port, 
                           zeroSignal(26) => X_Logic0_port, zeroSignal(25) => 
                           X_Logic0_port, zeroSignal(24) => X_Logic0_port, 
                           zeroSignal(23) => X_Logic0_port, zeroSignal(22) => 
                           X_Logic0_port, zeroSignal(21) => X_Logic0_port, 
                           zeroSignal(20) => X_Logic0_port, zeroSignal(19) => 
                           X_Logic0_port, zeroSignal(18) => X_Logic0_port, 
                           zeroSignal(17) => X_Logic0_port, zeroSignal(16) => 
                           X_Logic0_port, zeroSignal(15) => X_Logic0_port, 
                           zeroSignal(14) => X_Logic0_port, zeroSignal(13) => 
                           X_Logic0_port, zeroSignal(12) => X_Logic0_port, 
                           zeroSignal(11) => X_Logic0_port, zeroSignal(10) => 
                           X_Logic0_port, zeroSignal(9) => X_Logic0_port, 
                           zeroSignal(8) => X_Logic0_port, zeroSignal(7) => 
                           X_Logic0_port, zeroSignal(6) => X_Logic0_port, 
                           zeroSignal(5) => X_Logic0_port, zeroSignal(4) => 
                           X_Logic0_port, zeroSignal(3) => X_Logic0_port, 
                           zeroSignal(2) => X_Logic0_port, zeroSignal(1) => 
                           X_Logic0_port, zeroSignal(0) => X_Logic0_port, 
                           A_signal(63) => positive_inputs_26_63_port, 
                           A_signal(62) => positive_inputs_26_62_port, 
                           A_signal(61) => positive_inputs_26_61_port, 
                           A_signal(60) => positive_inputs_26_60_port, 
                           A_signal(59) => positive_inputs_26_59_port, 
                           A_signal(58) => positive_inputs_26_58_port, 
                           A_signal(57) => positive_inputs_26_57_port, 
                           A_signal(56) => positive_inputs_26_56_port, 
                           A_signal(55) => positive_inputs_26_55_port, 
                           A_signal(54) => positive_inputs_26_54_port, 
                           A_signal(53) => positive_inputs_26_53_port, 
                           A_signal(52) => positive_inputs_26_52_port, 
                           A_signal(51) => positive_inputs_26_51_port, 
                           A_signal(50) => positive_inputs_26_50_port, 
                           A_signal(49) => positive_inputs_26_49_port, 
                           A_signal(48) => positive_inputs_26_48_port, 
                           A_signal(47) => positive_inputs_26_47_port, 
                           A_signal(46) => positive_inputs_26_46_port, 
                           A_signal(45) => positive_inputs_26_45_port, 
                           A_signal(44) => positive_inputs_26_44_port, 
                           A_signal(43) => positive_inputs_26_43_port, 
                           A_signal(42) => positive_inputs_26_42_port, 
                           A_signal(41) => positive_inputs_26_41_port, 
                           A_signal(40) => positive_inputs_26_40_port, 
                           A_signal(39) => positive_inputs_26_39_port, 
                           A_signal(38) => positive_inputs_26_38_port, 
                           A_signal(37) => positive_inputs_26_37_port, 
                           A_signal(36) => positive_inputs_26_36_port, 
                           A_signal(35) => positive_inputs_26_35_port, 
                           A_signal(34) => positive_inputs_26_34_port, 
                           A_signal(33) => positive_inputs_26_33_port, 
                           A_signal(32) => positive_inputs_26_32_port, 
                           A_signal(31) => positive_inputs_26_31_port, 
                           A_signal(30) => positive_inputs_26_30_port, 
                           A_signal(29) => positive_inputs_26_29_port, 
                           A_signal(28) => positive_inputs_26_28_port, 
                           A_signal(27) => positive_inputs_26_27_port, 
                           A_signal(26) => positive_inputs_26_26_port, 
                           A_signal(25) => positive_inputs_26_25_port, 
                           A_signal(24) => positive_inputs_26_24_port, 
                           A_signal(23) => positive_inputs_26_23_port, 
                           A_signal(22) => positive_inputs_26_22_port, 
                           A_signal(21) => positive_inputs_26_21_port, 
                           A_signal(20) => positive_inputs_26_20_port, 
                           A_signal(19) => positive_inputs_26_19_port, 
                           A_signal(18) => positive_inputs_26_18_port, 
                           A_signal(17) => positive_inputs_26_17_port, 
                           A_signal(16) => positive_inputs_26_16_port, 
                           A_signal(15) => positive_inputs_26_15_port, 
                           A_signal(14) => positive_inputs_26_14_port, 
                           A_signal(13) => positive_inputs_26_13_port, 
                           A_signal(12) => positive_inputs_26_12_port, 
                           A_signal(11) => positive_inputs_26_11_port, 
                           A_signal(10) => positive_inputs_26_10_port, 
                           A_signal(9) => positive_inputs_26_9_port, 
                           A_signal(8) => positive_inputs_26_8_port, 
                           A_signal(7) => positive_inputs_26_7_port, 
                           A_signal(6) => positive_inputs_26_6_port, 
                           A_signal(5) => positive_inputs_26_5_port, 
                           A_signal(4) => positive_inputs_26_4_port, 
                           A_signal(3) => positive_inputs_26_3_port, 
                           A_signal(2) => positive_inputs_26_2_port, 
                           A_signal(1) => positive_inputs_26_1_port, 
                           A_signal(0) => n9, A_neg(63) => 
                           negative_inputs_26_63_port, A_neg(62) => 
                           negative_inputs_26_62_port, A_neg(61) => 
                           negative_inputs_26_61_port, A_neg(60) => 
                           negative_inputs_26_60_port, A_neg(59) => 
                           negative_inputs_26_59_port, A_neg(58) => 
                           negative_inputs_26_58_port, A_neg(57) => 
                           negative_inputs_26_57_port, A_neg(56) => 
                           negative_inputs_26_56_port, A_neg(55) => 
                           negative_inputs_26_55_port, A_neg(54) => 
                           negative_inputs_26_54_port, A_neg(53) => 
                           negative_inputs_26_53_port, A_neg(52) => 
                           negative_inputs_26_52_port, A_neg(51) => 
                           negative_inputs_26_51_port, A_neg(50) => 
                           negative_inputs_26_50_port, A_neg(49) => 
                           negative_inputs_26_49_port, A_neg(48) => 
                           negative_inputs_26_48_port, A_neg(47) => 
                           negative_inputs_26_47_port, A_neg(46) => 
                           negative_inputs_26_46_port, A_neg(45) => 
                           negative_inputs_26_45_port, A_neg(44) => 
                           negative_inputs_26_44_port, A_neg(43) => 
                           negative_inputs_26_43_port, A_neg(42) => 
                           negative_inputs_26_42_port, A_neg(41) => 
                           negative_inputs_26_41_port, A_neg(40) => 
                           negative_inputs_26_40_port, A_neg(39) => 
                           negative_inputs_26_39_port, A_neg(38) => 
                           negative_inputs_26_38_port, A_neg(37) => 
                           negative_inputs_26_37_port, A_neg(36) => 
                           negative_inputs_26_36_port, A_neg(35) => 
                           negative_inputs_26_35_port, A_neg(34) => 
                           negative_inputs_26_34_port, A_neg(33) => 
                           negative_inputs_26_33_port, A_neg(32) => 
                           negative_inputs_26_32_port, A_neg(31) => 
                           negative_inputs_26_31_port, A_neg(30) => 
                           negative_inputs_26_30_port, A_neg(29) => 
                           negative_inputs_26_29_port, A_neg(28) => 
                           negative_inputs_26_28_port, A_neg(27) => 
                           negative_inputs_26_27_port, A_neg(26) => 
                           negative_inputs_26_26_port, A_neg(25) => 
                           negative_inputs_26_25_port, A_neg(24) => 
                           negative_inputs_26_24_port, A_neg(23) => 
                           negative_inputs_26_23_port, A_neg(22) => 
                           negative_inputs_26_22_port, A_neg(21) => 
                           negative_inputs_26_21_port, A_neg(20) => 
                           negative_inputs_26_20_port, A_neg(19) => 
                           negative_inputs_26_19_port, A_neg(18) => 
                           negative_inputs_26_18_port, A_neg(17) => 
                           negative_inputs_26_17_port, A_neg(16) => 
                           negative_inputs_26_16_port, A_neg(15) => 
                           negative_inputs_26_15_port, A_neg(14) => 
                           negative_inputs_26_14_port, A_neg(13) => 
                           negative_inputs_26_13_port, A_neg(12) => 
                           negative_inputs_26_12_port, A_neg(11) => 
                           negative_inputs_26_11_port, A_neg(10) => 
                           negative_inputs_26_10_port, A_neg(9) => 
                           negative_inputs_26_9_port, A_neg(8) => 
                           negative_inputs_26_8_port, A_neg(7) => 
                           negative_inputs_26_7_port, A_neg(6) => 
                           negative_inputs_26_6_port, A_neg(5) => 
                           negative_inputs_26_5_port, A_neg(4) => 
                           negative_inputs_26_4_port, A_neg(3) => 
                           negative_inputs_26_3_port, A_neg(2) => 
                           negative_inputs_26_2_port, A_neg(1) => 
                           negative_inputs_26_1_port, A_neg(0) => n9, 
                           A_shifted(63) => positive_inputs_27_63_port, 
                           A_shifted(62) => positive_inputs_27_62_port, 
                           A_shifted(61) => positive_inputs_27_61_port, 
                           A_shifted(60) => positive_inputs_27_60_port, 
                           A_shifted(59) => positive_inputs_27_59_port, 
                           A_shifted(58) => positive_inputs_27_58_port, 
                           A_shifted(57) => positive_inputs_27_57_port, 
                           A_shifted(56) => positive_inputs_27_56_port, 
                           A_shifted(55) => positive_inputs_27_55_port, 
                           A_shifted(54) => positive_inputs_27_54_port, 
                           A_shifted(53) => positive_inputs_27_53_port, 
                           A_shifted(52) => positive_inputs_27_52_port, 
                           A_shifted(51) => positive_inputs_27_51_port, 
                           A_shifted(50) => positive_inputs_27_50_port, 
                           A_shifted(49) => positive_inputs_27_49_port, 
                           A_shifted(48) => positive_inputs_27_48_port, 
                           A_shifted(47) => positive_inputs_27_47_port, 
                           A_shifted(46) => positive_inputs_27_46_port, 
                           A_shifted(45) => positive_inputs_27_45_port, 
                           A_shifted(44) => positive_inputs_27_44_port, 
                           A_shifted(43) => positive_inputs_27_43_port, 
                           A_shifted(42) => positive_inputs_27_42_port, 
                           A_shifted(41) => positive_inputs_27_41_port, 
                           A_shifted(40) => positive_inputs_27_40_port, 
                           A_shifted(39) => positive_inputs_27_39_port, 
                           A_shifted(38) => positive_inputs_27_38_port, 
                           A_shifted(37) => positive_inputs_27_37_port, 
                           A_shifted(36) => positive_inputs_27_36_port, 
                           A_shifted(35) => positive_inputs_27_35_port, 
                           A_shifted(34) => positive_inputs_27_34_port, 
                           A_shifted(33) => positive_inputs_27_33_port, 
                           A_shifted(32) => positive_inputs_27_32_port, 
                           A_shifted(31) => positive_inputs_27_31_port, 
                           A_shifted(30) => positive_inputs_27_30_port, 
                           A_shifted(29) => positive_inputs_27_29_port, 
                           A_shifted(28) => positive_inputs_27_28_port, 
                           A_shifted(27) => positive_inputs_27_27_port, 
                           A_shifted(26) => positive_inputs_27_26_port, 
                           A_shifted(25) => positive_inputs_27_25_port, 
                           A_shifted(24) => positive_inputs_27_24_port, 
                           A_shifted(23) => positive_inputs_27_23_port, 
                           A_shifted(22) => positive_inputs_27_22_port, 
                           A_shifted(21) => positive_inputs_27_21_port, 
                           A_shifted(20) => positive_inputs_27_20_port, 
                           A_shifted(19) => positive_inputs_27_19_port, 
                           A_shifted(18) => positive_inputs_27_18_port, 
                           A_shifted(17) => positive_inputs_27_17_port, 
                           A_shifted(16) => positive_inputs_27_16_port, 
                           A_shifted(15) => positive_inputs_27_15_port, 
                           A_shifted(14) => positive_inputs_27_14_port, 
                           A_shifted(13) => positive_inputs_27_13_port, 
                           A_shifted(12) => positive_inputs_27_12_port, 
                           A_shifted(11) => positive_inputs_27_11_port, 
                           A_shifted(10) => positive_inputs_27_10_port, 
                           A_shifted(9) => positive_inputs_27_9_port, 
                           A_shifted(8) => positive_inputs_27_8_port, 
                           A_shifted(7) => positive_inputs_27_7_port, 
                           A_shifted(6) => positive_inputs_27_6_port, 
                           A_shifted(5) => positive_inputs_27_5_port, 
                           A_shifted(4) => positive_inputs_27_4_port, 
                           A_shifted(3) => positive_inputs_27_3_port, 
                           A_shifted(2) => positive_inputs_27_2_port, 
                           A_shifted(1) => positive_inputs_27_1_port, 
                           A_shifted(0) => n9, A_neg_shifted(63) => 
                           negative_inputs_27_63_port, A_neg_shifted(62) => 
                           negative_inputs_27_62_port, A_neg_shifted(61) => 
                           negative_inputs_27_61_port, A_neg_shifted(60) => 
                           negative_inputs_27_60_port, A_neg_shifted(59) => 
                           negative_inputs_27_59_port, A_neg_shifted(58) => 
                           negative_inputs_27_58_port, A_neg_shifted(57) => 
                           negative_inputs_27_57_port, A_neg_shifted(56) => 
                           negative_inputs_27_56_port, A_neg_shifted(55) => 
                           negative_inputs_27_55_port, A_neg_shifted(54) => 
                           negative_inputs_27_54_port, A_neg_shifted(53) => 
                           negative_inputs_27_53_port, A_neg_shifted(52) => 
                           negative_inputs_27_52_port, A_neg_shifted(51) => 
                           negative_inputs_27_51_port, A_neg_shifted(50) => 
                           negative_inputs_27_50_port, A_neg_shifted(49) => 
                           negative_inputs_27_49_port, A_neg_shifted(48) => 
                           negative_inputs_27_48_port, A_neg_shifted(47) => 
                           negative_inputs_27_47_port, A_neg_shifted(46) => 
                           negative_inputs_27_46_port, A_neg_shifted(45) => 
                           negative_inputs_27_45_port, A_neg_shifted(44) => 
                           negative_inputs_27_44_port, A_neg_shifted(43) => 
                           negative_inputs_27_43_port, A_neg_shifted(42) => 
                           negative_inputs_27_42_port, A_neg_shifted(41) => 
                           negative_inputs_27_41_port, A_neg_shifted(40) => 
                           negative_inputs_27_40_port, A_neg_shifted(39) => 
                           negative_inputs_27_39_port, A_neg_shifted(38) => 
                           negative_inputs_27_38_port, A_neg_shifted(37) => 
                           negative_inputs_27_37_port, A_neg_shifted(36) => 
                           negative_inputs_27_36_port, A_neg_shifted(35) => 
                           negative_inputs_27_35_port, A_neg_shifted(34) => 
                           negative_inputs_27_34_port, A_neg_shifted(33) => 
                           negative_inputs_27_33_port, A_neg_shifted(32) => 
                           negative_inputs_27_32_port, A_neg_shifted(31) => 
                           negative_inputs_27_31_port, A_neg_shifted(30) => 
                           negative_inputs_27_30_port, A_neg_shifted(29) => 
                           negative_inputs_27_29_port, A_neg_shifted(28) => 
                           negative_inputs_27_28_port, A_neg_shifted(27) => 
                           negative_inputs_27_27_port, A_neg_shifted(26) => 
                           negative_inputs_27_26_port, A_neg_shifted(25) => 
                           negative_inputs_27_25_port, A_neg_shifted(24) => 
                           negative_inputs_27_24_port, A_neg_shifted(23) => 
                           negative_inputs_27_23_port, A_neg_shifted(22) => 
                           negative_inputs_27_22_port, A_neg_shifted(21) => 
                           negative_inputs_27_21_port, A_neg_shifted(20) => 
                           negative_inputs_27_20_port, A_neg_shifted(19) => 
                           negative_inputs_27_19_port, A_neg_shifted(18) => 
                           negative_inputs_27_18_port, A_neg_shifted(17) => 
                           negative_inputs_27_17_port, A_neg_shifted(16) => 
                           negative_inputs_27_16_port, A_neg_shifted(15) => 
                           negative_inputs_27_15_port, A_neg_shifted(14) => 
                           negative_inputs_27_14_port, A_neg_shifted(13) => 
                           negative_inputs_27_13_port, A_neg_shifted(12) => 
                           negative_inputs_27_12_port, A_neg_shifted(11) => 
                           negative_inputs_27_11_port, A_neg_shifted(10) => 
                           negative_inputs_27_10_port, A_neg_shifted(9) => 
                           negative_inputs_27_9_port, A_neg_shifted(8) => 
                           negative_inputs_27_8_port, A_neg_shifted(7) => 
                           negative_inputs_27_7_port, A_neg_shifted(6) => 
                           negative_inputs_27_6_port, A_neg_shifted(5) => 
                           negative_inputs_27_5_port, A_neg_shifted(4) => 
                           negative_inputs_27_4_port, A_neg_shifted(3) => 
                           negative_inputs_27_3_port, A_neg_shifted(2) => 
                           negative_inputs_27_2_port, A_neg_shifted(1) => 
                           negative_inputs_27_1_port, A_neg_shifted(0) => n9, 
                           Sel(2) => sel_13_2_port, Sel(1) => sel_13_1_port, 
                           Sel(0) => sel_13_0_port, Y(63) => 
                           MuxOutputs_13_63_port, Y(62) => 
                           MuxOutputs_13_62_port, Y(61) => 
                           MuxOutputs_13_61_port, Y(60) => 
                           MuxOutputs_13_60_port, Y(59) => 
                           MuxOutputs_13_59_port, Y(58) => 
                           MuxOutputs_13_58_port, Y(57) => 
                           MuxOutputs_13_57_port, Y(56) => 
                           MuxOutputs_13_56_port, Y(55) => 
                           MuxOutputs_13_55_port, Y(54) => 
                           MuxOutputs_13_54_port, Y(53) => 
                           MuxOutputs_13_53_port, Y(52) => 
                           MuxOutputs_13_52_port, Y(51) => 
                           MuxOutputs_13_51_port, Y(50) => 
                           MuxOutputs_13_50_port, Y(49) => 
                           MuxOutputs_13_49_port, Y(48) => 
                           MuxOutputs_13_48_port, Y(47) => 
                           MuxOutputs_13_47_port, Y(46) => 
                           MuxOutputs_13_46_port, Y(45) => 
                           MuxOutputs_13_45_port, Y(44) => 
                           MuxOutputs_13_44_port, Y(43) => 
                           MuxOutputs_13_43_port, Y(42) => 
                           MuxOutputs_13_42_port, Y(41) => 
                           MuxOutputs_13_41_port, Y(40) => 
                           MuxOutputs_13_40_port, Y(39) => 
                           MuxOutputs_13_39_port, Y(38) => 
                           MuxOutputs_13_38_port, Y(37) => 
                           MuxOutputs_13_37_port, Y(36) => 
                           MuxOutputs_13_36_port, Y(35) => 
                           MuxOutputs_13_35_port, Y(34) => 
                           MuxOutputs_13_34_port, Y(33) => 
                           MuxOutputs_13_33_port, Y(32) => 
                           MuxOutputs_13_32_port, Y(31) => 
                           MuxOutputs_13_31_port, Y(30) => 
                           MuxOutputs_13_30_port, Y(29) => 
                           MuxOutputs_13_29_port, Y(28) => 
                           MuxOutputs_13_28_port, Y(27) => 
                           MuxOutputs_13_27_port, Y(26) => 
                           MuxOutputs_13_26_port, Y(25) => 
                           MuxOutputs_13_25_port, Y(24) => 
                           MuxOutputs_13_24_port, Y(23) => 
                           MuxOutputs_13_23_port, Y(22) => 
                           MuxOutputs_13_22_port, Y(21) => 
                           MuxOutputs_13_21_port, Y(20) => 
                           MuxOutputs_13_20_port, Y(19) => 
                           MuxOutputs_13_19_port, Y(18) => 
                           MuxOutputs_13_18_port, Y(17) => 
                           MuxOutputs_13_17_port, Y(16) => 
                           MuxOutputs_13_16_port, Y(15) => 
                           MuxOutputs_13_15_port, Y(14) => 
                           MuxOutputs_13_14_port, Y(13) => 
                           MuxOutputs_13_13_port, Y(12) => 
                           MuxOutputs_13_12_port, Y(11) => 
                           MuxOutputs_13_11_port, Y(10) => 
                           MuxOutputs_13_10_port, Y(9) => MuxOutputs_13_9_port,
                           Y(8) => MuxOutputs_13_8_port, Y(7) => 
                           MuxOutputs_13_7_port, Y(6) => MuxOutputs_13_6_port, 
                           Y(5) => MuxOutputs_13_5_port, Y(4) => 
                           MuxOutputs_13_4_port, Y(3) => MuxOutputs_13_3_port, 
                           Y(2) => MuxOutputs_13_2_port, Y(1) => 
                           MuxOutputs_13_1_port, Y(0) => MuxOutputs_13_0_port);
   encoderI_14 : encoder_2 port map( pieceofB(2) => B(29), pieceofB(1) => B(28)
                           , pieceofB(0) => B(27), sel(2) => sel_14_2_port, 
                           sel(1) => sel_14_1_port, sel(0) => sel_14_0_port);
   MUXI_14 : MUX51_MuxNbit64_2 port map( zeroSignal(63) => X_Logic0_port, 
                           zeroSignal(62) => X_Logic0_port, zeroSignal(61) => 
                           X_Logic0_port, zeroSignal(60) => X_Logic0_port, 
                           zeroSignal(59) => X_Logic0_port, zeroSignal(58) => 
                           X_Logic0_port, zeroSignal(57) => X_Logic0_port, 
                           zeroSignal(56) => X_Logic0_port, zeroSignal(55) => 
                           X_Logic0_port, zeroSignal(54) => X_Logic0_port, 
                           zeroSignal(53) => X_Logic0_port, zeroSignal(52) => 
                           X_Logic0_port, zeroSignal(51) => X_Logic0_port, 
                           zeroSignal(50) => X_Logic0_port, zeroSignal(49) => 
                           X_Logic0_port, zeroSignal(48) => X_Logic0_port, 
                           zeroSignal(47) => X_Logic0_port, zeroSignal(46) => 
                           X_Logic0_port, zeroSignal(45) => X_Logic0_port, 
                           zeroSignal(44) => X_Logic0_port, zeroSignal(43) => 
                           X_Logic0_port, zeroSignal(42) => X_Logic0_port, 
                           zeroSignal(41) => X_Logic0_port, zeroSignal(40) => 
                           X_Logic0_port, zeroSignal(39) => X_Logic0_port, 
                           zeroSignal(38) => X_Logic0_port, zeroSignal(37) => 
                           X_Logic0_port, zeroSignal(36) => X_Logic0_port, 
                           zeroSignal(35) => X_Logic0_port, zeroSignal(34) => 
                           X_Logic0_port, zeroSignal(33) => X_Logic0_port, 
                           zeroSignal(32) => X_Logic0_port, zeroSignal(31) => 
                           X_Logic0_port, zeroSignal(30) => X_Logic0_port, 
                           zeroSignal(29) => X_Logic0_port, zeroSignal(28) => 
                           X_Logic0_port, zeroSignal(27) => X_Logic0_port, 
                           zeroSignal(26) => X_Logic0_port, zeroSignal(25) => 
                           X_Logic0_port, zeroSignal(24) => X_Logic0_port, 
                           zeroSignal(23) => X_Logic0_port, zeroSignal(22) => 
                           X_Logic0_port, zeroSignal(21) => X_Logic0_port, 
                           zeroSignal(20) => X_Logic0_port, zeroSignal(19) => 
                           X_Logic0_port, zeroSignal(18) => X_Logic0_port, 
                           zeroSignal(17) => X_Logic0_port, zeroSignal(16) => 
                           X_Logic0_port, zeroSignal(15) => X_Logic0_port, 
                           zeroSignal(14) => X_Logic0_port, zeroSignal(13) => 
                           X_Logic0_port, zeroSignal(12) => X_Logic0_port, 
                           zeroSignal(11) => X_Logic0_port, zeroSignal(10) => 
                           X_Logic0_port, zeroSignal(9) => X_Logic0_port, 
                           zeroSignal(8) => X_Logic0_port, zeroSignal(7) => 
                           X_Logic0_port, zeroSignal(6) => X_Logic0_port, 
                           zeroSignal(5) => X_Logic0_port, zeroSignal(4) => 
                           X_Logic0_port, zeroSignal(3) => X_Logic0_port, 
                           zeroSignal(2) => X_Logic0_port, zeroSignal(1) => 
                           X_Logic0_port, zeroSignal(0) => X_Logic0_port, 
                           A_signal(63) => positive_inputs_28_63_port, 
                           A_signal(62) => positive_inputs_28_62_port, 
                           A_signal(61) => positive_inputs_28_61_port, 
                           A_signal(60) => positive_inputs_28_60_port, 
                           A_signal(59) => positive_inputs_28_59_port, 
                           A_signal(58) => positive_inputs_28_58_port, 
                           A_signal(57) => positive_inputs_28_57_port, 
                           A_signal(56) => positive_inputs_28_56_port, 
                           A_signal(55) => positive_inputs_28_55_port, 
                           A_signal(54) => positive_inputs_28_54_port, 
                           A_signal(53) => positive_inputs_28_53_port, 
                           A_signal(52) => positive_inputs_28_52_port, 
                           A_signal(51) => positive_inputs_28_51_port, 
                           A_signal(50) => positive_inputs_28_50_port, 
                           A_signal(49) => positive_inputs_28_49_port, 
                           A_signal(48) => positive_inputs_28_48_port, 
                           A_signal(47) => positive_inputs_28_47_port, 
                           A_signal(46) => positive_inputs_28_46_port, 
                           A_signal(45) => positive_inputs_28_45_port, 
                           A_signal(44) => positive_inputs_28_44_port, 
                           A_signal(43) => positive_inputs_28_43_port, 
                           A_signal(42) => positive_inputs_28_42_port, 
                           A_signal(41) => positive_inputs_28_41_port, 
                           A_signal(40) => positive_inputs_28_40_port, 
                           A_signal(39) => positive_inputs_28_39_port, 
                           A_signal(38) => positive_inputs_28_38_port, 
                           A_signal(37) => positive_inputs_28_37_port, 
                           A_signal(36) => positive_inputs_28_36_port, 
                           A_signal(35) => positive_inputs_28_35_port, 
                           A_signal(34) => positive_inputs_28_34_port, 
                           A_signal(33) => positive_inputs_28_33_port, 
                           A_signal(32) => positive_inputs_28_32_port, 
                           A_signal(31) => positive_inputs_28_31_port, 
                           A_signal(30) => positive_inputs_28_30_port, 
                           A_signal(29) => positive_inputs_28_29_port, 
                           A_signal(28) => positive_inputs_28_28_port, 
                           A_signal(27) => positive_inputs_28_27_port, 
                           A_signal(26) => positive_inputs_28_26_port, 
                           A_signal(25) => positive_inputs_28_25_port, 
                           A_signal(24) => positive_inputs_28_24_port, 
                           A_signal(23) => positive_inputs_28_23_port, 
                           A_signal(22) => positive_inputs_28_22_port, 
                           A_signal(21) => positive_inputs_28_21_port, 
                           A_signal(20) => positive_inputs_28_20_port, 
                           A_signal(19) => positive_inputs_28_19_port, 
                           A_signal(18) => positive_inputs_28_18_port, 
                           A_signal(17) => positive_inputs_28_17_port, 
                           A_signal(16) => positive_inputs_28_16_port, 
                           A_signal(15) => positive_inputs_28_15_port, 
                           A_signal(14) => positive_inputs_28_14_port, 
                           A_signal(13) => positive_inputs_28_13_port, 
                           A_signal(12) => positive_inputs_28_12_port, 
                           A_signal(11) => positive_inputs_28_11_port, 
                           A_signal(10) => positive_inputs_28_10_port, 
                           A_signal(9) => positive_inputs_28_9_port, 
                           A_signal(8) => positive_inputs_28_8_port, 
                           A_signal(7) => positive_inputs_28_7_port, 
                           A_signal(6) => positive_inputs_28_6_port, 
                           A_signal(5) => positive_inputs_28_5_port, 
                           A_signal(4) => positive_inputs_28_4_port, 
                           A_signal(3) => positive_inputs_28_3_port, 
                           A_signal(2) => positive_inputs_28_2_port, 
                           A_signal(1) => positive_inputs_28_1_port, 
                           A_signal(0) => n9, A_neg(63) => 
                           negative_inputs_28_63_port, A_neg(62) => 
                           negative_inputs_28_62_port, A_neg(61) => 
                           negative_inputs_28_61_port, A_neg(60) => 
                           negative_inputs_28_60_port, A_neg(59) => 
                           negative_inputs_28_59_port, A_neg(58) => 
                           negative_inputs_28_58_port, A_neg(57) => 
                           negative_inputs_28_57_port, A_neg(56) => 
                           negative_inputs_28_56_port, A_neg(55) => 
                           negative_inputs_28_55_port, A_neg(54) => 
                           negative_inputs_28_54_port, A_neg(53) => 
                           negative_inputs_28_53_port, A_neg(52) => 
                           negative_inputs_28_52_port, A_neg(51) => 
                           negative_inputs_28_51_port, A_neg(50) => 
                           negative_inputs_28_50_port, A_neg(49) => 
                           negative_inputs_28_49_port, A_neg(48) => 
                           negative_inputs_28_48_port, A_neg(47) => 
                           negative_inputs_28_47_port, A_neg(46) => 
                           negative_inputs_28_46_port, A_neg(45) => 
                           negative_inputs_28_45_port, A_neg(44) => 
                           negative_inputs_28_44_port, A_neg(43) => 
                           negative_inputs_28_43_port, A_neg(42) => 
                           negative_inputs_28_42_port, A_neg(41) => 
                           negative_inputs_28_41_port, A_neg(40) => 
                           negative_inputs_28_40_port, A_neg(39) => 
                           negative_inputs_28_39_port, A_neg(38) => 
                           negative_inputs_28_38_port, A_neg(37) => 
                           negative_inputs_28_37_port, A_neg(36) => 
                           negative_inputs_28_36_port, A_neg(35) => 
                           negative_inputs_28_35_port, A_neg(34) => 
                           negative_inputs_28_34_port, A_neg(33) => 
                           negative_inputs_28_33_port, A_neg(32) => 
                           negative_inputs_28_32_port, A_neg(31) => 
                           negative_inputs_28_31_port, A_neg(30) => 
                           negative_inputs_28_30_port, A_neg(29) => 
                           negative_inputs_28_29_port, A_neg(28) => 
                           negative_inputs_28_28_port, A_neg(27) => 
                           negative_inputs_28_27_port, A_neg(26) => 
                           negative_inputs_28_26_port, A_neg(25) => 
                           negative_inputs_28_25_port, A_neg(24) => 
                           negative_inputs_28_24_port, A_neg(23) => 
                           negative_inputs_28_23_port, A_neg(22) => 
                           negative_inputs_28_22_port, A_neg(21) => 
                           negative_inputs_28_21_port, A_neg(20) => 
                           negative_inputs_28_20_port, A_neg(19) => 
                           negative_inputs_28_19_port, A_neg(18) => 
                           negative_inputs_28_18_port, A_neg(17) => 
                           negative_inputs_28_17_port, A_neg(16) => 
                           negative_inputs_28_16_port, A_neg(15) => 
                           negative_inputs_28_15_port, A_neg(14) => 
                           negative_inputs_28_14_port, A_neg(13) => 
                           negative_inputs_28_13_port, A_neg(12) => 
                           negative_inputs_28_12_port, A_neg(11) => 
                           negative_inputs_28_11_port, A_neg(10) => 
                           negative_inputs_28_10_port, A_neg(9) => 
                           negative_inputs_28_9_port, A_neg(8) => 
                           negative_inputs_28_8_port, A_neg(7) => 
                           negative_inputs_28_7_port, A_neg(6) => 
                           negative_inputs_28_6_port, A_neg(5) => 
                           negative_inputs_28_5_port, A_neg(4) => 
                           negative_inputs_28_4_port, A_neg(3) => 
                           negative_inputs_28_3_port, A_neg(2) => 
                           negative_inputs_28_2_port, A_neg(1) => 
                           negative_inputs_28_1_port, A_neg(0) => n9, 
                           A_shifted(63) => positive_inputs_29_63_port, 
                           A_shifted(62) => positive_inputs_29_62_port, 
                           A_shifted(61) => positive_inputs_29_61_port, 
                           A_shifted(60) => positive_inputs_29_60_port, 
                           A_shifted(59) => positive_inputs_29_59_port, 
                           A_shifted(58) => positive_inputs_29_58_port, 
                           A_shifted(57) => positive_inputs_29_57_port, 
                           A_shifted(56) => positive_inputs_29_56_port, 
                           A_shifted(55) => positive_inputs_29_55_port, 
                           A_shifted(54) => positive_inputs_29_54_port, 
                           A_shifted(53) => positive_inputs_29_53_port, 
                           A_shifted(52) => positive_inputs_29_52_port, 
                           A_shifted(51) => positive_inputs_29_51_port, 
                           A_shifted(50) => positive_inputs_29_50_port, 
                           A_shifted(49) => positive_inputs_29_49_port, 
                           A_shifted(48) => positive_inputs_29_48_port, 
                           A_shifted(47) => positive_inputs_29_47_port, 
                           A_shifted(46) => positive_inputs_29_46_port, 
                           A_shifted(45) => positive_inputs_29_45_port, 
                           A_shifted(44) => positive_inputs_29_44_port, 
                           A_shifted(43) => positive_inputs_29_43_port, 
                           A_shifted(42) => positive_inputs_29_42_port, 
                           A_shifted(41) => positive_inputs_29_41_port, 
                           A_shifted(40) => positive_inputs_29_40_port, 
                           A_shifted(39) => positive_inputs_29_39_port, 
                           A_shifted(38) => positive_inputs_29_38_port, 
                           A_shifted(37) => positive_inputs_29_37_port, 
                           A_shifted(36) => positive_inputs_29_36_port, 
                           A_shifted(35) => positive_inputs_29_35_port, 
                           A_shifted(34) => positive_inputs_29_34_port, 
                           A_shifted(33) => positive_inputs_29_33_port, 
                           A_shifted(32) => positive_inputs_29_32_port, 
                           A_shifted(31) => positive_inputs_29_31_port, 
                           A_shifted(30) => positive_inputs_29_30_port, 
                           A_shifted(29) => positive_inputs_29_29_port, 
                           A_shifted(28) => positive_inputs_29_28_port, 
                           A_shifted(27) => positive_inputs_29_27_port, 
                           A_shifted(26) => positive_inputs_29_26_port, 
                           A_shifted(25) => positive_inputs_29_25_port, 
                           A_shifted(24) => positive_inputs_29_24_port, 
                           A_shifted(23) => positive_inputs_29_23_port, 
                           A_shifted(22) => positive_inputs_29_22_port, 
                           A_shifted(21) => positive_inputs_29_21_port, 
                           A_shifted(20) => positive_inputs_29_20_port, 
                           A_shifted(19) => positive_inputs_29_19_port, 
                           A_shifted(18) => positive_inputs_29_18_port, 
                           A_shifted(17) => positive_inputs_29_17_port, 
                           A_shifted(16) => positive_inputs_29_16_port, 
                           A_shifted(15) => positive_inputs_29_15_port, 
                           A_shifted(14) => positive_inputs_29_14_port, 
                           A_shifted(13) => positive_inputs_29_13_port, 
                           A_shifted(12) => positive_inputs_29_12_port, 
                           A_shifted(11) => positive_inputs_29_11_port, 
                           A_shifted(10) => positive_inputs_29_10_port, 
                           A_shifted(9) => positive_inputs_29_9_port, 
                           A_shifted(8) => positive_inputs_29_8_port, 
                           A_shifted(7) => positive_inputs_29_7_port, 
                           A_shifted(6) => positive_inputs_29_6_port, 
                           A_shifted(5) => positive_inputs_29_5_port, 
                           A_shifted(4) => positive_inputs_29_4_port, 
                           A_shifted(3) => positive_inputs_29_3_port, 
                           A_shifted(2) => positive_inputs_29_2_port, 
                           A_shifted(1) => positive_inputs_29_1_port, 
                           A_shifted(0) => n9, A_neg_shifted(63) => 
                           negative_inputs_29_63_port, A_neg_shifted(62) => 
                           negative_inputs_29_62_port, A_neg_shifted(61) => 
                           negative_inputs_29_61_port, A_neg_shifted(60) => 
                           negative_inputs_29_60_port, A_neg_shifted(59) => 
                           negative_inputs_29_59_port, A_neg_shifted(58) => 
                           negative_inputs_29_58_port, A_neg_shifted(57) => 
                           negative_inputs_29_57_port, A_neg_shifted(56) => 
                           negative_inputs_29_56_port, A_neg_shifted(55) => 
                           negative_inputs_29_55_port, A_neg_shifted(54) => 
                           negative_inputs_29_54_port, A_neg_shifted(53) => 
                           negative_inputs_29_53_port, A_neg_shifted(52) => 
                           negative_inputs_29_52_port, A_neg_shifted(51) => 
                           negative_inputs_29_51_port, A_neg_shifted(50) => 
                           negative_inputs_29_50_port, A_neg_shifted(49) => 
                           negative_inputs_29_49_port, A_neg_shifted(48) => 
                           negative_inputs_29_48_port, A_neg_shifted(47) => 
                           negative_inputs_29_47_port, A_neg_shifted(46) => 
                           negative_inputs_29_46_port, A_neg_shifted(45) => 
                           negative_inputs_29_45_port, A_neg_shifted(44) => 
                           negative_inputs_29_44_port, A_neg_shifted(43) => 
                           negative_inputs_29_43_port, A_neg_shifted(42) => 
                           negative_inputs_29_42_port, A_neg_shifted(41) => 
                           negative_inputs_29_41_port, A_neg_shifted(40) => 
                           negative_inputs_29_40_port, A_neg_shifted(39) => 
                           negative_inputs_29_39_port, A_neg_shifted(38) => 
                           negative_inputs_29_38_port, A_neg_shifted(37) => 
                           negative_inputs_29_37_port, A_neg_shifted(36) => 
                           negative_inputs_29_36_port, A_neg_shifted(35) => 
                           negative_inputs_29_35_port, A_neg_shifted(34) => 
                           negative_inputs_29_34_port, A_neg_shifted(33) => 
                           negative_inputs_29_33_port, A_neg_shifted(32) => 
                           negative_inputs_29_32_port, A_neg_shifted(31) => 
                           negative_inputs_29_31_port, A_neg_shifted(30) => 
                           negative_inputs_29_30_port, A_neg_shifted(29) => 
                           negative_inputs_29_29_port, A_neg_shifted(28) => 
                           negative_inputs_29_28_port, A_neg_shifted(27) => 
                           negative_inputs_29_27_port, A_neg_shifted(26) => 
                           negative_inputs_29_26_port, A_neg_shifted(25) => 
                           negative_inputs_29_25_port, A_neg_shifted(24) => 
                           negative_inputs_29_24_port, A_neg_shifted(23) => 
                           negative_inputs_29_23_port, A_neg_shifted(22) => 
                           negative_inputs_29_22_port, A_neg_shifted(21) => 
                           negative_inputs_29_21_port, A_neg_shifted(20) => 
                           negative_inputs_29_20_port, A_neg_shifted(19) => 
                           negative_inputs_29_19_port, A_neg_shifted(18) => 
                           negative_inputs_29_18_port, A_neg_shifted(17) => 
                           negative_inputs_29_17_port, A_neg_shifted(16) => 
                           negative_inputs_29_16_port, A_neg_shifted(15) => 
                           negative_inputs_29_15_port, A_neg_shifted(14) => 
                           negative_inputs_29_14_port, A_neg_shifted(13) => 
                           negative_inputs_29_13_port, A_neg_shifted(12) => 
                           negative_inputs_29_12_port, A_neg_shifted(11) => 
                           negative_inputs_29_11_port, A_neg_shifted(10) => 
                           negative_inputs_29_10_port, A_neg_shifted(9) => 
                           negative_inputs_29_9_port, A_neg_shifted(8) => 
                           negative_inputs_29_8_port, A_neg_shifted(7) => 
                           negative_inputs_29_7_port, A_neg_shifted(6) => 
                           negative_inputs_29_6_port, A_neg_shifted(5) => 
                           negative_inputs_29_5_port, A_neg_shifted(4) => 
                           negative_inputs_29_4_port, A_neg_shifted(3) => 
                           negative_inputs_29_3_port, A_neg_shifted(2) => 
                           negative_inputs_29_2_port, A_neg_shifted(1) => 
                           negative_inputs_29_1_port, A_neg_shifted(0) => n9, 
                           Sel(2) => sel_14_2_port, Sel(1) => sel_14_1_port, 
                           Sel(0) => sel_14_0_port, Y(63) => 
                           MuxOutputs_14_63_port, Y(62) => 
                           MuxOutputs_14_62_port, Y(61) => 
                           MuxOutputs_14_61_port, Y(60) => 
                           MuxOutputs_14_60_port, Y(59) => 
                           MuxOutputs_14_59_port, Y(58) => 
                           MuxOutputs_14_58_port, Y(57) => 
                           MuxOutputs_14_57_port, Y(56) => 
                           MuxOutputs_14_56_port, Y(55) => 
                           MuxOutputs_14_55_port, Y(54) => 
                           MuxOutputs_14_54_port, Y(53) => 
                           MuxOutputs_14_53_port, Y(52) => 
                           MuxOutputs_14_52_port, Y(51) => 
                           MuxOutputs_14_51_port, Y(50) => 
                           MuxOutputs_14_50_port, Y(49) => 
                           MuxOutputs_14_49_port, Y(48) => 
                           MuxOutputs_14_48_port, Y(47) => 
                           MuxOutputs_14_47_port, Y(46) => 
                           MuxOutputs_14_46_port, Y(45) => 
                           MuxOutputs_14_45_port, Y(44) => 
                           MuxOutputs_14_44_port, Y(43) => 
                           MuxOutputs_14_43_port, Y(42) => 
                           MuxOutputs_14_42_port, Y(41) => 
                           MuxOutputs_14_41_port, Y(40) => 
                           MuxOutputs_14_40_port, Y(39) => 
                           MuxOutputs_14_39_port, Y(38) => 
                           MuxOutputs_14_38_port, Y(37) => 
                           MuxOutputs_14_37_port, Y(36) => 
                           MuxOutputs_14_36_port, Y(35) => 
                           MuxOutputs_14_35_port, Y(34) => 
                           MuxOutputs_14_34_port, Y(33) => 
                           MuxOutputs_14_33_port, Y(32) => 
                           MuxOutputs_14_32_port, Y(31) => 
                           MuxOutputs_14_31_port, Y(30) => 
                           MuxOutputs_14_30_port, Y(29) => 
                           MuxOutputs_14_29_port, Y(28) => 
                           MuxOutputs_14_28_port, Y(27) => 
                           MuxOutputs_14_27_port, Y(26) => 
                           MuxOutputs_14_26_port, Y(25) => 
                           MuxOutputs_14_25_port, Y(24) => 
                           MuxOutputs_14_24_port, Y(23) => 
                           MuxOutputs_14_23_port, Y(22) => 
                           MuxOutputs_14_22_port, Y(21) => 
                           MuxOutputs_14_21_port, Y(20) => 
                           MuxOutputs_14_20_port, Y(19) => 
                           MuxOutputs_14_19_port, Y(18) => 
                           MuxOutputs_14_18_port, Y(17) => 
                           MuxOutputs_14_17_port, Y(16) => 
                           MuxOutputs_14_16_port, Y(15) => 
                           MuxOutputs_14_15_port, Y(14) => 
                           MuxOutputs_14_14_port, Y(13) => 
                           MuxOutputs_14_13_port, Y(12) => 
                           MuxOutputs_14_12_port, Y(11) => 
                           MuxOutputs_14_11_port, Y(10) => 
                           MuxOutputs_14_10_port, Y(9) => MuxOutputs_14_9_port,
                           Y(8) => MuxOutputs_14_8_port, Y(7) => 
                           MuxOutputs_14_7_port, Y(6) => MuxOutputs_14_6_port, 
                           Y(5) => MuxOutputs_14_5_port, Y(4) => 
                           MuxOutputs_14_4_port, Y(3) => MuxOutputs_14_3_port, 
                           Y(2) => MuxOutputs_14_2_port, Y(1) => 
                           MuxOutputs_14_1_port, Y(0) => MuxOutputs_14_0_port);
   encoderI_15 : encoder_1 port map( pieceofB(2) => B(31), pieceofB(1) => B(30)
                           , pieceofB(0) => B(29), sel(2) => sel_15_2_port, 
                           sel(1) => sel_15_1_port, sel(0) => sel_15_0_port);
   MUXI_15 : MUX51_MuxNbit64_1 port map( zeroSignal(63) => X_Logic0_port, 
                           zeroSignal(62) => X_Logic0_port, zeroSignal(61) => 
                           X_Logic0_port, zeroSignal(60) => X_Logic0_port, 
                           zeroSignal(59) => X_Logic0_port, zeroSignal(58) => 
                           X_Logic0_port, zeroSignal(57) => X_Logic0_port, 
                           zeroSignal(56) => X_Logic0_port, zeroSignal(55) => 
                           X_Logic0_port, zeroSignal(54) => X_Logic0_port, 
                           zeroSignal(53) => X_Logic0_port, zeroSignal(52) => 
                           X_Logic0_port, zeroSignal(51) => X_Logic0_port, 
                           zeroSignal(50) => X_Logic0_port, zeroSignal(49) => 
                           X_Logic0_port, zeroSignal(48) => X_Logic0_port, 
                           zeroSignal(47) => X_Logic0_port, zeroSignal(46) => 
                           X_Logic0_port, zeroSignal(45) => X_Logic0_port, 
                           zeroSignal(44) => X_Logic0_port, zeroSignal(43) => 
                           X_Logic0_port, zeroSignal(42) => X_Logic0_port, 
                           zeroSignal(41) => X_Logic0_port, zeroSignal(40) => 
                           X_Logic0_port, zeroSignal(39) => X_Logic0_port, 
                           zeroSignal(38) => X_Logic0_port, zeroSignal(37) => 
                           X_Logic0_port, zeroSignal(36) => X_Logic0_port, 
                           zeroSignal(35) => X_Logic0_port, zeroSignal(34) => 
                           X_Logic0_port, zeroSignal(33) => X_Logic0_port, 
                           zeroSignal(32) => X_Logic0_port, zeroSignal(31) => 
                           X_Logic0_port, zeroSignal(30) => X_Logic0_port, 
                           zeroSignal(29) => X_Logic0_port, zeroSignal(28) => 
                           X_Logic0_port, zeroSignal(27) => X_Logic0_port, 
                           zeroSignal(26) => X_Logic0_port, zeroSignal(25) => 
                           X_Logic0_port, zeroSignal(24) => X_Logic0_port, 
                           zeroSignal(23) => X_Logic0_port, zeroSignal(22) => 
                           X_Logic0_port, zeroSignal(21) => X_Logic0_port, 
                           zeroSignal(20) => X_Logic0_port, zeroSignal(19) => 
                           X_Logic0_port, zeroSignal(18) => X_Logic0_port, 
                           zeroSignal(17) => X_Logic0_port, zeroSignal(16) => 
                           X_Logic0_port, zeroSignal(15) => X_Logic0_port, 
                           zeroSignal(14) => X_Logic0_port, zeroSignal(13) => 
                           X_Logic0_port, zeroSignal(12) => X_Logic0_port, 
                           zeroSignal(11) => X_Logic0_port, zeroSignal(10) => 
                           X_Logic0_port, zeroSignal(9) => X_Logic0_port, 
                           zeroSignal(8) => X_Logic0_port, zeroSignal(7) => 
                           X_Logic0_port, zeroSignal(6) => X_Logic0_port, 
                           zeroSignal(5) => X_Logic0_port, zeroSignal(4) => 
                           X_Logic0_port, zeroSignal(3) => X_Logic0_port, 
                           zeroSignal(2) => X_Logic0_port, zeroSignal(1) => 
                           X_Logic0_port, zeroSignal(0) => X_Logic0_port, 
                           A_signal(63) => positive_inputs_30_63_port, 
                           A_signal(62) => positive_inputs_30_62_port, 
                           A_signal(61) => positive_inputs_30_61_port, 
                           A_signal(60) => positive_inputs_30_60_port, 
                           A_signal(59) => positive_inputs_30_59_port, 
                           A_signal(58) => positive_inputs_30_58_port, 
                           A_signal(57) => positive_inputs_30_57_port, 
                           A_signal(56) => positive_inputs_30_56_port, 
                           A_signal(55) => positive_inputs_30_55_port, 
                           A_signal(54) => positive_inputs_30_54_port, 
                           A_signal(53) => positive_inputs_30_53_port, 
                           A_signal(52) => positive_inputs_30_52_port, 
                           A_signal(51) => positive_inputs_30_51_port, 
                           A_signal(50) => positive_inputs_30_50_port, 
                           A_signal(49) => positive_inputs_30_49_port, 
                           A_signal(48) => positive_inputs_30_48_port, 
                           A_signal(47) => positive_inputs_30_47_port, 
                           A_signal(46) => positive_inputs_30_46_port, 
                           A_signal(45) => positive_inputs_30_45_port, 
                           A_signal(44) => positive_inputs_30_44_port, 
                           A_signal(43) => positive_inputs_30_43_port, 
                           A_signal(42) => positive_inputs_30_42_port, 
                           A_signal(41) => positive_inputs_30_41_port, 
                           A_signal(40) => positive_inputs_30_40_port, 
                           A_signal(39) => positive_inputs_30_39_port, 
                           A_signal(38) => positive_inputs_30_38_port, 
                           A_signal(37) => positive_inputs_30_37_port, 
                           A_signal(36) => positive_inputs_30_36_port, 
                           A_signal(35) => positive_inputs_30_35_port, 
                           A_signal(34) => positive_inputs_30_34_port, 
                           A_signal(33) => positive_inputs_30_33_port, 
                           A_signal(32) => positive_inputs_30_32_port, 
                           A_signal(31) => positive_inputs_30_31_port, 
                           A_signal(30) => positive_inputs_30_30_port, 
                           A_signal(29) => positive_inputs_30_29_port, 
                           A_signal(28) => positive_inputs_30_28_port, 
                           A_signal(27) => positive_inputs_30_27_port, 
                           A_signal(26) => positive_inputs_30_26_port, 
                           A_signal(25) => positive_inputs_30_25_port, 
                           A_signal(24) => positive_inputs_30_24_port, 
                           A_signal(23) => positive_inputs_30_23_port, 
                           A_signal(22) => positive_inputs_30_22_port, 
                           A_signal(21) => positive_inputs_30_21_port, 
                           A_signal(20) => positive_inputs_30_20_port, 
                           A_signal(19) => positive_inputs_30_19_port, 
                           A_signal(18) => positive_inputs_30_18_port, 
                           A_signal(17) => positive_inputs_30_17_port, 
                           A_signal(16) => positive_inputs_30_16_port, 
                           A_signal(15) => positive_inputs_30_15_port, 
                           A_signal(14) => positive_inputs_30_14_port, 
                           A_signal(13) => positive_inputs_30_13_port, 
                           A_signal(12) => positive_inputs_30_12_port, 
                           A_signal(11) => positive_inputs_30_11_port, 
                           A_signal(10) => positive_inputs_30_10_port, 
                           A_signal(9) => positive_inputs_30_9_port, 
                           A_signal(8) => positive_inputs_30_8_port, 
                           A_signal(7) => positive_inputs_30_7_port, 
                           A_signal(6) => positive_inputs_30_6_port, 
                           A_signal(5) => positive_inputs_30_5_port, 
                           A_signal(4) => positive_inputs_30_4_port, 
                           A_signal(3) => positive_inputs_30_3_port, 
                           A_signal(2) => positive_inputs_30_2_port, 
                           A_signal(1) => positive_inputs_30_1_port, 
                           A_signal(0) => n9, A_neg(63) => 
                           negative_inputs_30_63_port, A_neg(62) => 
                           negative_inputs_30_62_port, A_neg(61) => 
                           negative_inputs_30_61_port, A_neg(60) => 
                           negative_inputs_30_60_port, A_neg(59) => 
                           negative_inputs_30_59_port, A_neg(58) => 
                           negative_inputs_30_58_port, A_neg(57) => 
                           negative_inputs_30_57_port, A_neg(56) => 
                           negative_inputs_30_56_port, A_neg(55) => 
                           negative_inputs_30_55_port, A_neg(54) => 
                           negative_inputs_30_54_port, A_neg(53) => 
                           negative_inputs_30_53_port, A_neg(52) => 
                           negative_inputs_30_52_port, A_neg(51) => 
                           negative_inputs_30_51_port, A_neg(50) => 
                           negative_inputs_30_50_port, A_neg(49) => 
                           negative_inputs_30_49_port, A_neg(48) => 
                           negative_inputs_30_48_port, A_neg(47) => 
                           negative_inputs_30_47_port, A_neg(46) => 
                           negative_inputs_30_46_port, A_neg(45) => 
                           negative_inputs_30_45_port, A_neg(44) => 
                           negative_inputs_30_44_port, A_neg(43) => 
                           negative_inputs_30_43_port, A_neg(42) => 
                           negative_inputs_30_42_port, A_neg(41) => 
                           negative_inputs_30_41_port, A_neg(40) => 
                           negative_inputs_30_40_port, A_neg(39) => 
                           negative_inputs_30_39_port, A_neg(38) => 
                           negative_inputs_30_38_port, A_neg(37) => 
                           negative_inputs_30_37_port, A_neg(36) => 
                           negative_inputs_30_36_port, A_neg(35) => 
                           negative_inputs_30_35_port, A_neg(34) => 
                           negative_inputs_30_34_port, A_neg(33) => 
                           negative_inputs_30_33_port, A_neg(32) => 
                           negative_inputs_30_32_port, A_neg(31) => 
                           negative_inputs_30_31_port, A_neg(30) => 
                           negative_inputs_30_30_port, A_neg(29) => 
                           negative_inputs_30_29_port, A_neg(28) => 
                           negative_inputs_30_28_port, A_neg(27) => 
                           negative_inputs_30_27_port, A_neg(26) => 
                           negative_inputs_30_26_port, A_neg(25) => 
                           negative_inputs_30_25_port, A_neg(24) => 
                           negative_inputs_30_24_port, A_neg(23) => 
                           negative_inputs_30_23_port, A_neg(22) => 
                           negative_inputs_30_22_port, A_neg(21) => 
                           negative_inputs_30_21_port, A_neg(20) => 
                           negative_inputs_30_20_port, A_neg(19) => 
                           negative_inputs_30_19_port, A_neg(18) => 
                           negative_inputs_30_18_port, A_neg(17) => 
                           negative_inputs_30_17_port, A_neg(16) => 
                           negative_inputs_30_16_port, A_neg(15) => 
                           negative_inputs_30_15_port, A_neg(14) => 
                           negative_inputs_30_14_port, A_neg(13) => 
                           negative_inputs_30_13_port, A_neg(12) => 
                           negative_inputs_30_12_port, A_neg(11) => 
                           negative_inputs_30_11_port, A_neg(10) => 
                           negative_inputs_30_10_port, A_neg(9) => 
                           negative_inputs_30_9_port, A_neg(8) => 
                           negative_inputs_30_8_port, A_neg(7) => 
                           negative_inputs_30_7_port, A_neg(6) => 
                           negative_inputs_30_6_port, A_neg(5) => 
                           negative_inputs_30_5_port, A_neg(4) => 
                           negative_inputs_30_4_port, A_neg(3) => 
                           negative_inputs_30_3_port, A_neg(2) => 
                           negative_inputs_30_2_port, A_neg(1) => 
                           negative_inputs_30_1_port, A_neg(0) => n9, 
                           A_shifted(63) => positive_inputs_31_63_port, 
                           A_shifted(62) => positive_inputs_31_62_port, 
                           A_shifted(61) => positive_inputs_31_61_port, 
                           A_shifted(60) => positive_inputs_31_60_port, 
                           A_shifted(59) => positive_inputs_31_59_port, 
                           A_shifted(58) => positive_inputs_31_58_port, 
                           A_shifted(57) => positive_inputs_31_57_port, 
                           A_shifted(56) => positive_inputs_31_56_port, 
                           A_shifted(55) => positive_inputs_31_55_port, 
                           A_shifted(54) => positive_inputs_31_54_port, 
                           A_shifted(53) => positive_inputs_31_53_port, 
                           A_shifted(52) => positive_inputs_31_52_port, 
                           A_shifted(51) => positive_inputs_31_51_port, 
                           A_shifted(50) => positive_inputs_31_50_port, 
                           A_shifted(49) => positive_inputs_31_49_port, 
                           A_shifted(48) => positive_inputs_31_48_port, 
                           A_shifted(47) => positive_inputs_31_47_port, 
                           A_shifted(46) => positive_inputs_31_46_port, 
                           A_shifted(45) => positive_inputs_31_45_port, 
                           A_shifted(44) => positive_inputs_31_44_port, 
                           A_shifted(43) => positive_inputs_31_43_port, 
                           A_shifted(42) => positive_inputs_31_42_port, 
                           A_shifted(41) => positive_inputs_31_41_port, 
                           A_shifted(40) => positive_inputs_31_40_port, 
                           A_shifted(39) => positive_inputs_31_39_port, 
                           A_shifted(38) => positive_inputs_31_38_port, 
                           A_shifted(37) => positive_inputs_31_37_port, 
                           A_shifted(36) => positive_inputs_31_36_port, 
                           A_shifted(35) => positive_inputs_31_35_port, 
                           A_shifted(34) => positive_inputs_31_34_port, 
                           A_shifted(33) => positive_inputs_31_33_port, 
                           A_shifted(32) => positive_inputs_31_32_port, 
                           A_shifted(31) => positive_inputs_31_31_port, 
                           A_shifted(30) => positive_inputs_31_30_port, 
                           A_shifted(29) => positive_inputs_31_29_port, 
                           A_shifted(28) => positive_inputs_31_28_port, 
                           A_shifted(27) => positive_inputs_31_27_port, 
                           A_shifted(26) => positive_inputs_31_26_port, 
                           A_shifted(25) => positive_inputs_31_25_port, 
                           A_shifted(24) => positive_inputs_31_24_port, 
                           A_shifted(23) => positive_inputs_31_23_port, 
                           A_shifted(22) => positive_inputs_31_22_port, 
                           A_shifted(21) => positive_inputs_31_21_port, 
                           A_shifted(20) => positive_inputs_31_20_port, 
                           A_shifted(19) => positive_inputs_31_19_port, 
                           A_shifted(18) => positive_inputs_31_18_port, 
                           A_shifted(17) => positive_inputs_31_17_port, 
                           A_shifted(16) => positive_inputs_31_16_port, 
                           A_shifted(15) => positive_inputs_31_15_port, 
                           A_shifted(14) => positive_inputs_31_14_port, 
                           A_shifted(13) => positive_inputs_31_13_port, 
                           A_shifted(12) => positive_inputs_31_12_port, 
                           A_shifted(11) => positive_inputs_31_11_port, 
                           A_shifted(10) => positive_inputs_31_10_port, 
                           A_shifted(9) => positive_inputs_31_9_port, 
                           A_shifted(8) => positive_inputs_31_8_port, 
                           A_shifted(7) => positive_inputs_31_7_port, 
                           A_shifted(6) => positive_inputs_31_6_port, 
                           A_shifted(5) => positive_inputs_31_5_port, 
                           A_shifted(4) => positive_inputs_31_4_port, 
                           A_shifted(3) => positive_inputs_31_3_port, 
                           A_shifted(2) => positive_inputs_31_2_port, 
                           A_shifted(1) => positive_inputs_31_1_port, 
                           A_shifted(0) => n9, A_neg_shifted(63) => 
                           negative_inputs_31_63_port, A_neg_shifted(62) => 
                           negative_inputs_31_62_port, A_neg_shifted(61) => 
                           negative_inputs_31_61_port, A_neg_shifted(60) => 
                           negative_inputs_31_60_port, A_neg_shifted(59) => 
                           negative_inputs_31_59_port, A_neg_shifted(58) => 
                           negative_inputs_31_58_port, A_neg_shifted(57) => 
                           negative_inputs_31_57_port, A_neg_shifted(56) => 
                           negative_inputs_31_56_port, A_neg_shifted(55) => 
                           negative_inputs_31_55_port, A_neg_shifted(54) => 
                           negative_inputs_31_54_port, A_neg_shifted(53) => 
                           negative_inputs_31_53_port, A_neg_shifted(52) => 
                           negative_inputs_31_52_port, A_neg_shifted(51) => 
                           negative_inputs_31_51_port, A_neg_shifted(50) => 
                           negative_inputs_31_50_port, A_neg_shifted(49) => 
                           negative_inputs_31_49_port, A_neg_shifted(48) => 
                           negative_inputs_31_48_port, A_neg_shifted(47) => 
                           negative_inputs_31_47_port, A_neg_shifted(46) => 
                           negative_inputs_31_46_port, A_neg_shifted(45) => 
                           negative_inputs_31_45_port, A_neg_shifted(44) => 
                           negative_inputs_31_44_port, A_neg_shifted(43) => 
                           negative_inputs_31_43_port, A_neg_shifted(42) => 
                           negative_inputs_31_42_port, A_neg_shifted(41) => 
                           negative_inputs_31_41_port, A_neg_shifted(40) => 
                           negative_inputs_31_40_port, A_neg_shifted(39) => 
                           negative_inputs_31_39_port, A_neg_shifted(38) => 
                           negative_inputs_31_38_port, A_neg_shifted(37) => 
                           negative_inputs_31_37_port, A_neg_shifted(36) => 
                           negative_inputs_31_36_port, A_neg_shifted(35) => 
                           negative_inputs_31_35_port, A_neg_shifted(34) => 
                           negative_inputs_31_34_port, A_neg_shifted(33) => 
                           negative_inputs_31_33_port, A_neg_shifted(32) => 
                           negative_inputs_31_32_port, A_neg_shifted(31) => 
                           negative_inputs_31_31_port, A_neg_shifted(30) => 
                           negative_inputs_31_30_port, A_neg_shifted(29) => 
                           negative_inputs_31_29_port, A_neg_shifted(28) => 
                           negative_inputs_31_28_port, A_neg_shifted(27) => 
                           negative_inputs_31_27_port, A_neg_shifted(26) => 
                           negative_inputs_31_26_port, A_neg_shifted(25) => 
                           negative_inputs_31_25_port, A_neg_shifted(24) => 
                           negative_inputs_31_24_port, A_neg_shifted(23) => 
                           negative_inputs_31_23_port, A_neg_shifted(22) => 
                           negative_inputs_31_22_port, A_neg_shifted(21) => 
                           negative_inputs_31_21_port, A_neg_shifted(20) => 
                           negative_inputs_31_20_port, A_neg_shifted(19) => 
                           negative_inputs_31_19_port, A_neg_shifted(18) => 
                           negative_inputs_31_18_port, A_neg_shifted(17) => 
                           negative_inputs_31_17_port, A_neg_shifted(16) => 
                           negative_inputs_31_16_port, A_neg_shifted(15) => 
                           negative_inputs_31_15_port, A_neg_shifted(14) => 
                           negative_inputs_31_14_port, A_neg_shifted(13) => 
                           negative_inputs_31_13_port, A_neg_shifted(12) => 
                           negative_inputs_31_12_port, A_neg_shifted(11) => 
                           negative_inputs_31_11_port, A_neg_shifted(10) => 
                           negative_inputs_31_10_port, A_neg_shifted(9) => 
                           negative_inputs_31_9_port, A_neg_shifted(8) => 
                           negative_inputs_31_8_port, A_neg_shifted(7) => 
                           negative_inputs_31_7_port, A_neg_shifted(6) => 
                           negative_inputs_31_6_port, A_neg_shifted(5) => 
                           negative_inputs_31_5_port, A_neg_shifted(4) => 
                           negative_inputs_31_4_port, A_neg_shifted(3) => 
                           negative_inputs_31_3_port, A_neg_shifted(2) => 
                           negative_inputs_31_2_port, A_neg_shifted(1) => 
                           negative_inputs_31_1_port, A_neg_shifted(0) => n9, 
                           Sel(2) => sel_15_2_port, Sel(1) => sel_15_1_port, 
                           Sel(0) => sel_15_0_port, Y(63) => 
                           MuxOutputs_15_63_port, Y(62) => 
                           MuxOutputs_15_62_port, Y(61) => 
                           MuxOutputs_15_61_port, Y(60) => 
                           MuxOutputs_15_60_port, Y(59) => 
                           MuxOutputs_15_59_port, Y(58) => 
                           MuxOutputs_15_58_port, Y(57) => 
                           MuxOutputs_15_57_port, Y(56) => 
                           MuxOutputs_15_56_port, Y(55) => 
                           MuxOutputs_15_55_port, Y(54) => 
                           MuxOutputs_15_54_port, Y(53) => 
                           MuxOutputs_15_53_port, Y(52) => 
                           MuxOutputs_15_52_port, Y(51) => 
                           MuxOutputs_15_51_port, Y(50) => 
                           MuxOutputs_15_50_port, Y(49) => 
                           MuxOutputs_15_49_port, Y(48) => 
                           MuxOutputs_15_48_port, Y(47) => 
                           MuxOutputs_15_47_port, Y(46) => 
                           MuxOutputs_15_46_port, Y(45) => 
                           MuxOutputs_15_45_port, Y(44) => 
                           MuxOutputs_15_44_port, Y(43) => 
                           MuxOutputs_15_43_port, Y(42) => 
                           MuxOutputs_15_42_port, Y(41) => 
                           MuxOutputs_15_41_port, Y(40) => 
                           MuxOutputs_15_40_port, Y(39) => 
                           MuxOutputs_15_39_port, Y(38) => 
                           MuxOutputs_15_38_port, Y(37) => 
                           MuxOutputs_15_37_port, Y(36) => 
                           MuxOutputs_15_36_port, Y(35) => 
                           MuxOutputs_15_35_port, Y(34) => 
                           MuxOutputs_15_34_port, Y(33) => 
                           MuxOutputs_15_33_port, Y(32) => 
                           MuxOutputs_15_32_port, Y(31) => 
                           MuxOutputs_15_31_port, Y(30) => 
                           MuxOutputs_15_30_port, Y(29) => 
                           MuxOutputs_15_29_port, Y(28) => 
                           MuxOutputs_15_28_port, Y(27) => 
                           MuxOutputs_15_27_port, Y(26) => 
                           MuxOutputs_15_26_port, Y(25) => 
                           MuxOutputs_15_25_port, Y(24) => 
                           MuxOutputs_15_24_port, Y(23) => 
                           MuxOutputs_15_23_port, Y(22) => 
                           MuxOutputs_15_22_port, Y(21) => 
                           MuxOutputs_15_21_port, Y(20) => 
                           MuxOutputs_15_20_port, Y(19) => 
                           MuxOutputs_15_19_port, Y(18) => 
                           MuxOutputs_15_18_port, Y(17) => 
                           MuxOutputs_15_17_port, Y(16) => 
                           MuxOutputs_15_16_port, Y(15) => 
                           MuxOutputs_15_15_port, Y(14) => 
                           MuxOutputs_15_14_port, Y(13) => 
                           MuxOutputs_15_13_port, Y(12) => 
                           MuxOutputs_15_12_port, Y(11) => 
                           MuxOutputs_15_11_port, Y(10) => 
                           MuxOutputs_15_10_port, Y(9) => MuxOutputs_15_9_port,
                           Y(8) => MuxOutputs_15_8_port, Y(7) => 
                           MuxOutputs_15_7_port, Y(6) => MuxOutputs_15_6_port, 
                           Y(5) => MuxOutputs_15_5_port, Y(4) => 
                           MuxOutputs_15_4_port, Y(3) => MuxOutputs_15_3_port, 
                           Y(2) => MuxOutputs_15_2_port, Y(1) => 
                           MuxOutputs_15_1_port, Y(0) => MuxOutputs_15_0_port);
   SUM0 : RCA_NbitRca64_15 port map( A(63) => MuxOutputs_0_63_port, A(62) => 
                           MuxOutputs_0_62_port, A(61) => MuxOutputs_0_61_port,
                           A(60) => MuxOutputs_0_60_port, A(59) => 
                           MuxOutputs_0_59_port, A(58) => MuxOutputs_0_58_port,
                           A(57) => MuxOutputs_0_57_port, A(56) => 
                           MuxOutputs_0_56_port, A(55) => MuxOutputs_0_55_port,
                           A(54) => MuxOutputs_0_54_port, A(53) => 
                           MuxOutputs_0_53_port, A(52) => MuxOutputs_0_52_port,
                           A(51) => MuxOutputs_0_51_port, A(50) => 
                           MuxOutputs_0_50_port, A(49) => MuxOutputs_0_49_port,
                           A(48) => MuxOutputs_0_48_port, A(47) => 
                           MuxOutputs_0_47_port, A(46) => MuxOutputs_0_46_port,
                           A(45) => MuxOutputs_0_45_port, A(44) => 
                           MuxOutputs_0_44_port, A(43) => MuxOutputs_0_43_port,
                           A(42) => MuxOutputs_0_42_port, A(41) => 
                           MuxOutputs_0_41_port, A(40) => MuxOutputs_0_40_port,
                           A(39) => MuxOutputs_0_39_port, A(38) => 
                           MuxOutputs_0_38_port, A(37) => MuxOutputs_0_37_port,
                           A(36) => MuxOutputs_0_36_port, A(35) => 
                           MuxOutputs_0_35_port, A(34) => MuxOutputs_0_34_port,
                           A(33) => MuxOutputs_0_33_port, A(32) => 
                           MuxOutputs_0_32_port, A(31) => MuxOutputs_0_31_port,
                           A(30) => MuxOutputs_0_30_port, A(29) => 
                           MuxOutputs_0_29_port, A(28) => MuxOutputs_0_28_port,
                           A(27) => MuxOutputs_0_27_port, A(26) => 
                           MuxOutputs_0_26_port, A(25) => MuxOutputs_0_25_port,
                           A(24) => MuxOutputs_0_24_port, A(23) => 
                           MuxOutputs_0_23_port, A(22) => MuxOutputs_0_22_port,
                           A(21) => MuxOutputs_0_21_port, A(20) => 
                           MuxOutputs_0_20_port, A(19) => MuxOutputs_0_19_port,
                           A(18) => MuxOutputs_0_18_port, A(17) => 
                           MuxOutputs_0_17_port, A(16) => MuxOutputs_0_16_port,
                           A(15) => MuxOutputs_0_15_port, A(14) => 
                           MuxOutputs_0_14_port, A(13) => MuxOutputs_0_13_port,
                           A(12) => MuxOutputs_0_12_port, A(11) => 
                           MuxOutputs_0_11_port, A(10) => MuxOutputs_0_10_port,
                           A(9) => MuxOutputs_0_9_port, A(8) => 
                           MuxOutputs_0_8_port, A(7) => MuxOutputs_0_7_port, 
                           A(6) => MuxOutputs_0_6_port, A(5) => 
                           MuxOutputs_0_5_port, A(4) => MuxOutputs_0_4_port, 
                           A(3) => MuxOutputs_0_3_port, A(2) => 
                           MuxOutputs_0_2_port, A(1) => MuxOutputs_0_1_port, 
                           A(0) => MuxOutputs_0_0_port, B(63) => 
                           MuxOutputs_1_63_port, B(62) => MuxOutputs_1_62_port,
                           B(61) => MuxOutputs_1_61_port, B(60) => 
                           MuxOutputs_1_60_port, B(59) => MuxOutputs_1_59_port,
                           B(58) => MuxOutputs_1_58_port, B(57) => 
                           MuxOutputs_1_57_port, B(56) => MuxOutputs_1_56_port,
                           B(55) => MuxOutputs_1_55_port, B(54) => 
                           MuxOutputs_1_54_port, B(53) => MuxOutputs_1_53_port,
                           B(52) => MuxOutputs_1_52_port, B(51) => 
                           MuxOutputs_1_51_port, B(50) => MuxOutputs_1_50_port,
                           B(49) => MuxOutputs_1_49_port, B(48) => 
                           MuxOutputs_1_48_port, B(47) => MuxOutputs_1_47_port,
                           B(46) => MuxOutputs_1_46_port, B(45) => 
                           MuxOutputs_1_45_port, B(44) => MuxOutputs_1_44_port,
                           B(43) => MuxOutputs_1_43_port, B(42) => 
                           MuxOutputs_1_42_port, B(41) => MuxOutputs_1_41_port,
                           B(40) => MuxOutputs_1_40_port, B(39) => 
                           MuxOutputs_1_39_port, B(38) => MuxOutputs_1_38_port,
                           B(37) => MuxOutputs_1_37_port, B(36) => 
                           MuxOutputs_1_36_port, B(35) => MuxOutputs_1_35_port,
                           B(34) => MuxOutputs_1_34_port, B(33) => 
                           MuxOutputs_1_33_port, B(32) => MuxOutputs_1_32_port,
                           B(31) => MuxOutputs_1_31_port, B(30) => 
                           MuxOutputs_1_30_port, B(29) => MuxOutputs_1_29_port,
                           B(28) => MuxOutputs_1_28_port, B(27) => 
                           MuxOutputs_1_27_port, B(26) => MuxOutputs_1_26_port,
                           B(25) => MuxOutputs_1_25_port, B(24) => 
                           MuxOutputs_1_24_port, B(23) => MuxOutputs_1_23_port,
                           B(22) => MuxOutputs_1_22_port, B(21) => 
                           MuxOutputs_1_21_port, B(20) => MuxOutputs_1_20_port,
                           B(19) => MuxOutputs_1_19_port, B(18) => 
                           MuxOutputs_1_18_port, B(17) => MuxOutputs_1_17_port,
                           B(16) => MuxOutputs_1_16_port, B(15) => 
                           MuxOutputs_1_15_port, B(14) => MuxOutputs_1_14_port,
                           B(13) => MuxOutputs_1_13_port, B(12) => 
                           MuxOutputs_1_12_port, B(11) => MuxOutputs_1_11_port,
                           B(10) => MuxOutputs_1_10_port, B(9) => 
                           MuxOutputs_1_9_port, B(8) => MuxOutputs_1_8_port, 
                           B(7) => MuxOutputs_1_7_port, B(6) => 
                           MuxOutputs_1_6_port, B(5) => MuxOutputs_1_5_port, 
                           B(4) => MuxOutputs_1_4_port, B(3) => 
                           MuxOutputs_1_3_port, B(2) => MuxOutputs_1_2_port, 
                           B(1) => MuxOutputs_1_1_port, B(0) => 
                           MuxOutputs_1_0_port, Ci => X_Logic0_port, S(63) => 
                           SumOutputs_0_63_port, S(62) => SumOutputs_0_62_port,
                           S(61) => SumOutputs_0_61_port, S(60) => 
                           SumOutputs_0_60_port, S(59) => SumOutputs_0_59_port,
                           S(58) => SumOutputs_0_58_port, S(57) => 
                           SumOutputs_0_57_port, S(56) => SumOutputs_0_56_port,
                           S(55) => SumOutputs_0_55_port, S(54) => 
                           SumOutputs_0_54_port, S(53) => SumOutputs_0_53_port,
                           S(52) => SumOutputs_0_52_port, S(51) => 
                           SumOutputs_0_51_port, S(50) => SumOutputs_0_50_port,
                           S(49) => SumOutputs_0_49_port, S(48) => 
                           SumOutputs_0_48_port, S(47) => SumOutputs_0_47_port,
                           S(46) => SumOutputs_0_46_port, S(45) => 
                           SumOutputs_0_45_port, S(44) => SumOutputs_0_44_port,
                           S(43) => SumOutputs_0_43_port, S(42) => 
                           SumOutputs_0_42_port, S(41) => SumOutputs_0_41_port,
                           S(40) => SumOutputs_0_40_port, S(39) => 
                           SumOutputs_0_39_port, S(38) => SumOutputs_0_38_port,
                           S(37) => SumOutputs_0_37_port, S(36) => 
                           SumOutputs_0_36_port, S(35) => SumOutputs_0_35_port,
                           S(34) => SumOutputs_0_34_port, S(33) => 
                           SumOutputs_0_33_port, S(32) => SumOutputs_0_32_port,
                           S(31) => SumOutputs_0_31_port, S(30) => 
                           SumOutputs_0_30_port, S(29) => SumOutputs_0_29_port,
                           S(28) => SumOutputs_0_28_port, S(27) => 
                           SumOutputs_0_27_port, S(26) => SumOutputs_0_26_port,
                           S(25) => SumOutputs_0_25_port, S(24) => 
                           SumOutputs_0_24_port, S(23) => SumOutputs_0_23_port,
                           S(22) => SumOutputs_0_22_port, S(21) => 
                           SumOutputs_0_21_port, S(20) => SumOutputs_0_20_port,
                           S(19) => SumOutputs_0_19_port, S(18) => 
                           SumOutputs_0_18_port, S(17) => SumOutputs_0_17_port,
                           S(16) => SumOutputs_0_16_port, S(15) => 
                           SumOutputs_0_15_port, S(14) => SumOutputs_0_14_port,
                           S(13) => SumOutputs_0_13_port, S(12) => 
                           SumOutputs_0_12_port, S(11) => SumOutputs_0_11_port,
                           S(10) => SumOutputs_0_10_port, S(9) => 
                           SumOutputs_0_9_port, S(8) => SumOutputs_0_8_port, 
                           S(7) => SumOutputs_0_7_port, S(6) => 
                           SumOutputs_0_6_port, S(5) => SumOutputs_0_5_port, 
                           S(4) => SumOutputs_0_4_port, S(3) => 
                           SumOutputs_0_3_port, S(2) => SumOutputs_0_2_port, 
                           S(1) => SumOutputs_0_1_port, S(0) => 
                           SumOutputs_0_0_port, Co => n_1127);
   SUMI_1 : RCA_NbitRca64_14 port map( A(63) => MuxOutputs_2_63_port, A(62) => 
                           MuxOutputs_2_62_port, A(61) => MuxOutputs_2_61_port,
                           A(60) => MuxOutputs_2_60_port, A(59) => 
                           MuxOutputs_2_59_port, A(58) => MuxOutputs_2_58_port,
                           A(57) => MuxOutputs_2_57_port, A(56) => 
                           MuxOutputs_2_56_port, A(55) => MuxOutputs_2_55_port,
                           A(54) => MuxOutputs_2_54_port, A(53) => 
                           MuxOutputs_2_53_port, A(52) => MuxOutputs_2_52_port,
                           A(51) => MuxOutputs_2_51_port, A(50) => 
                           MuxOutputs_2_50_port, A(49) => MuxOutputs_2_49_port,
                           A(48) => MuxOutputs_2_48_port, A(47) => 
                           MuxOutputs_2_47_port, A(46) => MuxOutputs_2_46_port,
                           A(45) => MuxOutputs_2_45_port, A(44) => 
                           MuxOutputs_2_44_port, A(43) => MuxOutputs_2_43_port,
                           A(42) => MuxOutputs_2_42_port, A(41) => 
                           MuxOutputs_2_41_port, A(40) => MuxOutputs_2_40_port,
                           A(39) => MuxOutputs_2_39_port, A(38) => 
                           MuxOutputs_2_38_port, A(37) => MuxOutputs_2_37_port,
                           A(36) => MuxOutputs_2_36_port, A(35) => 
                           MuxOutputs_2_35_port, A(34) => MuxOutputs_2_34_port,
                           A(33) => MuxOutputs_2_33_port, A(32) => 
                           MuxOutputs_2_32_port, A(31) => MuxOutputs_2_31_port,
                           A(30) => MuxOutputs_2_30_port, A(29) => 
                           MuxOutputs_2_29_port, A(28) => MuxOutputs_2_28_port,
                           A(27) => MuxOutputs_2_27_port, A(26) => 
                           MuxOutputs_2_26_port, A(25) => MuxOutputs_2_25_port,
                           A(24) => MuxOutputs_2_24_port, A(23) => 
                           MuxOutputs_2_23_port, A(22) => MuxOutputs_2_22_port,
                           A(21) => MuxOutputs_2_21_port, A(20) => 
                           MuxOutputs_2_20_port, A(19) => MuxOutputs_2_19_port,
                           A(18) => MuxOutputs_2_18_port, A(17) => 
                           MuxOutputs_2_17_port, A(16) => MuxOutputs_2_16_port,
                           A(15) => MuxOutputs_2_15_port, A(14) => 
                           MuxOutputs_2_14_port, A(13) => MuxOutputs_2_13_port,
                           A(12) => MuxOutputs_2_12_port, A(11) => 
                           MuxOutputs_2_11_port, A(10) => MuxOutputs_2_10_port,
                           A(9) => MuxOutputs_2_9_port, A(8) => 
                           MuxOutputs_2_8_port, A(7) => MuxOutputs_2_7_port, 
                           A(6) => MuxOutputs_2_6_port, A(5) => 
                           MuxOutputs_2_5_port, A(4) => MuxOutputs_2_4_port, 
                           A(3) => MuxOutputs_2_3_port, A(2) => 
                           MuxOutputs_2_2_port, A(1) => MuxOutputs_2_1_port, 
                           A(0) => MuxOutputs_2_0_port, B(63) => 
                           SumOutputs_0_63_port, B(62) => SumOutputs_0_62_port,
                           B(61) => SumOutputs_0_61_port, B(60) => 
                           SumOutputs_0_60_port, B(59) => SumOutputs_0_59_port,
                           B(58) => SumOutputs_0_58_port, B(57) => 
                           SumOutputs_0_57_port, B(56) => SumOutputs_0_56_port,
                           B(55) => SumOutputs_0_55_port, B(54) => 
                           SumOutputs_0_54_port, B(53) => SumOutputs_0_53_port,
                           B(52) => SumOutputs_0_52_port, B(51) => 
                           SumOutputs_0_51_port, B(50) => SumOutputs_0_50_port,
                           B(49) => SumOutputs_0_49_port, B(48) => 
                           SumOutputs_0_48_port, B(47) => SumOutputs_0_47_port,
                           B(46) => SumOutputs_0_46_port, B(45) => 
                           SumOutputs_0_45_port, B(44) => SumOutputs_0_44_port,
                           B(43) => SumOutputs_0_43_port, B(42) => 
                           SumOutputs_0_42_port, B(41) => SumOutputs_0_41_port,
                           B(40) => SumOutputs_0_40_port, B(39) => 
                           SumOutputs_0_39_port, B(38) => SumOutputs_0_38_port,
                           B(37) => SumOutputs_0_37_port, B(36) => 
                           SumOutputs_0_36_port, B(35) => SumOutputs_0_35_port,
                           B(34) => SumOutputs_0_34_port, B(33) => 
                           SumOutputs_0_33_port, B(32) => SumOutputs_0_32_port,
                           B(31) => SumOutputs_0_31_port, B(30) => 
                           SumOutputs_0_30_port, B(29) => SumOutputs_0_29_port,
                           B(28) => SumOutputs_0_28_port, B(27) => 
                           SumOutputs_0_27_port, B(26) => SumOutputs_0_26_port,
                           B(25) => SumOutputs_0_25_port, B(24) => 
                           SumOutputs_0_24_port, B(23) => SumOutputs_0_23_port,
                           B(22) => SumOutputs_0_22_port, B(21) => 
                           SumOutputs_0_21_port, B(20) => SumOutputs_0_20_port,
                           B(19) => SumOutputs_0_19_port, B(18) => 
                           SumOutputs_0_18_port, B(17) => SumOutputs_0_17_port,
                           B(16) => SumOutputs_0_16_port, B(15) => 
                           SumOutputs_0_15_port, B(14) => SumOutputs_0_14_port,
                           B(13) => SumOutputs_0_13_port, B(12) => 
                           SumOutputs_0_12_port, B(11) => SumOutputs_0_11_port,
                           B(10) => SumOutputs_0_10_port, B(9) => 
                           SumOutputs_0_9_port, B(8) => SumOutputs_0_8_port, 
                           B(7) => SumOutputs_0_7_port, B(6) => 
                           SumOutputs_0_6_port, B(5) => SumOutputs_0_5_port, 
                           B(4) => SumOutputs_0_4_port, B(3) => 
                           SumOutputs_0_3_port, B(2) => SumOutputs_0_2_port, 
                           B(1) => SumOutputs_0_1_port, B(0) => 
                           SumOutputs_0_0_port, Ci => X_Logic0_port, S(63) => 
                           SumOutputs_1_63_port, S(62) => SumOutputs_1_62_port,
                           S(61) => SumOutputs_1_61_port, S(60) => 
                           SumOutputs_1_60_port, S(59) => SumOutputs_1_59_port,
                           S(58) => SumOutputs_1_58_port, S(57) => 
                           SumOutputs_1_57_port, S(56) => SumOutputs_1_56_port,
                           S(55) => SumOutputs_1_55_port, S(54) => 
                           SumOutputs_1_54_port, S(53) => SumOutputs_1_53_port,
                           S(52) => SumOutputs_1_52_port, S(51) => 
                           SumOutputs_1_51_port, S(50) => SumOutputs_1_50_port,
                           S(49) => SumOutputs_1_49_port, S(48) => 
                           SumOutputs_1_48_port, S(47) => SumOutputs_1_47_port,
                           S(46) => SumOutputs_1_46_port, S(45) => 
                           SumOutputs_1_45_port, S(44) => SumOutputs_1_44_port,
                           S(43) => SumOutputs_1_43_port, S(42) => 
                           SumOutputs_1_42_port, S(41) => SumOutputs_1_41_port,
                           S(40) => SumOutputs_1_40_port, S(39) => 
                           SumOutputs_1_39_port, S(38) => SumOutputs_1_38_port,
                           S(37) => SumOutputs_1_37_port, S(36) => 
                           SumOutputs_1_36_port, S(35) => SumOutputs_1_35_port,
                           S(34) => SumOutputs_1_34_port, S(33) => 
                           SumOutputs_1_33_port, S(32) => SumOutputs_1_32_port,
                           S(31) => SumOutputs_1_31_port, S(30) => 
                           SumOutputs_1_30_port, S(29) => SumOutputs_1_29_port,
                           S(28) => SumOutputs_1_28_port, S(27) => 
                           SumOutputs_1_27_port, S(26) => SumOutputs_1_26_port,
                           S(25) => SumOutputs_1_25_port, S(24) => 
                           SumOutputs_1_24_port, S(23) => SumOutputs_1_23_port,
                           S(22) => SumOutputs_1_22_port, S(21) => 
                           SumOutputs_1_21_port, S(20) => SumOutputs_1_20_port,
                           S(19) => SumOutputs_1_19_port, S(18) => 
                           SumOutputs_1_18_port, S(17) => SumOutputs_1_17_port,
                           S(16) => SumOutputs_1_16_port, S(15) => 
                           SumOutputs_1_15_port, S(14) => SumOutputs_1_14_port,
                           S(13) => SumOutputs_1_13_port, S(12) => 
                           SumOutputs_1_12_port, S(11) => SumOutputs_1_11_port,
                           S(10) => SumOutputs_1_10_port, S(9) => 
                           SumOutputs_1_9_port, S(8) => SumOutputs_1_8_port, 
                           S(7) => SumOutputs_1_7_port, S(6) => 
                           SumOutputs_1_6_port, S(5) => SumOutputs_1_5_port, 
                           S(4) => SumOutputs_1_4_port, S(3) => 
                           SumOutputs_1_3_port, S(2) => SumOutputs_1_2_port, 
                           S(1) => SumOutputs_1_1_port, S(0) => 
                           SumOutputs_1_0_port, Co => n_1128);
   SUMI_2 : RCA_NbitRca64_13 port map( A(63) => MuxOutputs_3_63_port, A(62) => 
                           MuxOutputs_3_62_port, A(61) => MuxOutputs_3_61_port,
                           A(60) => MuxOutputs_3_60_port, A(59) => 
                           MuxOutputs_3_59_port, A(58) => MuxOutputs_3_58_port,
                           A(57) => MuxOutputs_3_57_port, A(56) => 
                           MuxOutputs_3_56_port, A(55) => MuxOutputs_3_55_port,
                           A(54) => MuxOutputs_3_54_port, A(53) => 
                           MuxOutputs_3_53_port, A(52) => MuxOutputs_3_52_port,
                           A(51) => MuxOutputs_3_51_port, A(50) => 
                           MuxOutputs_3_50_port, A(49) => MuxOutputs_3_49_port,
                           A(48) => MuxOutputs_3_48_port, A(47) => 
                           MuxOutputs_3_47_port, A(46) => MuxOutputs_3_46_port,
                           A(45) => MuxOutputs_3_45_port, A(44) => 
                           MuxOutputs_3_44_port, A(43) => MuxOutputs_3_43_port,
                           A(42) => MuxOutputs_3_42_port, A(41) => 
                           MuxOutputs_3_41_port, A(40) => MuxOutputs_3_40_port,
                           A(39) => MuxOutputs_3_39_port, A(38) => 
                           MuxOutputs_3_38_port, A(37) => MuxOutputs_3_37_port,
                           A(36) => MuxOutputs_3_36_port, A(35) => 
                           MuxOutputs_3_35_port, A(34) => MuxOutputs_3_34_port,
                           A(33) => MuxOutputs_3_33_port, A(32) => 
                           MuxOutputs_3_32_port, A(31) => MuxOutputs_3_31_port,
                           A(30) => MuxOutputs_3_30_port, A(29) => 
                           MuxOutputs_3_29_port, A(28) => MuxOutputs_3_28_port,
                           A(27) => MuxOutputs_3_27_port, A(26) => 
                           MuxOutputs_3_26_port, A(25) => MuxOutputs_3_25_port,
                           A(24) => MuxOutputs_3_24_port, A(23) => 
                           MuxOutputs_3_23_port, A(22) => MuxOutputs_3_22_port,
                           A(21) => MuxOutputs_3_21_port, A(20) => 
                           MuxOutputs_3_20_port, A(19) => MuxOutputs_3_19_port,
                           A(18) => MuxOutputs_3_18_port, A(17) => 
                           MuxOutputs_3_17_port, A(16) => MuxOutputs_3_16_port,
                           A(15) => MuxOutputs_3_15_port, A(14) => 
                           MuxOutputs_3_14_port, A(13) => MuxOutputs_3_13_port,
                           A(12) => MuxOutputs_3_12_port, A(11) => 
                           MuxOutputs_3_11_port, A(10) => MuxOutputs_3_10_port,
                           A(9) => MuxOutputs_3_9_port, A(8) => 
                           MuxOutputs_3_8_port, A(7) => MuxOutputs_3_7_port, 
                           A(6) => MuxOutputs_3_6_port, A(5) => 
                           MuxOutputs_3_5_port, A(4) => MuxOutputs_3_4_port, 
                           A(3) => MuxOutputs_3_3_port, A(2) => 
                           MuxOutputs_3_2_port, A(1) => MuxOutputs_3_1_port, 
                           A(0) => MuxOutputs_3_0_port, B(63) => 
                           SumOutputs_1_63_port, B(62) => SumOutputs_1_62_port,
                           B(61) => SumOutputs_1_61_port, B(60) => 
                           SumOutputs_1_60_port, B(59) => SumOutputs_1_59_port,
                           B(58) => SumOutputs_1_58_port, B(57) => 
                           SumOutputs_1_57_port, B(56) => SumOutputs_1_56_port,
                           B(55) => SumOutputs_1_55_port, B(54) => 
                           SumOutputs_1_54_port, B(53) => SumOutputs_1_53_port,
                           B(52) => SumOutputs_1_52_port, B(51) => 
                           SumOutputs_1_51_port, B(50) => SumOutputs_1_50_port,
                           B(49) => SumOutputs_1_49_port, B(48) => 
                           SumOutputs_1_48_port, B(47) => SumOutputs_1_47_port,
                           B(46) => SumOutputs_1_46_port, B(45) => 
                           SumOutputs_1_45_port, B(44) => SumOutputs_1_44_port,
                           B(43) => SumOutputs_1_43_port, B(42) => 
                           SumOutputs_1_42_port, B(41) => SumOutputs_1_41_port,
                           B(40) => SumOutputs_1_40_port, B(39) => 
                           SumOutputs_1_39_port, B(38) => SumOutputs_1_38_port,
                           B(37) => SumOutputs_1_37_port, B(36) => 
                           SumOutputs_1_36_port, B(35) => SumOutputs_1_35_port,
                           B(34) => SumOutputs_1_34_port, B(33) => 
                           SumOutputs_1_33_port, B(32) => SumOutputs_1_32_port,
                           B(31) => SumOutputs_1_31_port, B(30) => 
                           SumOutputs_1_30_port, B(29) => SumOutputs_1_29_port,
                           B(28) => SumOutputs_1_28_port, B(27) => 
                           SumOutputs_1_27_port, B(26) => SumOutputs_1_26_port,
                           B(25) => SumOutputs_1_25_port, B(24) => 
                           SumOutputs_1_24_port, B(23) => SumOutputs_1_23_port,
                           B(22) => SumOutputs_1_22_port, B(21) => 
                           SumOutputs_1_21_port, B(20) => SumOutputs_1_20_port,
                           B(19) => SumOutputs_1_19_port, B(18) => 
                           SumOutputs_1_18_port, B(17) => SumOutputs_1_17_port,
                           B(16) => SumOutputs_1_16_port, B(15) => 
                           SumOutputs_1_15_port, B(14) => SumOutputs_1_14_port,
                           B(13) => SumOutputs_1_13_port, B(12) => 
                           SumOutputs_1_12_port, B(11) => SumOutputs_1_11_port,
                           B(10) => SumOutputs_1_10_port, B(9) => 
                           SumOutputs_1_9_port, B(8) => SumOutputs_1_8_port, 
                           B(7) => SumOutputs_1_7_port, B(6) => 
                           SumOutputs_1_6_port, B(5) => SumOutputs_1_5_port, 
                           B(4) => SumOutputs_1_4_port, B(3) => 
                           SumOutputs_1_3_port, B(2) => SumOutputs_1_2_port, 
                           B(1) => SumOutputs_1_1_port, B(0) => 
                           SumOutputs_1_0_port, Ci => X_Logic0_port, S(63) => 
                           SumOutputs_2_63_port, S(62) => SumOutputs_2_62_port,
                           S(61) => SumOutputs_2_61_port, S(60) => 
                           SumOutputs_2_60_port, S(59) => SumOutputs_2_59_port,
                           S(58) => SumOutputs_2_58_port, S(57) => 
                           SumOutputs_2_57_port, S(56) => SumOutputs_2_56_port,
                           S(55) => SumOutputs_2_55_port, S(54) => 
                           SumOutputs_2_54_port, S(53) => SumOutputs_2_53_port,
                           S(52) => SumOutputs_2_52_port, S(51) => 
                           SumOutputs_2_51_port, S(50) => SumOutputs_2_50_port,
                           S(49) => SumOutputs_2_49_port, S(48) => 
                           SumOutputs_2_48_port, S(47) => SumOutputs_2_47_port,
                           S(46) => SumOutputs_2_46_port, S(45) => 
                           SumOutputs_2_45_port, S(44) => SumOutputs_2_44_port,
                           S(43) => SumOutputs_2_43_port, S(42) => 
                           SumOutputs_2_42_port, S(41) => SumOutputs_2_41_port,
                           S(40) => SumOutputs_2_40_port, S(39) => 
                           SumOutputs_2_39_port, S(38) => SumOutputs_2_38_port,
                           S(37) => SumOutputs_2_37_port, S(36) => 
                           SumOutputs_2_36_port, S(35) => SumOutputs_2_35_port,
                           S(34) => SumOutputs_2_34_port, S(33) => 
                           SumOutputs_2_33_port, S(32) => SumOutputs_2_32_port,
                           S(31) => SumOutputs_2_31_port, S(30) => 
                           SumOutputs_2_30_port, S(29) => SumOutputs_2_29_port,
                           S(28) => SumOutputs_2_28_port, S(27) => 
                           SumOutputs_2_27_port, S(26) => SumOutputs_2_26_port,
                           S(25) => SumOutputs_2_25_port, S(24) => 
                           SumOutputs_2_24_port, S(23) => SumOutputs_2_23_port,
                           S(22) => SumOutputs_2_22_port, S(21) => 
                           SumOutputs_2_21_port, S(20) => SumOutputs_2_20_port,
                           S(19) => SumOutputs_2_19_port, S(18) => 
                           SumOutputs_2_18_port, S(17) => SumOutputs_2_17_port,
                           S(16) => SumOutputs_2_16_port, S(15) => 
                           SumOutputs_2_15_port, S(14) => SumOutputs_2_14_port,
                           S(13) => SumOutputs_2_13_port, S(12) => 
                           SumOutputs_2_12_port, S(11) => SumOutputs_2_11_port,
                           S(10) => SumOutputs_2_10_port, S(9) => 
                           SumOutputs_2_9_port, S(8) => SumOutputs_2_8_port, 
                           S(7) => SumOutputs_2_7_port, S(6) => 
                           SumOutputs_2_6_port, S(5) => SumOutputs_2_5_port, 
                           S(4) => SumOutputs_2_4_port, S(3) => 
                           SumOutputs_2_3_port, S(2) => SumOutputs_2_2_port, 
                           S(1) => SumOutputs_2_1_port, S(0) => 
                           SumOutputs_2_0_port, Co => n_1129);
   SUMI_3 : RCA_NbitRca64_12 port map( A(63) => MuxOutputs_4_63_port, A(62) => 
                           MuxOutputs_4_62_port, A(61) => MuxOutputs_4_61_port,
                           A(60) => MuxOutputs_4_60_port, A(59) => 
                           MuxOutputs_4_59_port, A(58) => MuxOutputs_4_58_port,
                           A(57) => MuxOutputs_4_57_port, A(56) => 
                           MuxOutputs_4_56_port, A(55) => MuxOutputs_4_55_port,
                           A(54) => MuxOutputs_4_54_port, A(53) => 
                           MuxOutputs_4_53_port, A(52) => MuxOutputs_4_52_port,
                           A(51) => MuxOutputs_4_51_port, A(50) => 
                           MuxOutputs_4_50_port, A(49) => MuxOutputs_4_49_port,
                           A(48) => MuxOutputs_4_48_port, A(47) => 
                           MuxOutputs_4_47_port, A(46) => MuxOutputs_4_46_port,
                           A(45) => MuxOutputs_4_45_port, A(44) => 
                           MuxOutputs_4_44_port, A(43) => MuxOutputs_4_43_port,
                           A(42) => MuxOutputs_4_42_port, A(41) => 
                           MuxOutputs_4_41_port, A(40) => MuxOutputs_4_40_port,
                           A(39) => MuxOutputs_4_39_port, A(38) => 
                           MuxOutputs_4_38_port, A(37) => MuxOutputs_4_37_port,
                           A(36) => MuxOutputs_4_36_port, A(35) => 
                           MuxOutputs_4_35_port, A(34) => MuxOutputs_4_34_port,
                           A(33) => MuxOutputs_4_33_port, A(32) => 
                           MuxOutputs_4_32_port, A(31) => MuxOutputs_4_31_port,
                           A(30) => MuxOutputs_4_30_port, A(29) => 
                           MuxOutputs_4_29_port, A(28) => MuxOutputs_4_28_port,
                           A(27) => MuxOutputs_4_27_port, A(26) => 
                           MuxOutputs_4_26_port, A(25) => MuxOutputs_4_25_port,
                           A(24) => MuxOutputs_4_24_port, A(23) => 
                           MuxOutputs_4_23_port, A(22) => MuxOutputs_4_22_port,
                           A(21) => MuxOutputs_4_21_port, A(20) => 
                           MuxOutputs_4_20_port, A(19) => MuxOutputs_4_19_port,
                           A(18) => MuxOutputs_4_18_port, A(17) => 
                           MuxOutputs_4_17_port, A(16) => MuxOutputs_4_16_port,
                           A(15) => MuxOutputs_4_15_port, A(14) => 
                           MuxOutputs_4_14_port, A(13) => MuxOutputs_4_13_port,
                           A(12) => MuxOutputs_4_12_port, A(11) => 
                           MuxOutputs_4_11_port, A(10) => MuxOutputs_4_10_port,
                           A(9) => MuxOutputs_4_9_port, A(8) => 
                           MuxOutputs_4_8_port, A(7) => MuxOutputs_4_7_port, 
                           A(6) => MuxOutputs_4_6_port, A(5) => 
                           MuxOutputs_4_5_port, A(4) => MuxOutputs_4_4_port, 
                           A(3) => MuxOutputs_4_3_port, A(2) => 
                           MuxOutputs_4_2_port, A(1) => MuxOutputs_4_1_port, 
                           A(0) => MuxOutputs_4_0_port, B(63) => 
                           SumOutputs_2_63_port, B(62) => SumOutputs_2_62_port,
                           B(61) => SumOutputs_2_61_port, B(60) => 
                           SumOutputs_2_60_port, B(59) => SumOutputs_2_59_port,
                           B(58) => SumOutputs_2_58_port, B(57) => 
                           SumOutputs_2_57_port, B(56) => SumOutputs_2_56_port,
                           B(55) => SumOutputs_2_55_port, B(54) => 
                           SumOutputs_2_54_port, B(53) => SumOutputs_2_53_port,
                           B(52) => SumOutputs_2_52_port, B(51) => 
                           SumOutputs_2_51_port, B(50) => SumOutputs_2_50_port,
                           B(49) => SumOutputs_2_49_port, B(48) => 
                           SumOutputs_2_48_port, B(47) => SumOutputs_2_47_port,
                           B(46) => SumOutputs_2_46_port, B(45) => 
                           SumOutputs_2_45_port, B(44) => SumOutputs_2_44_port,
                           B(43) => SumOutputs_2_43_port, B(42) => 
                           SumOutputs_2_42_port, B(41) => SumOutputs_2_41_port,
                           B(40) => SumOutputs_2_40_port, B(39) => 
                           SumOutputs_2_39_port, B(38) => SumOutputs_2_38_port,
                           B(37) => SumOutputs_2_37_port, B(36) => 
                           SumOutputs_2_36_port, B(35) => SumOutputs_2_35_port,
                           B(34) => SumOutputs_2_34_port, B(33) => 
                           SumOutputs_2_33_port, B(32) => SumOutputs_2_32_port,
                           B(31) => SumOutputs_2_31_port, B(30) => 
                           SumOutputs_2_30_port, B(29) => SumOutputs_2_29_port,
                           B(28) => SumOutputs_2_28_port, B(27) => 
                           SumOutputs_2_27_port, B(26) => SumOutputs_2_26_port,
                           B(25) => SumOutputs_2_25_port, B(24) => 
                           SumOutputs_2_24_port, B(23) => SumOutputs_2_23_port,
                           B(22) => SumOutputs_2_22_port, B(21) => 
                           SumOutputs_2_21_port, B(20) => SumOutputs_2_20_port,
                           B(19) => SumOutputs_2_19_port, B(18) => 
                           SumOutputs_2_18_port, B(17) => SumOutputs_2_17_port,
                           B(16) => SumOutputs_2_16_port, B(15) => 
                           SumOutputs_2_15_port, B(14) => SumOutputs_2_14_port,
                           B(13) => SumOutputs_2_13_port, B(12) => 
                           SumOutputs_2_12_port, B(11) => SumOutputs_2_11_port,
                           B(10) => SumOutputs_2_10_port, B(9) => 
                           SumOutputs_2_9_port, B(8) => SumOutputs_2_8_port, 
                           B(7) => SumOutputs_2_7_port, B(6) => 
                           SumOutputs_2_6_port, B(5) => SumOutputs_2_5_port, 
                           B(4) => SumOutputs_2_4_port, B(3) => 
                           SumOutputs_2_3_port, B(2) => SumOutputs_2_2_port, 
                           B(1) => SumOutputs_2_1_port, B(0) => 
                           SumOutputs_2_0_port, Ci => X_Logic0_port, S(63) => 
                           SumOutputs_3_63_port, S(62) => SumOutputs_3_62_port,
                           S(61) => SumOutputs_3_61_port, S(60) => 
                           SumOutputs_3_60_port, S(59) => SumOutputs_3_59_port,
                           S(58) => SumOutputs_3_58_port, S(57) => 
                           SumOutputs_3_57_port, S(56) => SumOutputs_3_56_port,
                           S(55) => SumOutputs_3_55_port, S(54) => 
                           SumOutputs_3_54_port, S(53) => SumOutputs_3_53_port,
                           S(52) => SumOutputs_3_52_port, S(51) => 
                           SumOutputs_3_51_port, S(50) => SumOutputs_3_50_port,
                           S(49) => SumOutputs_3_49_port, S(48) => 
                           SumOutputs_3_48_port, S(47) => SumOutputs_3_47_port,
                           S(46) => SumOutputs_3_46_port, S(45) => 
                           SumOutputs_3_45_port, S(44) => SumOutputs_3_44_port,
                           S(43) => SumOutputs_3_43_port, S(42) => 
                           SumOutputs_3_42_port, S(41) => SumOutputs_3_41_port,
                           S(40) => SumOutputs_3_40_port, S(39) => 
                           SumOutputs_3_39_port, S(38) => SumOutputs_3_38_port,
                           S(37) => SumOutputs_3_37_port, S(36) => 
                           SumOutputs_3_36_port, S(35) => SumOutputs_3_35_port,
                           S(34) => SumOutputs_3_34_port, S(33) => 
                           SumOutputs_3_33_port, S(32) => SumOutputs_3_32_port,
                           S(31) => SumOutputs_3_31_port, S(30) => 
                           SumOutputs_3_30_port, S(29) => SumOutputs_3_29_port,
                           S(28) => SumOutputs_3_28_port, S(27) => 
                           SumOutputs_3_27_port, S(26) => SumOutputs_3_26_port,
                           S(25) => SumOutputs_3_25_port, S(24) => 
                           SumOutputs_3_24_port, S(23) => SumOutputs_3_23_port,
                           S(22) => SumOutputs_3_22_port, S(21) => 
                           SumOutputs_3_21_port, S(20) => SumOutputs_3_20_port,
                           S(19) => SumOutputs_3_19_port, S(18) => 
                           SumOutputs_3_18_port, S(17) => SumOutputs_3_17_port,
                           S(16) => SumOutputs_3_16_port, S(15) => 
                           SumOutputs_3_15_port, S(14) => SumOutputs_3_14_port,
                           S(13) => SumOutputs_3_13_port, S(12) => 
                           SumOutputs_3_12_port, S(11) => SumOutputs_3_11_port,
                           S(10) => SumOutputs_3_10_port, S(9) => 
                           SumOutputs_3_9_port, S(8) => SumOutputs_3_8_port, 
                           S(7) => SumOutputs_3_7_port, S(6) => 
                           SumOutputs_3_6_port, S(5) => SumOutputs_3_5_port, 
                           S(4) => SumOutputs_3_4_port, S(3) => 
                           SumOutputs_3_3_port, S(2) => SumOutputs_3_2_port, 
                           S(1) => SumOutputs_3_1_port, S(0) => 
                           SumOutputs_3_0_port, Co => n_1130);
   SUMI_4 : RCA_NbitRca64_11 port map( A(63) => MuxOutputs_5_63_port, A(62) => 
                           MuxOutputs_5_62_port, A(61) => MuxOutputs_5_61_port,
                           A(60) => MuxOutputs_5_60_port, A(59) => 
                           MuxOutputs_5_59_port, A(58) => MuxOutputs_5_58_port,
                           A(57) => MuxOutputs_5_57_port, A(56) => 
                           MuxOutputs_5_56_port, A(55) => MuxOutputs_5_55_port,
                           A(54) => MuxOutputs_5_54_port, A(53) => 
                           MuxOutputs_5_53_port, A(52) => MuxOutputs_5_52_port,
                           A(51) => MuxOutputs_5_51_port, A(50) => 
                           MuxOutputs_5_50_port, A(49) => MuxOutputs_5_49_port,
                           A(48) => MuxOutputs_5_48_port, A(47) => 
                           MuxOutputs_5_47_port, A(46) => MuxOutputs_5_46_port,
                           A(45) => MuxOutputs_5_45_port, A(44) => 
                           MuxOutputs_5_44_port, A(43) => MuxOutputs_5_43_port,
                           A(42) => MuxOutputs_5_42_port, A(41) => 
                           MuxOutputs_5_41_port, A(40) => MuxOutputs_5_40_port,
                           A(39) => MuxOutputs_5_39_port, A(38) => 
                           MuxOutputs_5_38_port, A(37) => MuxOutputs_5_37_port,
                           A(36) => MuxOutputs_5_36_port, A(35) => 
                           MuxOutputs_5_35_port, A(34) => MuxOutputs_5_34_port,
                           A(33) => MuxOutputs_5_33_port, A(32) => 
                           MuxOutputs_5_32_port, A(31) => MuxOutputs_5_31_port,
                           A(30) => MuxOutputs_5_30_port, A(29) => 
                           MuxOutputs_5_29_port, A(28) => MuxOutputs_5_28_port,
                           A(27) => MuxOutputs_5_27_port, A(26) => 
                           MuxOutputs_5_26_port, A(25) => MuxOutputs_5_25_port,
                           A(24) => MuxOutputs_5_24_port, A(23) => 
                           MuxOutputs_5_23_port, A(22) => MuxOutputs_5_22_port,
                           A(21) => MuxOutputs_5_21_port, A(20) => 
                           MuxOutputs_5_20_port, A(19) => MuxOutputs_5_19_port,
                           A(18) => MuxOutputs_5_18_port, A(17) => 
                           MuxOutputs_5_17_port, A(16) => MuxOutputs_5_16_port,
                           A(15) => MuxOutputs_5_15_port, A(14) => 
                           MuxOutputs_5_14_port, A(13) => MuxOutputs_5_13_port,
                           A(12) => MuxOutputs_5_12_port, A(11) => 
                           MuxOutputs_5_11_port, A(10) => MuxOutputs_5_10_port,
                           A(9) => MuxOutputs_5_9_port, A(8) => 
                           MuxOutputs_5_8_port, A(7) => MuxOutputs_5_7_port, 
                           A(6) => MuxOutputs_5_6_port, A(5) => 
                           MuxOutputs_5_5_port, A(4) => MuxOutputs_5_4_port, 
                           A(3) => MuxOutputs_5_3_port, A(2) => 
                           MuxOutputs_5_2_port, A(1) => MuxOutputs_5_1_port, 
                           A(0) => MuxOutputs_5_0_port, B(63) => 
                           SumOutputs_3_63_port, B(62) => SumOutputs_3_62_port,
                           B(61) => SumOutputs_3_61_port, B(60) => 
                           SumOutputs_3_60_port, B(59) => SumOutputs_3_59_port,
                           B(58) => SumOutputs_3_58_port, B(57) => 
                           SumOutputs_3_57_port, B(56) => SumOutputs_3_56_port,
                           B(55) => SumOutputs_3_55_port, B(54) => 
                           SumOutputs_3_54_port, B(53) => SumOutputs_3_53_port,
                           B(52) => SumOutputs_3_52_port, B(51) => 
                           SumOutputs_3_51_port, B(50) => SumOutputs_3_50_port,
                           B(49) => SumOutputs_3_49_port, B(48) => 
                           SumOutputs_3_48_port, B(47) => SumOutputs_3_47_port,
                           B(46) => SumOutputs_3_46_port, B(45) => 
                           SumOutputs_3_45_port, B(44) => SumOutputs_3_44_port,
                           B(43) => SumOutputs_3_43_port, B(42) => 
                           SumOutputs_3_42_port, B(41) => SumOutputs_3_41_port,
                           B(40) => SumOutputs_3_40_port, B(39) => 
                           SumOutputs_3_39_port, B(38) => SumOutputs_3_38_port,
                           B(37) => SumOutputs_3_37_port, B(36) => 
                           SumOutputs_3_36_port, B(35) => SumOutputs_3_35_port,
                           B(34) => SumOutputs_3_34_port, B(33) => 
                           SumOutputs_3_33_port, B(32) => SumOutputs_3_32_port,
                           B(31) => SumOutputs_3_31_port, B(30) => 
                           SumOutputs_3_30_port, B(29) => SumOutputs_3_29_port,
                           B(28) => SumOutputs_3_28_port, B(27) => 
                           SumOutputs_3_27_port, B(26) => SumOutputs_3_26_port,
                           B(25) => SumOutputs_3_25_port, B(24) => 
                           SumOutputs_3_24_port, B(23) => SumOutputs_3_23_port,
                           B(22) => SumOutputs_3_22_port, B(21) => 
                           SumOutputs_3_21_port, B(20) => SumOutputs_3_20_port,
                           B(19) => SumOutputs_3_19_port, B(18) => 
                           SumOutputs_3_18_port, B(17) => SumOutputs_3_17_port,
                           B(16) => SumOutputs_3_16_port, B(15) => 
                           SumOutputs_3_15_port, B(14) => SumOutputs_3_14_port,
                           B(13) => SumOutputs_3_13_port, B(12) => 
                           SumOutputs_3_12_port, B(11) => SumOutputs_3_11_port,
                           B(10) => SumOutputs_3_10_port, B(9) => 
                           SumOutputs_3_9_port, B(8) => SumOutputs_3_8_port, 
                           B(7) => SumOutputs_3_7_port, B(6) => 
                           SumOutputs_3_6_port, B(5) => SumOutputs_3_5_port, 
                           B(4) => SumOutputs_3_4_port, B(3) => 
                           SumOutputs_3_3_port, B(2) => SumOutputs_3_2_port, 
                           B(1) => SumOutputs_3_1_port, B(0) => 
                           SumOutputs_3_0_port, Ci => X_Logic0_port, S(63) => 
                           SumOutputs_4_63_port, S(62) => SumOutputs_4_62_port,
                           S(61) => SumOutputs_4_61_port, S(60) => 
                           SumOutputs_4_60_port, S(59) => SumOutputs_4_59_port,
                           S(58) => SumOutputs_4_58_port, S(57) => 
                           SumOutputs_4_57_port, S(56) => SumOutputs_4_56_port,
                           S(55) => SumOutputs_4_55_port, S(54) => 
                           SumOutputs_4_54_port, S(53) => SumOutputs_4_53_port,
                           S(52) => SumOutputs_4_52_port, S(51) => 
                           SumOutputs_4_51_port, S(50) => SumOutputs_4_50_port,
                           S(49) => SumOutputs_4_49_port, S(48) => 
                           SumOutputs_4_48_port, S(47) => SumOutputs_4_47_port,
                           S(46) => SumOutputs_4_46_port, S(45) => 
                           SumOutputs_4_45_port, S(44) => SumOutputs_4_44_port,
                           S(43) => SumOutputs_4_43_port, S(42) => 
                           SumOutputs_4_42_port, S(41) => SumOutputs_4_41_port,
                           S(40) => SumOutputs_4_40_port, S(39) => 
                           SumOutputs_4_39_port, S(38) => SumOutputs_4_38_port,
                           S(37) => SumOutputs_4_37_port, S(36) => 
                           SumOutputs_4_36_port, S(35) => SumOutputs_4_35_port,
                           S(34) => SumOutputs_4_34_port, S(33) => 
                           SumOutputs_4_33_port, S(32) => SumOutputs_4_32_port,
                           S(31) => SumOutputs_4_31_port, S(30) => 
                           SumOutputs_4_30_port, S(29) => SumOutputs_4_29_port,
                           S(28) => SumOutputs_4_28_port, S(27) => 
                           SumOutputs_4_27_port, S(26) => SumOutputs_4_26_port,
                           S(25) => SumOutputs_4_25_port, S(24) => 
                           SumOutputs_4_24_port, S(23) => SumOutputs_4_23_port,
                           S(22) => SumOutputs_4_22_port, S(21) => 
                           SumOutputs_4_21_port, S(20) => SumOutputs_4_20_port,
                           S(19) => SumOutputs_4_19_port, S(18) => 
                           SumOutputs_4_18_port, S(17) => SumOutputs_4_17_port,
                           S(16) => SumOutputs_4_16_port, S(15) => 
                           SumOutputs_4_15_port, S(14) => SumOutputs_4_14_port,
                           S(13) => SumOutputs_4_13_port, S(12) => 
                           SumOutputs_4_12_port, S(11) => SumOutputs_4_11_port,
                           S(10) => SumOutputs_4_10_port, S(9) => 
                           SumOutputs_4_9_port, S(8) => SumOutputs_4_8_port, 
                           S(7) => SumOutputs_4_7_port, S(6) => 
                           SumOutputs_4_6_port, S(5) => SumOutputs_4_5_port, 
                           S(4) => SumOutputs_4_4_port, S(3) => 
                           SumOutputs_4_3_port, S(2) => SumOutputs_4_2_port, 
                           S(1) => SumOutputs_4_1_port, S(0) => 
                           SumOutputs_4_0_port, Co => n_1131);
   SUMI_5 : RCA_NbitRca64_10 port map( A(63) => MuxOutputs_6_63_port, A(62) => 
                           MuxOutputs_6_62_port, A(61) => MuxOutputs_6_61_port,
                           A(60) => MuxOutputs_6_60_port, A(59) => 
                           MuxOutputs_6_59_port, A(58) => MuxOutputs_6_58_port,
                           A(57) => MuxOutputs_6_57_port, A(56) => 
                           MuxOutputs_6_56_port, A(55) => MuxOutputs_6_55_port,
                           A(54) => MuxOutputs_6_54_port, A(53) => 
                           MuxOutputs_6_53_port, A(52) => MuxOutputs_6_52_port,
                           A(51) => MuxOutputs_6_51_port, A(50) => 
                           MuxOutputs_6_50_port, A(49) => MuxOutputs_6_49_port,
                           A(48) => MuxOutputs_6_48_port, A(47) => 
                           MuxOutputs_6_47_port, A(46) => MuxOutputs_6_46_port,
                           A(45) => MuxOutputs_6_45_port, A(44) => 
                           MuxOutputs_6_44_port, A(43) => MuxOutputs_6_43_port,
                           A(42) => MuxOutputs_6_42_port, A(41) => 
                           MuxOutputs_6_41_port, A(40) => MuxOutputs_6_40_port,
                           A(39) => MuxOutputs_6_39_port, A(38) => 
                           MuxOutputs_6_38_port, A(37) => MuxOutputs_6_37_port,
                           A(36) => MuxOutputs_6_36_port, A(35) => 
                           MuxOutputs_6_35_port, A(34) => MuxOutputs_6_34_port,
                           A(33) => MuxOutputs_6_33_port, A(32) => 
                           MuxOutputs_6_32_port, A(31) => MuxOutputs_6_31_port,
                           A(30) => MuxOutputs_6_30_port, A(29) => 
                           MuxOutputs_6_29_port, A(28) => MuxOutputs_6_28_port,
                           A(27) => MuxOutputs_6_27_port, A(26) => 
                           MuxOutputs_6_26_port, A(25) => MuxOutputs_6_25_port,
                           A(24) => MuxOutputs_6_24_port, A(23) => 
                           MuxOutputs_6_23_port, A(22) => MuxOutputs_6_22_port,
                           A(21) => MuxOutputs_6_21_port, A(20) => 
                           MuxOutputs_6_20_port, A(19) => MuxOutputs_6_19_port,
                           A(18) => MuxOutputs_6_18_port, A(17) => 
                           MuxOutputs_6_17_port, A(16) => MuxOutputs_6_16_port,
                           A(15) => MuxOutputs_6_15_port, A(14) => 
                           MuxOutputs_6_14_port, A(13) => MuxOutputs_6_13_port,
                           A(12) => MuxOutputs_6_12_port, A(11) => 
                           MuxOutputs_6_11_port, A(10) => MuxOutputs_6_10_port,
                           A(9) => MuxOutputs_6_9_port, A(8) => 
                           MuxOutputs_6_8_port, A(7) => MuxOutputs_6_7_port, 
                           A(6) => MuxOutputs_6_6_port, A(5) => 
                           MuxOutputs_6_5_port, A(4) => MuxOutputs_6_4_port, 
                           A(3) => MuxOutputs_6_3_port, A(2) => 
                           MuxOutputs_6_2_port, A(1) => MuxOutputs_6_1_port, 
                           A(0) => MuxOutputs_6_0_port, B(63) => 
                           SumOutputs_4_63_port, B(62) => SumOutputs_4_62_port,
                           B(61) => SumOutputs_4_61_port, B(60) => 
                           SumOutputs_4_60_port, B(59) => SumOutputs_4_59_port,
                           B(58) => SumOutputs_4_58_port, B(57) => 
                           SumOutputs_4_57_port, B(56) => SumOutputs_4_56_port,
                           B(55) => SumOutputs_4_55_port, B(54) => 
                           SumOutputs_4_54_port, B(53) => SumOutputs_4_53_port,
                           B(52) => SumOutputs_4_52_port, B(51) => 
                           SumOutputs_4_51_port, B(50) => SumOutputs_4_50_port,
                           B(49) => SumOutputs_4_49_port, B(48) => 
                           SumOutputs_4_48_port, B(47) => SumOutputs_4_47_port,
                           B(46) => SumOutputs_4_46_port, B(45) => 
                           SumOutputs_4_45_port, B(44) => SumOutputs_4_44_port,
                           B(43) => SumOutputs_4_43_port, B(42) => 
                           SumOutputs_4_42_port, B(41) => SumOutputs_4_41_port,
                           B(40) => SumOutputs_4_40_port, B(39) => 
                           SumOutputs_4_39_port, B(38) => SumOutputs_4_38_port,
                           B(37) => SumOutputs_4_37_port, B(36) => 
                           SumOutputs_4_36_port, B(35) => SumOutputs_4_35_port,
                           B(34) => SumOutputs_4_34_port, B(33) => 
                           SumOutputs_4_33_port, B(32) => SumOutputs_4_32_port,
                           B(31) => SumOutputs_4_31_port, B(30) => 
                           SumOutputs_4_30_port, B(29) => SumOutputs_4_29_port,
                           B(28) => SumOutputs_4_28_port, B(27) => 
                           SumOutputs_4_27_port, B(26) => SumOutputs_4_26_port,
                           B(25) => SumOutputs_4_25_port, B(24) => 
                           SumOutputs_4_24_port, B(23) => SumOutputs_4_23_port,
                           B(22) => SumOutputs_4_22_port, B(21) => 
                           SumOutputs_4_21_port, B(20) => SumOutputs_4_20_port,
                           B(19) => SumOutputs_4_19_port, B(18) => 
                           SumOutputs_4_18_port, B(17) => SumOutputs_4_17_port,
                           B(16) => SumOutputs_4_16_port, B(15) => 
                           SumOutputs_4_15_port, B(14) => SumOutputs_4_14_port,
                           B(13) => SumOutputs_4_13_port, B(12) => 
                           SumOutputs_4_12_port, B(11) => SumOutputs_4_11_port,
                           B(10) => SumOutputs_4_10_port, B(9) => 
                           SumOutputs_4_9_port, B(8) => SumOutputs_4_8_port, 
                           B(7) => SumOutputs_4_7_port, B(6) => 
                           SumOutputs_4_6_port, B(5) => SumOutputs_4_5_port, 
                           B(4) => SumOutputs_4_4_port, B(3) => 
                           SumOutputs_4_3_port, B(2) => SumOutputs_4_2_port, 
                           B(1) => SumOutputs_4_1_port, B(0) => 
                           SumOutputs_4_0_port, Ci => X_Logic0_port, S(63) => 
                           SumOutputs_5_63_port, S(62) => SumOutputs_5_62_port,
                           S(61) => SumOutputs_5_61_port, S(60) => 
                           SumOutputs_5_60_port, S(59) => SumOutputs_5_59_port,
                           S(58) => SumOutputs_5_58_port, S(57) => 
                           SumOutputs_5_57_port, S(56) => SumOutputs_5_56_port,
                           S(55) => SumOutputs_5_55_port, S(54) => 
                           SumOutputs_5_54_port, S(53) => SumOutputs_5_53_port,
                           S(52) => SumOutputs_5_52_port, S(51) => 
                           SumOutputs_5_51_port, S(50) => SumOutputs_5_50_port,
                           S(49) => SumOutputs_5_49_port, S(48) => 
                           SumOutputs_5_48_port, S(47) => SumOutputs_5_47_port,
                           S(46) => SumOutputs_5_46_port, S(45) => 
                           SumOutputs_5_45_port, S(44) => SumOutputs_5_44_port,
                           S(43) => SumOutputs_5_43_port, S(42) => 
                           SumOutputs_5_42_port, S(41) => SumOutputs_5_41_port,
                           S(40) => SumOutputs_5_40_port, S(39) => 
                           SumOutputs_5_39_port, S(38) => SumOutputs_5_38_port,
                           S(37) => SumOutputs_5_37_port, S(36) => 
                           SumOutputs_5_36_port, S(35) => SumOutputs_5_35_port,
                           S(34) => SumOutputs_5_34_port, S(33) => 
                           SumOutputs_5_33_port, S(32) => SumOutputs_5_32_port,
                           S(31) => SumOutputs_5_31_port, S(30) => 
                           SumOutputs_5_30_port, S(29) => SumOutputs_5_29_port,
                           S(28) => SumOutputs_5_28_port, S(27) => 
                           SumOutputs_5_27_port, S(26) => SumOutputs_5_26_port,
                           S(25) => SumOutputs_5_25_port, S(24) => 
                           SumOutputs_5_24_port, S(23) => SumOutputs_5_23_port,
                           S(22) => SumOutputs_5_22_port, S(21) => 
                           SumOutputs_5_21_port, S(20) => SumOutputs_5_20_port,
                           S(19) => SumOutputs_5_19_port, S(18) => 
                           SumOutputs_5_18_port, S(17) => SumOutputs_5_17_port,
                           S(16) => SumOutputs_5_16_port, S(15) => 
                           SumOutputs_5_15_port, S(14) => SumOutputs_5_14_port,
                           S(13) => SumOutputs_5_13_port, S(12) => 
                           SumOutputs_5_12_port, S(11) => SumOutputs_5_11_port,
                           S(10) => SumOutputs_5_10_port, S(9) => 
                           SumOutputs_5_9_port, S(8) => SumOutputs_5_8_port, 
                           S(7) => SumOutputs_5_7_port, S(6) => 
                           SumOutputs_5_6_port, S(5) => SumOutputs_5_5_port, 
                           S(4) => SumOutputs_5_4_port, S(3) => 
                           SumOutputs_5_3_port, S(2) => SumOutputs_5_2_port, 
                           S(1) => SumOutputs_5_1_port, S(0) => 
                           SumOutputs_5_0_port, Co => n_1132);
   SUMI_6 : RCA_NbitRca64_9 port map( A(63) => MuxOutputs_7_63_port, A(62) => 
                           MuxOutputs_7_62_port, A(61) => MuxOutputs_7_61_port,
                           A(60) => MuxOutputs_7_60_port, A(59) => 
                           MuxOutputs_7_59_port, A(58) => MuxOutputs_7_58_port,
                           A(57) => MuxOutputs_7_57_port, A(56) => 
                           MuxOutputs_7_56_port, A(55) => MuxOutputs_7_55_port,
                           A(54) => MuxOutputs_7_54_port, A(53) => 
                           MuxOutputs_7_53_port, A(52) => MuxOutputs_7_52_port,
                           A(51) => MuxOutputs_7_51_port, A(50) => 
                           MuxOutputs_7_50_port, A(49) => MuxOutputs_7_49_port,
                           A(48) => MuxOutputs_7_48_port, A(47) => 
                           MuxOutputs_7_47_port, A(46) => MuxOutputs_7_46_port,
                           A(45) => MuxOutputs_7_45_port, A(44) => 
                           MuxOutputs_7_44_port, A(43) => MuxOutputs_7_43_port,
                           A(42) => MuxOutputs_7_42_port, A(41) => 
                           MuxOutputs_7_41_port, A(40) => MuxOutputs_7_40_port,
                           A(39) => MuxOutputs_7_39_port, A(38) => 
                           MuxOutputs_7_38_port, A(37) => MuxOutputs_7_37_port,
                           A(36) => MuxOutputs_7_36_port, A(35) => 
                           MuxOutputs_7_35_port, A(34) => MuxOutputs_7_34_port,
                           A(33) => MuxOutputs_7_33_port, A(32) => 
                           MuxOutputs_7_32_port, A(31) => MuxOutputs_7_31_port,
                           A(30) => MuxOutputs_7_30_port, A(29) => 
                           MuxOutputs_7_29_port, A(28) => MuxOutputs_7_28_port,
                           A(27) => MuxOutputs_7_27_port, A(26) => 
                           MuxOutputs_7_26_port, A(25) => MuxOutputs_7_25_port,
                           A(24) => MuxOutputs_7_24_port, A(23) => 
                           MuxOutputs_7_23_port, A(22) => MuxOutputs_7_22_port,
                           A(21) => MuxOutputs_7_21_port, A(20) => 
                           MuxOutputs_7_20_port, A(19) => MuxOutputs_7_19_port,
                           A(18) => MuxOutputs_7_18_port, A(17) => 
                           MuxOutputs_7_17_port, A(16) => MuxOutputs_7_16_port,
                           A(15) => MuxOutputs_7_15_port, A(14) => 
                           MuxOutputs_7_14_port, A(13) => MuxOutputs_7_13_port,
                           A(12) => MuxOutputs_7_12_port, A(11) => 
                           MuxOutputs_7_11_port, A(10) => MuxOutputs_7_10_port,
                           A(9) => MuxOutputs_7_9_port, A(8) => 
                           MuxOutputs_7_8_port, A(7) => MuxOutputs_7_7_port, 
                           A(6) => MuxOutputs_7_6_port, A(5) => 
                           MuxOutputs_7_5_port, A(4) => MuxOutputs_7_4_port, 
                           A(3) => MuxOutputs_7_3_port, A(2) => 
                           MuxOutputs_7_2_port, A(1) => MuxOutputs_7_1_port, 
                           A(0) => MuxOutputs_7_0_port, B(63) => 
                           SumOutputs_5_63_port, B(62) => SumOutputs_5_62_port,
                           B(61) => SumOutputs_5_61_port, B(60) => 
                           SumOutputs_5_60_port, B(59) => SumOutputs_5_59_port,
                           B(58) => SumOutputs_5_58_port, B(57) => 
                           SumOutputs_5_57_port, B(56) => SumOutputs_5_56_port,
                           B(55) => SumOutputs_5_55_port, B(54) => 
                           SumOutputs_5_54_port, B(53) => SumOutputs_5_53_port,
                           B(52) => SumOutputs_5_52_port, B(51) => 
                           SumOutputs_5_51_port, B(50) => SumOutputs_5_50_port,
                           B(49) => SumOutputs_5_49_port, B(48) => 
                           SumOutputs_5_48_port, B(47) => SumOutputs_5_47_port,
                           B(46) => SumOutputs_5_46_port, B(45) => 
                           SumOutputs_5_45_port, B(44) => SumOutputs_5_44_port,
                           B(43) => SumOutputs_5_43_port, B(42) => 
                           SumOutputs_5_42_port, B(41) => SumOutputs_5_41_port,
                           B(40) => SumOutputs_5_40_port, B(39) => 
                           SumOutputs_5_39_port, B(38) => SumOutputs_5_38_port,
                           B(37) => SumOutputs_5_37_port, B(36) => 
                           SumOutputs_5_36_port, B(35) => SumOutputs_5_35_port,
                           B(34) => SumOutputs_5_34_port, B(33) => 
                           SumOutputs_5_33_port, B(32) => SumOutputs_5_32_port,
                           B(31) => SumOutputs_5_31_port, B(30) => 
                           SumOutputs_5_30_port, B(29) => SumOutputs_5_29_port,
                           B(28) => SumOutputs_5_28_port, B(27) => 
                           SumOutputs_5_27_port, B(26) => SumOutputs_5_26_port,
                           B(25) => SumOutputs_5_25_port, B(24) => 
                           SumOutputs_5_24_port, B(23) => SumOutputs_5_23_port,
                           B(22) => SumOutputs_5_22_port, B(21) => 
                           SumOutputs_5_21_port, B(20) => SumOutputs_5_20_port,
                           B(19) => SumOutputs_5_19_port, B(18) => 
                           SumOutputs_5_18_port, B(17) => SumOutputs_5_17_port,
                           B(16) => SumOutputs_5_16_port, B(15) => 
                           SumOutputs_5_15_port, B(14) => SumOutputs_5_14_port,
                           B(13) => SumOutputs_5_13_port, B(12) => 
                           SumOutputs_5_12_port, B(11) => SumOutputs_5_11_port,
                           B(10) => SumOutputs_5_10_port, B(9) => 
                           SumOutputs_5_9_port, B(8) => SumOutputs_5_8_port, 
                           B(7) => SumOutputs_5_7_port, B(6) => 
                           SumOutputs_5_6_port, B(5) => SumOutputs_5_5_port, 
                           B(4) => SumOutputs_5_4_port, B(3) => 
                           SumOutputs_5_3_port, B(2) => SumOutputs_5_2_port, 
                           B(1) => SumOutputs_5_1_port, B(0) => 
                           SumOutputs_5_0_port, Ci => X_Logic0_port, S(63) => 
                           SumOutputs_6_63_port, S(62) => SumOutputs_6_62_port,
                           S(61) => SumOutputs_6_61_port, S(60) => 
                           SumOutputs_6_60_port, S(59) => SumOutputs_6_59_port,
                           S(58) => SumOutputs_6_58_port, S(57) => 
                           SumOutputs_6_57_port, S(56) => SumOutputs_6_56_port,
                           S(55) => SumOutputs_6_55_port, S(54) => 
                           SumOutputs_6_54_port, S(53) => SumOutputs_6_53_port,
                           S(52) => SumOutputs_6_52_port, S(51) => 
                           SumOutputs_6_51_port, S(50) => SumOutputs_6_50_port,
                           S(49) => SumOutputs_6_49_port, S(48) => 
                           SumOutputs_6_48_port, S(47) => SumOutputs_6_47_port,
                           S(46) => SumOutputs_6_46_port, S(45) => 
                           SumOutputs_6_45_port, S(44) => SumOutputs_6_44_port,
                           S(43) => SumOutputs_6_43_port, S(42) => 
                           SumOutputs_6_42_port, S(41) => SumOutputs_6_41_port,
                           S(40) => SumOutputs_6_40_port, S(39) => 
                           SumOutputs_6_39_port, S(38) => SumOutputs_6_38_port,
                           S(37) => SumOutputs_6_37_port, S(36) => 
                           SumOutputs_6_36_port, S(35) => SumOutputs_6_35_port,
                           S(34) => SumOutputs_6_34_port, S(33) => 
                           SumOutputs_6_33_port, S(32) => SumOutputs_6_32_port,
                           S(31) => SumOutputs_6_31_port, S(30) => 
                           SumOutputs_6_30_port, S(29) => SumOutputs_6_29_port,
                           S(28) => SumOutputs_6_28_port, S(27) => 
                           SumOutputs_6_27_port, S(26) => SumOutputs_6_26_port,
                           S(25) => SumOutputs_6_25_port, S(24) => 
                           SumOutputs_6_24_port, S(23) => SumOutputs_6_23_port,
                           S(22) => SumOutputs_6_22_port, S(21) => 
                           SumOutputs_6_21_port, S(20) => SumOutputs_6_20_port,
                           S(19) => SumOutputs_6_19_port, S(18) => 
                           SumOutputs_6_18_port, S(17) => SumOutputs_6_17_port,
                           S(16) => SumOutputs_6_16_port, S(15) => 
                           SumOutputs_6_15_port, S(14) => SumOutputs_6_14_port,
                           S(13) => SumOutputs_6_13_port, S(12) => 
                           SumOutputs_6_12_port, S(11) => SumOutputs_6_11_port,
                           S(10) => SumOutputs_6_10_port, S(9) => 
                           SumOutputs_6_9_port, S(8) => SumOutputs_6_8_port, 
                           S(7) => SumOutputs_6_7_port, S(6) => 
                           SumOutputs_6_6_port, S(5) => SumOutputs_6_5_port, 
                           S(4) => SumOutputs_6_4_port, S(3) => 
                           SumOutputs_6_3_port, S(2) => SumOutputs_6_2_port, 
                           S(1) => SumOutputs_6_1_port, S(0) => 
                           SumOutputs_6_0_port, Co => n_1133);
   SUMI_7 : RCA_NbitRca64_8 port map( A(63) => MuxOutputs_8_63_port, A(62) => 
                           MuxOutputs_8_62_port, A(61) => MuxOutputs_8_61_port,
                           A(60) => MuxOutputs_8_60_port, A(59) => 
                           MuxOutputs_8_59_port, A(58) => MuxOutputs_8_58_port,
                           A(57) => MuxOutputs_8_57_port, A(56) => 
                           MuxOutputs_8_56_port, A(55) => MuxOutputs_8_55_port,
                           A(54) => MuxOutputs_8_54_port, A(53) => 
                           MuxOutputs_8_53_port, A(52) => MuxOutputs_8_52_port,
                           A(51) => MuxOutputs_8_51_port, A(50) => 
                           MuxOutputs_8_50_port, A(49) => MuxOutputs_8_49_port,
                           A(48) => MuxOutputs_8_48_port, A(47) => 
                           MuxOutputs_8_47_port, A(46) => MuxOutputs_8_46_port,
                           A(45) => MuxOutputs_8_45_port, A(44) => 
                           MuxOutputs_8_44_port, A(43) => MuxOutputs_8_43_port,
                           A(42) => MuxOutputs_8_42_port, A(41) => 
                           MuxOutputs_8_41_port, A(40) => MuxOutputs_8_40_port,
                           A(39) => MuxOutputs_8_39_port, A(38) => 
                           MuxOutputs_8_38_port, A(37) => MuxOutputs_8_37_port,
                           A(36) => MuxOutputs_8_36_port, A(35) => 
                           MuxOutputs_8_35_port, A(34) => MuxOutputs_8_34_port,
                           A(33) => MuxOutputs_8_33_port, A(32) => 
                           MuxOutputs_8_32_port, A(31) => MuxOutputs_8_31_port,
                           A(30) => MuxOutputs_8_30_port, A(29) => 
                           MuxOutputs_8_29_port, A(28) => MuxOutputs_8_28_port,
                           A(27) => MuxOutputs_8_27_port, A(26) => 
                           MuxOutputs_8_26_port, A(25) => MuxOutputs_8_25_port,
                           A(24) => MuxOutputs_8_24_port, A(23) => 
                           MuxOutputs_8_23_port, A(22) => MuxOutputs_8_22_port,
                           A(21) => MuxOutputs_8_21_port, A(20) => 
                           MuxOutputs_8_20_port, A(19) => MuxOutputs_8_19_port,
                           A(18) => MuxOutputs_8_18_port, A(17) => 
                           MuxOutputs_8_17_port, A(16) => MuxOutputs_8_16_port,
                           A(15) => MuxOutputs_8_15_port, A(14) => 
                           MuxOutputs_8_14_port, A(13) => MuxOutputs_8_13_port,
                           A(12) => MuxOutputs_8_12_port, A(11) => 
                           MuxOutputs_8_11_port, A(10) => MuxOutputs_8_10_port,
                           A(9) => MuxOutputs_8_9_port, A(8) => 
                           MuxOutputs_8_8_port, A(7) => MuxOutputs_8_7_port, 
                           A(6) => MuxOutputs_8_6_port, A(5) => 
                           MuxOutputs_8_5_port, A(4) => MuxOutputs_8_4_port, 
                           A(3) => MuxOutputs_8_3_port, A(2) => 
                           MuxOutputs_8_2_port, A(1) => MuxOutputs_8_1_port, 
                           A(0) => MuxOutputs_8_0_port, B(63) => 
                           SumOutputs_6_63_port, B(62) => SumOutputs_6_62_port,
                           B(61) => SumOutputs_6_61_port, B(60) => 
                           SumOutputs_6_60_port, B(59) => SumOutputs_6_59_port,
                           B(58) => SumOutputs_6_58_port, B(57) => 
                           SumOutputs_6_57_port, B(56) => SumOutputs_6_56_port,
                           B(55) => SumOutputs_6_55_port, B(54) => 
                           SumOutputs_6_54_port, B(53) => SumOutputs_6_53_port,
                           B(52) => SumOutputs_6_52_port, B(51) => 
                           SumOutputs_6_51_port, B(50) => SumOutputs_6_50_port,
                           B(49) => SumOutputs_6_49_port, B(48) => 
                           SumOutputs_6_48_port, B(47) => SumOutputs_6_47_port,
                           B(46) => SumOutputs_6_46_port, B(45) => 
                           SumOutputs_6_45_port, B(44) => SumOutputs_6_44_port,
                           B(43) => SumOutputs_6_43_port, B(42) => 
                           SumOutputs_6_42_port, B(41) => SumOutputs_6_41_port,
                           B(40) => SumOutputs_6_40_port, B(39) => 
                           SumOutputs_6_39_port, B(38) => SumOutputs_6_38_port,
                           B(37) => SumOutputs_6_37_port, B(36) => 
                           SumOutputs_6_36_port, B(35) => SumOutputs_6_35_port,
                           B(34) => SumOutputs_6_34_port, B(33) => 
                           SumOutputs_6_33_port, B(32) => SumOutputs_6_32_port,
                           B(31) => SumOutputs_6_31_port, B(30) => 
                           SumOutputs_6_30_port, B(29) => SumOutputs_6_29_port,
                           B(28) => SumOutputs_6_28_port, B(27) => 
                           SumOutputs_6_27_port, B(26) => SumOutputs_6_26_port,
                           B(25) => SumOutputs_6_25_port, B(24) => 
                           SumOutputs_6_24_port, B(23) => SumOutputs_6_23_port,
                           B(22) => SumOutputs_6_22_port, B(21) => 
                           SumOutputs_6_21_port, B(20) => SumOutputs_6_20_port,
                           B(19) => SumOutputs_6_19_port, B(18) => 
                           SumOutputs_6_18_port, B(17) => SumOutputs_6_17_port,
                           B(16) => SumOutputs_6_16_port, B(15) => 
                           SumOutputs_6_15_port, B(14) => SumOutputs_6_14_port,
                           B(13) => SumOutputs_6_13_port, B(12) => 
                           SumOutputs_6_12_port, B(11) => SumOutputs_6_11_port,
                           B(10) => SumOutputs_6_10_port, B(9) => 
                           SumOutputs_6_9_port, B(8) => SumOutputs_6_8_port, 
                           B(7) => SumOutputs_6_7_port, B(6) => 
                           SumOutputs_6_6_port, B(5) => SumOutputs_6_5_port, 
                           B(4) => SumOutputs_6_4_port, B(3) => 
                           SumOutputs_6_3_port, B(2) => SumOutputs_6_2_port, 
                           B(1) => SumOutputs_6_1_port, B(0) => 
                           SumOutputs_6_0_port, Ci => X_Logic0_port, S(63) => 
                           SumOutputs_7_63_port, S(62) => SumOutputs_7_62_port,
                           S(61) => SumOutputs_7_61_port, S(60) => 
                           SumOutputs_7_60_port, S(59) => SumOutputs_7_59_port,
                           S(58) => SumOutputs_7_58_port, S(57) => 
                           SumOutputs_7_57_port, S(56) => SumOutputs_7_56_port,
                           S(55) => SumOutputs_7_55_port, S(54) => 
                           SumOutputs_7_54_port, S(53) => SumOutputs_7_53_port,
                           S(52) => SumOutputs_7_52_port, S(51) => 
                           SumOutputs_7_51_port, S(50) => SumOutputs_7_50_port,
                           S(49) => SumOutputs_7_49_port, S(48) => 
                           SumOutputs_7_48_port, S(47) => SumOutputs_7_47_port,
                           S(46) => SumOutputs_7_46_port, S(45) => 
                           SumOutputs_7_45_port, S(44) => SumOutputs_7_44_port,
                           S(43) => SumOutputs_7_43_port, S(42) => 
                           SumOutputs_7_42_port, S(41) => SumOutputs_7_41_port,
                           S(40) => SumOutputs_7_40_port, S(39) => 
                           SumOutputs_7_39_port, S(38) => SumOutputs_7_38_port,
                           S(37) => SumOutputs_7_37_port, S(36) => 
                           SumOutputs_7_36_port, S(35) => SumOutputs_7_35_port,
                           S(34) => SumOutputs_7_34_port, S(33) => 
                           SumOutputs_7_33_port, S(32) => SumOutputs_7_32_port,
                           S(31) => SumOutputs_7_31_port, S(30) => 
                           SumOutputs_7_30_port, S(29) => SumOutputs_7_29_port,
                           S(28) => SumOutputs_7_28_port, S(27) => 
                           SumOutputs_7_27_port, S(26) => SumOutputs_7_26_port,
                           S(25) => SumOutputs_7_25_port, S(24) => 
                           SumOutputs_7_24_port, S(23) => SumOutputs_7_23_port,
                           S(22) => SumOutputs_7_22_port, S(21) => 
                           SumOutputs_7_21_port, S(20) => SumOutputs_7_20_port,
                           S(19) => SumOutputs_7_19_port, S(18) => 
                           SumOutputs_7_18_port, S(17) => SumOutputs_7_17_port,
                           S(16) => SumOutputs_7_16_port, S(15) => 
                           SumOutputs_7_15_port, S(14) => SumOutputs_7_14_port,
                           S(13) => SumOutputs_7_13_port, S(12) => 
                           SumOutputs_7_12_port, S(11) => SumOutputs_7_11_port,
                           S(10) => SumOutputs_7_10_port, S(9) => 
                           SumOutputs_7_9_port, S(8) => SumOutputs_7_8_port, 
                           S(7) => SumOutputs_7_7_port, S(6) => 
                           SumOutputs_7_6_port, S(5) => SumOutputs_7_5_port, 
                           S(4) => SumOutputs_7_4_port, S(3) => 
                           SumOutputs_7_3_port, S(2) => SumOutputs_7_2_port, 
                           S(1) => SumOutputs_7_1_port, S(0) => 
                           SumOutputs_7_0_port, Co => n_1134);
   SUMI_8 : RCA_NbitRca64_7 port map( A(63) => MuxOutputs_9_63_port, A(62) => 
                           MuxOutputs_9_62_port, A(61) => MuxOutputs_9_61_port,
                           A(60) => MuxOutputs_9_60_port, A(59) => 
                           MuxOutputs_9_59_port, A(58) => MuxOutputs_9_58_port,
                           A(57) => MuxOutputs_9_57_port, A(56) => 
                           MuxOutputs_9_56_port, A(55) => MuxOutputs_9_55_port,
                           A(54) => MuxOutputs_9_54_port, A(53) => 
                           MuxOutputs_9_53_port, A(52) => MuxOutputs_9_52_port,
                           A(51) => MuxOutputs_9_51_port, A(50) => 
                           MuxOutputs_9_50_port, A(49) => MuxOutputs_9_49_port,
                           A(48) => MuxOutputs_9_48_port, A(47) => 
                           MuxOutputs_9_47_port, A(46) => MuxOutputs_9_46_port,
                           A(45) => MuxOutputs_9_45_port, A(44) => 
                           MuxOutputs_9_44_port, A(43) => MuxOutputs_9_43_port,
                           A(42) => MuxOutputs_9_42_port, A(41) => 
                           MuxOutputs_9_41_port, A(40) => MuxOutputs_9_40_port,
                           A(39) => MuxOutputs_9_39_port, A(38) => 
                           MuxOutputs_9_38_port, A(37) => MuxOutputs_9_37_port,
                           A(36) => MuxOutputs_9_36_port, A(35) => 
                           MuxOutputs_9_35_port, A(34) => MuxOutputs_9_34_port,
                           A(33) => MuxOutputs_9_33_port, A(32) => 
                           MuxOutputs_9_32_port, A(31) => MuxOutputs_9_31_port,
                           A(30) => MuxOutputs_9_30_port, A(29) => 
                           MuxOutputs_9_29_port, A(28) => MuxOutputs_9_28_port,
                           A(27) => MuxOutputs_9_27_port, A(26) => 
                           MuxOutputs_9_26_port, A(25) => MuxOutputs_9_25_port,
                           A(24) => MuxOutputs_9_24_port, A(23) => 
                           MuxOutputs_9_23_port, A(22) => MuxOutputs_9_22_port,
                           A(21) => MuxOutputs_9_21_port, A(20) => 
                           MuxOutputs_9_20_port, A(19) => MuxOutputs_9_19_port,
                           A(18) => MuxOutputs_9_18_port, A(17) => 
                           MuxOutputs_9_17_port, A(16) => MuxOutputs_9_16_port,
                           A(15) => MuxOutputs_9_15_port, A(14) => 
                           MuxOutputs_9_14_port, A(13) => MuxOutputs_9_13_port,
                           A(12) => MuxOutputs_9_12_port, A(11) => 
                           MuxOutputs_9_11_port, A(10) => MuxOutputs_9_10_port,
                           A(9) => MuxOutputs_9_9_port, A(8) => 
                           MuxOutputs_9_8_port, A(7) => MuxOutputs_9_7_port, 
                           A(6) => MuxOutputs_9_6_port, A(5) => 
                           MuxOutputs_9_5_port, A(4) => MuxOutputs_9_4_port, 
                           A(3) => MuxOutputs_9_3_port, A(2) => 
                           MuxOutputs_9_2_port, A(1) => MuxOutputs_9_1_port, 
                           A(0) => MuxOutputs_9_0_port, B(63) => 
                           SumOutputs_7_63_port, B(62) => SumOutputs_7_62_port,
                           B(61) => SumOutputs_7_61_port, B(60) => 
                           SumOutputs_7_60_port, B(59) => SumOutputs_7_59_port,
                           B(58) => SumOutputs_7_58_port, B(57) => 
                           SumOutputs_7_57_port, B(56) => SumOutputs_7_56_port,
                           B(55) => SumOutputs_7_55_port, B(54) => 
                           SumOutputs_7_54_port, B(53) => SumOutputs_7_53_port,
                           B(52) => SumOutputs_7_52_port, B(51) => 
                           SumOutputs_7_51_port, B(50) => SumOutputs_7_50_port,
                           B(49) => SumOutputs_7_49_port, B(48) => 
                           SumOutputs_7_48_port, B(47) => SumOutputs_7_47_port,
                           B(46) => SumOutputs_7_46_port, B(45) => 
                           SumOutputs_7_45_port, B(44) => SumOutputs_7_44_port,
                           B(43) => SumOutputs_7_43_port, B(42) => 
                           SumOutputs_7_42_port, B(41) => SumOutputs_7_41_port,
                           B(40) => SumOutputs_7_40_port, B(39) => 
                           SumOutputs_7_39_port, B(38) => SumOutputs_7_38_port,
                           B(37) => SumOutputs_7_37_port, B(36) => 
                           SumOutputs_7_36_port, B(35) => SumOutputs_7_35_port,
                           B(34) => SumOutputs_7_34_port, B(33) => 
                           SumOutputs_7_33_port, B(32) => SumOutputs_7_32_port,
                           B(31) => SumOutputs_7_31_port, B(30) => 
                           SumOutputs_7_30_port, B(29) => SumOutputs_7_29_port,
                           B(28) => SumOutputs_7_28_port, B(27) => 
                           SumOutputs_7_27_port, B(26) => SumOutputs_7_26_port,
                           B(25) => SumOutputs_7_25_port, B(24) => 
                           SumOutputs_7_24_port, B(23) => SumOutputs_7_23_port,
                           B(22) => SumOutputs_7_22_port, B(21) => 
                           SumOutputs_7_21_port, B(20) => SumOutputs_7_20_port,
                           B(19) => SumOutputs_7_19_port, B(18) => 
                           SumOutputs_7_18_port, B(17) => SumOutputs_7_17_port,
                           B(16) => SumOutputs_7_16_port, B(15) => 
                           SumOutputs_7_15_port, B(14) => SumOutputs_7_14_port,
                           B(13) => SumOutputs_7_13_port, B(12) => 
                           SumOutputs_7_12_port, B(11) => SumOutputs_7_11_port,
                           B(10) => SumOutputs_7_10_port, B(9) => 
                           SumOutputs_7_9_port, B(8) => SumOutputs_7_8_port, 
                           B(7) => SumOutputs_7_7_port, B(6) => 
                           SumOutputs_7_6_port, B(5) => SumOutputs_7_5_port, 
                           B(4) => SumOutputs_7_4_port, B(3) => 
                           SumOutputs_7_3_port, B(2) => SumOutputs_7_2_port, 
                           B(1) => SumOutputs_7_1_port, B(0) => 
                           SumOutputs_7_0_port, Ci => X_Logic0_port, S(63) => 
                           SumOutputs_8_63_port, S(62) => SumOutputs_8_62_port,
                           S(61) => SumOutputs_8_61_port, S(60) => 
                           SumOutputs_8_60_port, S(59) => SumOutputs_8_59_port,
                           S(58) => SumOutputs_8_58_port, S(57) => 
                           SumOutputs_8_57_port, S(56) => SumOutputs_8_56_port,
                           S(55) => SumOutputs_8_55_port, S(54) => 
                           SumOutputs_8_54_port, S(53) => SumOutputs_8_53_port,
                           S(52) => SumOutputs_8_52_port, S(51) => 
                           SumOutputs_8_51_port, S(50) => SumOutputs_8_50_port,
                           S(49) => SumOutputs_8_49_port, S(48) => 
                           SumOutputs_8_48_port, S(47) => SumOutputs_8_47_port,
                           S(46) => SumOutputs_8_46_port, S(45) => 
                           SumOutputs_8_45_port, S(44) => SumOutputs_8_44_port,
                           S(43) => SumOutputs_8_43_port, S(42) => 
                           SumOutputs_8_42_port, S(41) => SumOutputs_8_41_port,
                           S(40) => SumOutputs_8_40_port, S(39) => 
                           SumOutputs_8_39_port, S(38) => SumOutputs_8_38_port,
                           S(37) => SumOutputs_8_37_port, S(36) => 
                           SumOutputs_8_36_port, S(35) => SumOutputs_8_35_port,
                           S(34) => SumOutputs_8_34_port, S(33) => 
                           SumOutputs_8_33_port, S(32) => SumOutputs_8_32_port,
                           S(31) => SumOutputs_8_31_port, S(30) => 
                           SumOutputs_8_30_port, S(29) => SumOutputs_8_29_port,
                           S(28) => SumOutputs_8_28_port, S(27) => 
                           SumOutputs_8_27_port, S(26) => SumOutputs_8_26_port,
                           S(25) => SumOutputs_8_25_port, S(24) => 
                           SumOutputs_8_24_port, S(23) => SumOutputs_8_23_port,
                           S(22) => SumOutputs_8_22_port, S(21) => 
                           SumOutputs_8_21_port, S(20) => SumOutputs_8_20_port,
                           S(19) => SumOutputs_8_19_port, S(18) => 
                           SumOutputs_8_18_port, S(17) => SumOutputs_8_17_port,
                           S(16) => SumOutputs_8_16_port, S(15) => 
                           SumOutputs_8_15_port, S(14) => SumOutputs_8_14_port,
                           S(13) => SumOutputs_8_13_port, S(12) => 
                           SumOutputs_8_12_port, S(11) => SumOutputs_8_11_port,
                           S(10) => SumOutputs_8_10_port, S(9) => 
                           SumOutputs_8_9_port, S(8) => SumOutputs_8_8_port, 
                           S(7) => SumOutputs_8_7_port, S(6) => 
                           SumOutputs_8_6_port, S(5) => SumOutputs_8_5_port, 
                           S(4) => SumOutputs_8_4_port, S(3) => 
                           SumOutputs_8_3_port, S(2) => SumOutputs_8_2_port, 
                           S(1) => SumOutputs_8_1_port, S(0) => 
                           SumOutputs_8_0_port, Co => n_1135);
   SUMI_9 : RCA_NbitRca64_6 port map( A(63) => MuxOutputs_10_63_port, A(62) => 
                           MuxOutputs_10_62_port, A(61) => 
                           MuxOutputs_10_61_port, A(60) => 
                           MuxOutputs_10_60_port, A(59) => 
                           MuxOutputs_10_59_port, A(58) => 
                           MuxOutputs_10_58_port, A(57) => 
                           MuxOutputs_10_57_port, A(56) => 
                           MuxOutputs_10_56_port, A(55) => 
                           MuxOutputs_10_55_port, A(54) => 
                           MuxOutputs_10_54_port, A(53) => 
                           MuxOutputs_10_53_port, A(52) => 
                           MuxOutputs_10_52_port, A(51) => 
                           MuxOutputs_10_51_port, A(50) => 
                           MuxOutputs_10_50_port, A(49) => 
                           MuxOutputs_10_49_port, A(48) => 
                           MuxOutputs_10_48_port, A(47) => 
                           MuxOutputs_10_47_port, A(46) => 
                           MuxOutputs_10_46_port, A(45) => 
                           MuxOutputs_10_45_port, A(44) => 
                           MuxOutputs_10_44_port, A(43) => 
                           MuxOutputs_10_43_port, A(42) => 
                           MuxOutputs_10_42_port, A(41) => 
                           MuxOutputs_10_41_port, A(40) => 
                           MuxOutputs_10_40_port, A(39) => 
                           MuxOutputs_10_39_port, A(38) => 
                           MuxOutputs_10_38_port, A(37) => 
                           MuxOutputs_10_37_port, A(36) => 
                           MuxOutputs_10_36_port, A(35) => 
                           MuxOutputs_10_35_port, A(34) => 
                           MuxOutputs_10_34_port, A(33) => 
                           MuxOutputs_10_33_port, A(32) => 
                           MuxOutputs_10_32_port, A(31) => 
                           MuxOutputs_10_31_port, A(30) => 
                           MuxOutputs_10_30_port, A(29) => 
                           MuxOutputs_10_29_port, A(28) => 
                           MuxOutputs_10_28_port, A(27) => 
                           MuxOutputs_10_27_port, A(26) => 
                           MuxOutputs_10_26_port, A(25) => 
                           MuxOutputs_10_25_port, A(24) => 
                           MuxOutputs_10_24_port, A(23) => 
                           MuxOutputs_10_23_port, A(22) => 
                           MuxOutputs_10_22_port, A(21) => 
                           MuxOutputs_10_21_port, A(20) => 
                           MuxOutputs_10_20_port, A(19) => 
                           MuxOutputs_10_19_port, A(18) => 
                           MuxOutputs_10_18_port, A(17) => 
                           MuxOutputs_10_17_port, A(16) => 
                           MuxOutputs_10_16_port, A(15) => 
                           MuxOutputs_10_15_port, A(14) => 
                           MuxOutputs_10_14_port, A(13) => 
                           MuxOutputs_10_13_port, A(12) => 
                           MuxOutputs_10_12_port, A(11) => 
                           MuxOutputs_10_11_port, A(10) => 
                           MuxOutputs_10_10_port, A(9) => MuxOutputs_10_9_port,
                           A(8) => MuxOutputs_10_8_port, A(7) => 
                           MuxOutputs_10_7_port, A(6) => MuxOutputs_10_6_port, 
                           A(5) => MuxOutputs_10_5_port, A(4) => 
                           MuxOutputs_10_4_port, A(3) => MuxOutputs_10_3_port, 
                           A(2) => MuxOutputs_10_2_port, A(1) => 
                           MuxOutputs_10_1_port, A(0) => MuxOutputs_10_0_port, 
                           B(63) => SumOutputs_8_63_port, B(62) => 
                           SumOutputs_8_62_port, B(61) => SumOutputs_8_61_port,
                           B(60) => SumOutputs_8_60_port, B(59) => 
                           SumOutputs_8_59_port, B(58) => SumOutputs_8_58_port,
                           B(57) => SumOutputs_8_57_port, B(56) => 
                           SumOutputs_8_56_port, B(55) => SumOutputs_8_55_port,
                           B(54) => SumOutputs_8_54_port, B(53) => 
                           SumOutputs_8_53_port, B(52) => SumOutputs_8_52_port,
                           B(51) => SumOutputs_8_51_port, B(50) => 
                           SumOutputs_8_50_port, B(49) => SumOutputs_8_49_port,
                           B(48) => SumOutputs_8_48_port, B(47) => 
                           SumOutputs_8_47_port, B(46) => SumOutputs_8_46_port,
                           B(45) => SumOutputs_8_45_port, B(44) => 
                           SumOutputs_8_44_port, B(43) => SumOutputs_8_43_port,
                           B(42) => SumOutputs_8_42_port, B(41) => 
                           SumOutputs_8_41_port, B(40) => SumOutputs_8_40_port,
                           B(39) => SumOutputs_8_39_port, B(38) => 
                           SumOutputs_8_38_port, B(37) => SumOutputs_8_37_port,
                           B(36) => SumOutputs_8_36_port, B(35) => 
                           SumOutputs_8_35_port, B(34) => SumOutputs_8_34_port,
                           B(33) => SumOutputs_8_33_port, B(32) => 
                           SumOutputs_8_32_port, B(31) => SumOutputs_8_31_port,
                           B(30) => SumOutputs_8_30_port, B(29) => 
                           SumOutputs_8_29_port, B(28) => SumOutputs_8_28_port,
                           B(27) => SumOutputs_8_27_port, B(26) => 
                           SumOutputs_8_26_port, B(25) => SumOutputs_8_25_port,
                           B(24) => SumOutputs_8_24_port, B(23) => 
                           SumOutputs_8_23_port, B(22) => SumOutputs_8_22_port,
                           B(21) => SumOutputs_8_21_port, B(20) => 
                           SumOutputs_8_20_port, B(19) => SumOutputs_8_19_port,
                           B(18) => SumOutputs_8_18_port, B(17) => 
                           SumOutputs_8_17_port, B(16) => SumOutputs_8_16_port,
                           B(15) => SumOutputs_8_15_port, B(14) => 
                           SumOutputs_8_14_port, B(13) => SumOutputs_8_13_port,
                           B(12) => SumOutputs_8_12_port, B(11) => 
                           SumOutputs_8_11_port, B(10) => SumOutputs_8_10_port,
                           B(9) => SumOutputs_8_9_port, B(8) => 
                           SumOutputs_8_8_port, B(7) => SumOutputs_8_7_port, 
                           B(6) => SumOutputs_8_6_port, B(5) => 
                           SumOutputs_8_5_port, B(4) => SumOutputs_8_4_port, 
                           B(3) => SumOutputs_8_3_port, B(2) => 
                           SumOutputs_8_2_port, B(1) => SumOutputs_8_1_port, 
                           B(0) => SumOutputs_8_0_port, Ci => X_Logic0_port, 
                           S(63) => SumOutputs_9_63_port, S(62) => 
                           SumOutputs_9_62_port, S(61) => SumOutputs_9_61_port,
                           S(60) => SumOutputs_9_60_port, S(59) => 
                           SumOutputs_9_59_port, S(58) => SumOutputs_9_58_port,
                           S(57) => SumOutputs_9_57_port, S(56) => 
                           SumOutputs_9_56_port, S(55) => SumOutputs_9_55_port,
                           S(54) => SumOutputs_9_54_port, S(53) => 
                           SumOutputs_9_53_port, S(52) => SumOutputs_9_52_port,
                           S(51) => SumOutputs_9_51_port, S(50) => 
                           SumOutputs_9_50_port, S(49) => SumOutputs_9_49_port,
                           S(48) => SumOutputs_9_48_port, S(47) => 
                           SumOutputs_9_47_port, S(46) => SumOutputs_9_46_port,
                           S(45) => SumOutputs_9_45_port, S(44) => 
                           SumOutputs_9_44_port, S(43) => SumOutputs_9_43_port,
                           S(42) => SumOutputs_9_42_port, S(41) => 
                           SumOutputs_9_41_port, S(40) => SumOutputs_9_40_port,
                           S(39) => SumOutputs_9_39_port, S(38) => 
                           SumOutputs_9_38_port, S(37) => SumOutputs_9_37_port,
                           S(36) => SumOutputs_9_36_port, S(35) => 
                           SumOutputs_9_35_port, S(34) => SumOutputs_9_34_port,
                           S(33) => SumOutputs_9_33_port, S(32) => 
                           SumOutputs_9_32_port, S(31) => SumOutputs_9_31_port,
                           S(30) => SumOutputs_9_30_port, S(29) => 
                           SumOutputs_9_29_port, S(28) => SumOutputs_9_28_port,
                           S(27) => SumOutputs_9_27_port, S(26) => 
                           SumOutputs_9_26_port, S(25) => SumOutputs_9_25_port,
                           S(24) => SumOutputs_9_24_port, S(23) => 
                           SumOutputs_9_23_port, S(22) => SumOutputs_9_22_port,
                           S(21) => SumOutputs_9_21_port, S(20) => 
                           SumOutputs_9_20_port, S(19) => SumOutputs_9_19_port,
                           S(18) => SumOutputs_9_18_port, S(17) => 
                           SumOutputs_9_17_port, S(16) => SumOutputs_9_16_port,
                           S(15) => SumOutputs_9_15_port, S(14) => 
                           SumOutputs_9_14_port, S(13) => SumOutputs_9_13_port,
                           S(12) => SumOutputs_9_12_port, S(11) => 
                           SumOutputs_9_11_port, S(10) => SumOutputs_9_10_port,
                           S(9) => SumOutputs_9_9_port, S(8) => 
                           SumOutputs_9_8_port, S(7) => SumOutputs_9_7_port, 
                           S(6) => SumOutputs_9_6_port, S(5) => 
                           SumOutputs_9_5_port, S(4) => SumOutputs_9_4_port, 
                           S(3) => SumOutputs_9_3_port, S(2) => 
                           SumOutputs_9_2_port, S(1) => SumOutputs_9_1_port, 
                           S(0) => SumOutputs_9_0_port, Co => n_1136);
   SUMI_10 : RCA_NbitRca64_5 port map( A(63) => MuxOutputs_11_63_port, A(62) =>
                           MuxOutputs_11_62_port, A(61) => 
                           MuxOutputs_11_61_port, A(60) => 
                           MuxOutputs_11_60_port, A(59) => 
                           MuxOutputs_11_59_port, A(58) => 
                           MuxOutputs_11_58_port, A(57) => 
                           MuxOutputs_11_57_port, A(56) => 
                           MuxOutputs_11_56_port, A(55) => 
                           MuxOutputs_11_55_port, A(54) => 
                           MuxOutputs_11_54_port, A(53) => 
                           MuxOutputs_11_53_port, A(52) => 
                           MuxOutputs_11_52_port, A(51) => 
                           MuxOutputs_11_51_port, A(50) => 
                           MuxOutputs_11_50_port, A(49) => 
                           MuxOutputs_11_49_port, A(48) => 
                           MuxOutputs_11_48_port, A(47) => 
                           MuxOutputs_11_47_port, A(46) => 
                           MuxOutputs_11_46_port, A(45) => 
                           MuxOutputs_11_45_port, A(44) => 
                           MuxOutputs_11_44_port, A(43) => 
                           MuxOutputs_11_43_port, A(42) => 
                           MuxOutputs_11_42_port, A(41) => 
                           MuxOutputs_11_41_port, A(40) => 
                           MuxOutputs_11_40_port, A(39) => 
                           MuxOutputs_11_39_port, A(38) => 
                           MuxOutputs_11_38_port, A(37) => 
                           MuxOutputs_11_37_port, A(36) => 
                           MuxOutputs_11_36_port, A(35) => 
                           MuxOutputs_11_35_port, A(34) => 
                           MuxOutputs_11_34_port, A(33) => 
                           MuxOutputs_11_33_port, A(32) => 
                           MuxOutputs_11_32_port, A(31) => 
                           MuxOutputs_11_31_port, A(30) => 
                           MuxOutputs_11_30_port, A(29) => 
                           MuxOutputs_11_29_port, A(28) => 
                           MuxOutputs_11_28_port, A(27) => 
                           MuxOutputs_11_27_port, A(26) => 
                           MuxOutputs_11_26_port, A(25) => 
                           MuxOutputs_11_25_port, A(24) => 
                           MuxOutputs_11_24_port, A(23) => 
                           MuxOutputs_11_23_port, A(22) => 
                           MuxOutputs_11_22_port, A(21) => 
                           MuxOutputs_11_21_port, A(20) => 
                           MuxOutputs_11_20_port, A(19) => 
                           MuxOutputs_11_19_port, A(18) => 
                           MuxOutputs_11_18_port, A(17) => 
                           MuxOutputs_11_17_port, A(16) => 
                           MuxOutputs_11_16_port, A(15) => 
                           MuxOutputs_11_15_port, A(14) => 
                           MuxOutputs_11_14_port, A(13) => 
                           MuxOutputs_11_13_port, A(12) => 
                           MuxOutputs_11_12_port, A(11) => 
                           MuxOutputs_11_11_port, A(10) => 
                           MuxOutputs_11_10_port, A(9) => MuxOutputs_11_9_port,
                           A(8) => MuxOutputs_11_8_port, A(7) => 
                           MuxOutputs_11_7_port, A(6) => MuxOutputs_11_6_port, 
                           A(5) => MuxOutputs_11_5_port, A(4) => 
                           MuxOutputs_11_4_port, A(3) => MuxOutputs_11_3_port, 
                           A(2) => MuxOutputs_11_2_port, A(1) => 
                           MuxOutputs_11_1_port, A(0) => MuxOutputs_11_0_port, 
                           B(63) => SumOutputs_9_63_port, B(62) => 
                           SumOutputs_9_62_port, B(61) => SumOutputs_9_61_port,
                           B(60) => SumOutputs_9_60_port, B(59) => 
                           SumOutputs_9_59_port, B(58) => SumOutputs_9_58_port,
                           B(57) => SumOutputs_9_57_port, B(56) => 
                           SumOutputs_9_56_port, B(55) => SumOutputs_9_55_port,
                           B(54) => SumOutputs_9_54_port, B(53) => 
                           SumOutputs_9_53_port, B(52) => SumOutputs_9_52_port,
                           B(51) => SumOutputs_9_51_port, B(50) => 
                           SumOutputs_9_50_port, B(49) => SumOutputs_9_49_port,
                           B(48) => SumOutputs_9_48_port, B(47) => 
                           SumOutputs_9_47_port, B(46) => SumOutputs_9_46_port,
                           B(45) => SumOutputs_9_45_port, B(44) => 
                           SumOutputs_9_44_port, B(43) => SumOutputs_9_43_port,
                           B(42) => SumOutputs_9_42_port, B(41) => 
                           SumOutputs_9_41_port, B(40) => SumOutputs_9_40_port,
                           B(39) => SumOutputs_9_39_port, B(38) => 
                           SumOutputs_9_38_port, B(37) => SumOutputs_9_37_port,
                           B(36) => SumOutputs_9_36_port, B(35) => 
                           SumOutputs_9_35_port, B(34) => SumOutputs_9_34_port,
                           B(33) => SumOutputs_9_33_port, B(32) => 
                           SumOutputs_9_32_port, B(31) => SumOutputs_9_31_port,
                           B(30) => SumOutputs_9_30_port, B(29) => 
                           SumOutputs_9_29_port, B(28) => SumOutputs_9_28_port,
                           B(27) => SumOutputs_9_27_port, B(26) => 
                           SumOutputs_9_26_port, B(25) => SumOutputs_9_25_port,
                           B(24) => SumOutputs_9_24_port, B(23) => 
                           SumOutputs_9_23_port, B(22) => SumOutputs_9_22_port,
                           B(21) => SumOutputs_9_21_port, B(20) => 
                           SumOutputs_9_20_port, B(19) => SumOutputs_9_19_port,
                           B(18) => SumOutputs_9_18_port, B(17) => 
                           SumOutputs_9_17_port, B(16) => SumOutputs_9_16_port,
                           B(15) => SumOutputs_9_15_port, B(14) => 
                           SumOutputs_9_14_port, B(13) => SumOutputs_9_13_port,
                           B(12) => SumOutputs_9_12_port, B(11) => 
                           SumOutputs_9_11_port, B(10) => SumOutputs_9_10_port,
                           B(9) => SumOutputs_9_9_port, B(8) => 
                           SumOutputs_9_8_port, B(7) => SumOutputs_9_7_port, 
                           B(6) => SumOutputs_9_6_port, B(5) => 
                           SumOutputs_9_5_port, B(4) => SumOutputs_9_4_port, 
                           B(3) => SumOutputs_9_3_port, B(2) => 
                           SumOutputs_9_2_port, B(1) => SumOutputs_9_1_port, 
                           B(0) => SumOutputs_9_0_port, Ci => X_Logic0_port, 
                           S(63) => SumOutputs_10_63_port, S(62) => 
                           SumOutputs_10_62_port, S(61) => 
                           SumOutputs_10_61_port, S(60) => 
                           SumOutputs_10_60_port, S(59) => 
                           SumOutputs_10_59_port, S(58) => 
                           SumOutputs_10_58_port, S(57) => 
                           SumOutputs_10_57_port, S(56) => 
                           SumOutputs_10_56_port, S(55) => 
                           SumOutputs_10_55_port, S(54) => 
                           SumOutputs_10_54_port, S(53) => 
                           SumOutputs_10_53_port, S(52) => 
                           SumOutputs_10_52_port, S(51) => 
                           SumOutputs_10_51_port, S(50) => 
                           SumOutputs_10_50_port, S(49) => 
                           SumOutputs_10_49_port, S(48) => 
                           SumOutputs_10_48_port, S(47) => 
                           SumOutputs_10_47_port, S(46) => 
                           SumOutputs_10_46_port, S(45) => 
                           SumOutputs_10_45_port, S(44) => 
                           SumOutputs_10_44_port, S(43) => 
                           SumOutputs_10_43_port, S(42) => 
                           SumOutputs_10_42_port, S(41) => 
                           SumOutputs_10_41_port, S(40) => 
                           SumOutputs_10_40_port, S(39) => 
                           SumOutputs_10_39_port, S(38) => 
                           SumOutputs_10_38_port, S(37) => 
                           SumOutputs_10_37_port, S(36) => 
                           SumOutputs_10_36_port, S(35) => 
                           SumOutputs_10_35_port, S(34) => 
                           SumOutputs_10_34_port, S(33) => 
                           SumOutputs_10_33_port, S(32) => 
                           SumOutputs_10_32_port, S(31) => 
                           SumOutputs_10_31_port, S(30) => 
                           SumOutputs_10_30_port, S(29) => 
                           SumOutputs_10_29_port, S(28) => 
                           SumOutputs_10_28_port, S(27) => 
                           SumOutputs_10_27_port, S(26) => 
                           SumOutputs_10_26_port, S(25) => 
                           SumOutputs_10_25_port, S(24) => 
                           SumOutputs_10_24_port, S(23) => 
                           SumOutputs_10_23_port, S(22) => 
                           SumOutputs_10_22_port, S(21) => 
                           SumOutputs_10_21_port, S(20) => 
                           SumOutputs_10_20_port, S(19) => 
                           SumOutputs_10_19_port, S(18) => 
                           SumOutputs_10_18_port, S(17) => 
                           SumOutputs_10_17_port, S(16) => 
                           SumOutputs_10_16_port, S(15) => 
                           SumOutputs_10_15_port, S(14) => 
                           SumOutputs_10_14_port, S(13) => 
                           SumOutputs_10_13_port, S(12) => 
                           SumOutputs_10_12_port, S(11) => 
                           SumOutputs_10_11_port, S(10) => 
                           SumOutputs_10_10_port, S(9) => SumOutputs_10_9_port,
                           S(8) => SumOutputs_10_8_port, S(7) => 
                           SumOutputs_10_7_port, S(6) => SumOutputs_10_6_port, 
                           S(5) => SumOutputs_10_5_port, S(4) => 
                           SumOutputs_10_4_port, S(3) => SumOutputs_10_3_port, 
                           S(2) => SumOutputs_10_2_port, S(1) => 
                           SumOutputs_10_1_port, S(0) => SumOutputs_10_0_port, 
                           Co => n_1137);
   SUMI_11 : RCA_NbitRca64_4 port map( A(63) => MuxOutputs_12_63_port, A(62) =>
                           MuxOutputs_12_62_port, A(61) => 
                           MuxOutputs_12_61_port, A(60) => 
                           MuxOutputs_12_60_port, A(59) => 
                           MuxOutputs_12_59_port, A(58) => 
                           MuxOutputs_12_58_port, A(57) => 
                           MuxOutputs_12_57_port, A(56) => 
                           MuxOutputs_12_56_port, A(55) => 
                           MuxOutputs_12_55_port, A(54) => 
                           MuxOutputs_12_54_port, A(53) => 
                           MuxOutputs_12_53_port, A(52) => 
                           MuxOutputs_12_52_port, A(51) => 
                           MuxOutputs_12_51_port, A(50) => 
                           MuxOutputs_12_50_port, A(49) => 
                           MuxOutputs_12_49_port, A(48) => 
                           MuxOutputs_12_48_port, A(47) => 
                           MuxOutputs_12_47_port, A(46) => 
                           MuxOutputs_12_46_port, A(45) => 
                           MuxOutputs_12_45_port, A(44) => 
                           MuxOutputs_12_44_port, A(43) => 
                           MuxOutputs_12_43_port, A(42) => 
                           MuxOutputs_12_42_port, A(41) => 
                           MuxOutputs_12_41_port, A(40) => 
                           MuxOutputs_12_40_port, A(39) => 
                           MuxOutputs_12_39_port, A(38) => 
                           MuxOutputs_12_38_port, A(37) => 
                           MuxOutputs_12_37_port, A(36) => 
                           MuxOutputs_12_36_port, A(35) => 
                           MuxOutputs_12_35_port, A(34) => 
                           MuxOutputs_12_34_port, A(33) => 
                           MuxOutputs_12_33_port, A(32) => 
                           MuxOutputs_12_32_port, A(31) => 
                           MuxOutputs_12_31_port, A(30) => 
                           MuxOutputs_12_30_port, A(29) => 
                           MuxOutputs_12_29_port, A(28) => 
                           MuxOutputs_12_28_port, A(27) => 
                           MuxOutputs_12_27_port, A(26) => 
                           MuxOutputs_12_26_port, A(25) => 
                           MuxOutputs_12_25_port, A(24) => 
                           MuxOutputs_12_24_port, A(23) => 
                           MuxOutputs_12_23_port, A(22) => 
                           MuxOutputs_12_22_port, A(21) => 
                           MuxOutputs_12_21_port, A(20) => 
                           MuxOutputs_12_20_port, A(19) => 
                           MuxOutputs_12_19_port, A(18) => 
                           MuxOutputs_12_18_port, A(17) => 
                           MuxOutputs_12_17_port, A(16) => 
                           MuxOutputs_12_16_port, A(15) => 
                           MuxOutputs_12_15_port, A(14) => 
                           MuxOutputs_12_14_port, A(13) => 
                           MuxOutputs_12_13_port, A(12) => 
                           MuxOutputs_12_12_port, A(11) => 
                           MuxOutputs_12_11_port, A(10) => 
                           MuxOutputs_12_10_port, A(9) => MuxOutputs_12_9_port,
                           A(8) => MuxOutputs_12_8_port, A(7) => 
                           MuxOutputs_12_7_port, A(6) => MuxOutputs_12_6_port, 
                           A(5) => MuxOutputs_12_5_port, A(4) => 
                           MuxOutputs_12_4_port, A(3) => MuxOutputs_12_3_port, 
                           A(2) => MuxOutputs_12_2_port, A(1) => 
                           MuxOutputs_12_1_port, A(0) => MuxOutputs_12_0_port, 
                           B(63) => SumOutputs_10_63_port, B(62) => 
                           SumOutputs_10_62_port, B(61) => 
                           SumOutputs_10_61_port, B(60) => 
                           SumOutputs_10_60_port, B(59) => 
                           SumOutputs_10_59_port, B(58) => 
                           SumOutputs_10_58_port, B(57) => 
                           SumOutputs_10_57_port, B(56) => 
                           SumOutputs_10_56_port, B(55) => 
                           SumOutputs_10_55_port, B(54) => 
                           SumOutputs_10_54_port, B(53) => 
                           SumOutputs_10_53_port, B(52) => 
                           SumOutputs_10_52_port, B(51) => 
                           SumOutputs_10_51_port, B(50) => 
                           SumOutputs_10_50_port, B(49) => 
                           SumOutputs_10_49_port, B(48) => 
                           SumOutputs_10_48_port, B(47) => 
                           SumOutputs_10_47_port, B(46) => 
                           SumOutputs_10_46_port, B(45) => 
                           SumOutputs_10_45_port, B(44) => 
                           SumOutputs_10_44_port, B(43) => 
                           SumOutputs_10_43_port, B(42) => 
                           SumOutputs_10_42_port, B(41) => 
                           SumOutputs_10_41_port, B(40) => 
                           SumOutputs_10_40_port, B(39) => 
                           SumOutputs_10_39_port, B(38) => 
                           SumOutputs_10_38_port, B(37) => 
                           SumOutputs_10_37_port, B(36) => 
                           SumOutputs_10_36_port, B(35) => 
                           SumOutputs_10_35_port, B(34) => 
                           SumOutputs_10_34_port, B(33) => 
                           SumOutputs_10_33_port, B(32) => 
                           SumOutputs_10_32_port, B(31) => 
                           SumOutputs_10_31_port, B(30) => 
                           SumOutputs_10_30_port, B(29) => 
                           SumOutputs_10_29_port, B(28) => 
                           SumOutputs_10_28_port, B(27) => 
                           SumOutputs_10_27_port, B(26) => 
                           SumOutputs_10_26_port, B(25) => 
                           SumOutputs_10_25_port, B(24) => 
                           SumOutputs_10_24_port, B(23) => 
                           SumOutputs_10_23_port, B(22) => 
                           SumOutputs_10_22_port, B(21) => 
                           SumOutputs_10_21_port, B(20) => 
                           SumOutputs_10_20_port, B(19) => 
                           SumOutputs_10_19_port, B(18) => 
                           SumOutputs_10_18_port, B(17) => 
                           SumOutputs_10_17_port, B(16) => 
                           SumOutputs_10_16_port, B(15) => 
                           SumOutputs_10_15_port, B(14) => 
                           SumOutputs_10_14_port, B(13) => 
                           SumOutputs_10_13_port, B(12) => 
                           SumOutputs_10_12_port, B(11) => 
                           SumOutputs_10_11_port, B(10) => 
                           SumOutputs_10_10_port, B(9) => SumOutputs_10_9_port,
                           B(8) => SumOutputs_10_8_port, B(7) => 
                           SumOutputs_10_7_port, B(6) => SumOutputs_10_6_port, 
                           B(5) => SumOutputs_10_5_port, B(4) => 
                           SumOutputs_10_4_port, B(3) => SumOutputs_10_3_port, 
                           B(2) => SumOutputs_10_2_port, B(1) => 
                           SumOutputs_10_1_port, B(0) => SumOutputs_10_0_port, 
                           Ci => X_Logic0_port, S(63) => SumOutputs_11_63_port,
                           S(62) => SumOutputs_11_62_port, S(61) => 
                           SumOutputs_11_61_port, S(60) => 
                           SumOutputs_11_60_port, S(59) => 
                           SumOutputs_11_59_port, S(58) => 
                           SumOutputs_11_58_port, S(57) => 
                           SumOutputs_11_57_port, S(56) => 
                           SumOutputs_11_56_port, S(55) => 
                           SumOutputs_11_55_port, S(54) => 
                           SumOutputs_11_54_port, S(53) => 
                           SumOutputs_11_53_port, S(52) => 
                           SumOutputs_11_52_port, S(51) => 
                           SumOutputs_11_51_port, S(50) => 
                           SumOutputs_11_50_port, S(49) => 
                           SumOutputs_11_49_port, S(48) => 
                           SumOutputs_11_48_port, S(47) => 
                           SumOutputs_11_47_port, S(46) => 
                           SumOutputs_11_46_port, S(45) => 
                           SumOutputs_11_45_port, S(44) => 
                           SumOutputs_11_44_port, S(43) => 
                           SumOutputs_11_43_port, S(42) => 
                           SumOutputs_11_42_port, S(41) => 
                           SumOutputs_11_41_port, S(40) => 
                           SumOutputs_11_40_port, S(39) => 
                           SumOutputs_11_39_port, S(38) => 
                           SumOutputs_11_38_port, S(37) => 
                           SumOutputs_11_37_port, S(36) => 
                           SumOutputs_11_36_port, S(35) => 
                           SumOutputs_11_35_port, S(34) => 
                           SumOutputs_11_34_port, S(33) => 
                           SumOutputs_11_33_port, S(32) => 
                           SumOutputs_11_32_port, S(31) => 
                           SumOutputs_11_31_port, S(30) => 
                           SumOutputs_11_30_port, S(29) => 
                           SumOutputs_11_29_port, S(28) => 
                           SumOutputs_11_28_port, S(27) => 
                           SumOutputs_11_27_port, S(26) => 
                           SumOutputs_11_26_port, S(25) => 
                           SumOutputs_11_25_port, S(24) => 
                           SumOutputs_11_24_port, S(23) => 
                           SumOutputs_11_23_port, S(22) => 
                           SumOutputs_11_22_port, S(21) => 
                           SumOutputs_11_21_port, S(20) => 
                           SumOutputs_11_20_port, S(19) => 
                           SumOutputs_11_19_port, S(18) => 
                           SumOutputs_11_18_port, S(17) => 
                           SumOutputs_11_17_port, S(16) => 
                           SumOutputs_11_16_port, S(15) => 
                           SumOutputs_11_15_port, S(14) => 
                           SumOutputs_11_14_port, S(13) => 
                           SumOutputs_11_13_port, S(12) => 
                           SumOutputs_11_12_port, S(11) => 
                           SumOutputs_11_11_port, S(10) => 
                           SumOutputs_11_10_port, S(9) => SumOutputs_11_9_port,
                           S(8) => SumOutputs_11_8_port, S(7) => 
                           SumOutputs_11_7_port, S(6) => SumOutputs_11_6_port, 
                           S(5) => SumOutputs_11_5_port, S(4) => 
                           SumOutputs_11_4_port, S(3) => SumOutputs_11_3_port, 
                           S(2) => SumOutputs_11_2_port, S(1) => 
                           SumOutputs_11_1_port, S(0) => SumOutputs_11_0_port, 
                           Co => n_1138);
   SUMI_12 : RCA_NbitRca64_3 port map( A(63) => MuxOutputs_13_63_port, A(62) =>
                           MuxOutputs_13_62_port, A(61) => 
                           MuxOutputs_13_61_port, A(60) => 
                           MuxOutputs_13_60_port, A(59) => 
                           MuxOutputs_13_59_port, A(58) => 
                           MuxOutputs_13_58_port, A(57) => 
                           MuxOutputs_13_57_port, A(56) => 
                           MuxOutputs_13_56_port, A(55) => 
                           MuxOutputs_13_55_port, A(54) => 
                           MuxOutputs_13_54_port, A(53) => 
                           MuxOutputs_13_53_port, A(52) => 
                           MuxOutputs_13_52_port, A(51) => 
                           MuxOutputs_13_51_port, A(50) => 
                           MuxOutputs_13_50_port, A(49) => 
                           MuxOutputs_13_49_port, A(48) => 
                           MuxOutputs_13_48_port, A(47) => 
                           MuxOutputs_13_47_port, A(46) => 
                           MuxOutputs_13_46_port, A(45) => 
                           MuxOutputs_13_45_port, A(44) => 
                           MuxOutputs_13_44_port, A(43) => 
                           MuxOutputs_13_43_port, A(42) => 
                           MuxOutputs_13_42_port, A(41) => 
                           MuxOutputs_13_41_port, A(40) => 
                           MuxOutputs_13_40_port, A(39) => 
                           MuxOutputs_13_39_port, A(38) => 
                           MuxOutputs_13_38_port, A(37) => 
                           MuxOutputs_13_37_port, A(36) => 
                           MuxOutputs_13_36_port, A(35) => 
                           MuxOutputs_13_35_port, A(34) => 
                           MuxOutputs_13_34_port, A(33) => 
                           MuxOutputs_13_33_port, A(32) => 
                           MuxOutputs_13_32_port, A(31) => 
                           MuxOutputs_13_31_port, A(30) => 
                           MuxOutputs_13_30_port, A(29) => 
                           MuxOutputs_13_29_port, A(28) => 
                           MuxOutputs_13_28_port, A(27) => 
                           MuxOutputs_13_27_port, A(26) => 
                           MuxOutputs_13_26_port, A(25) => 
                           MuxOutputs_13_25_port, A(24) => 
                           MuxOutputs_13_24_port, A(23) => 
                           MuxOutputs_13_23_port, A(22) => 
                           MuxOutputs_13_22_port, A(21) => 
                           MuxOutputs_13_21_port, A(20) => 
                           MuxOutputs_13_20_port, A(19) => 
                           MuxOutputs_13_19_port, A(18) => 
                           MuxOutputs_13_18_port, A(17) => 
                           MuxOutputs_13_17_port, A(16) => 
                           MuxOutputs_13_16_port, A(15) => 
                           MuxOutputs_13_15_port, A(14) => 
                           MuxOutputs_13_14_port, A(13) => 
                           MuxOutputs_13_13_port, A(12) => 
                           MuxOutputs_13_12_port, A(11) => 
                           MuxOutputs_13_11_port, A(10) => 
                           MuxOutputs_13_10_port, A(9) => MuxOutputs_13_9_port,
                           A(8) => MuxOutputs_13_8_port, A(7) => 
                           MuxOutputs_13_7_port, A(6) => MuxOutputs_13_6_port, 
                           A(5) => MuxOutputs_13_5_port, A(4) => 
                           MuxOutputs_13_4_port, A(3) => MuxOutputs_13_3_port, 
                           A(2) => MuxOutputs_13_2_port, A(1) => 
                           MuxOutputs_13_1_port, A(0) => MuxOutputs_13_0_port, 
                           B(63) => SumOutputs_11_63_port, B(62) => 
                           SumOutputs_11_62_port, B(61) => 
                           SumOutputs_11_61_port, B(60) => 
                           SumOutputs_11_60_port, B(59) => 
                           SumOutputs_11_59_port, B(58) => 
                           SumOutputs_11_58_port, B(57) => 
                           SumOutputs_11_57_port, B(56) => 
                           SumOutputs_11_56_port, B(55) => 
                           SumOutputs_11_55_port, B(54) => 
                           SumOutputs_11_54_port, B(53) => 
                           SumOutputs_11_53_port, B(52) => 
                           SumOutputs_11_52_port, B(51) => 
                           SumOutputs_11_51_port, B(50) => 
                           SumOutputs_11_50_port, B(49) => 
                           SumOutputs_11_49_port, B(48) => 
                           SumOutputs_11_48_port, B(47) => 
                           SumOutputs_11_47_port, B(46) => 
                           SumOutputs_11_46_port, B(45) => 
                           SumOutputs_11_45_port, B(44) => 
                           SumOutputs_11_44_port, B(43) => 
                           SumOutputs_11_43_port, B(42) => 
                           SumOutputs_11_42_port, B(41) => 
                           SumOutputs_11_41_port, B(40) => 
                           SumOutputs_11_40_port, B(39) => 
                           SumOutputs_11_39_port, B(38) => 
                           SumOutputs_11_38_port, B(37) => 
                           SumOutputs_11_37_port, B(36) => 
                           SumOutputs_11_36_port, B(35) => 
                           SumOutputs_11_35_port, B(34) => 
                           SumOutputs_11_34_port, B(33) => 
                           SumOutputs_11_33_port, B(32) => 
                           SumOutputs_11_32_port, B(31) => 
                           SumOutputs_11_31_port, B(30) => 
                           SumOutputs_11_30_port, B(29) => 
                           SumOutputs_11_29_port, B(28) => 
                           SumOutputs_11_28_port, B(27) => 
                           SumOutputs_11_27_port, B(26) => 
                           SumOutputs_11_26_port, B(25) => 
                           SumOutputs_11_25_port, B(24) => 
                           SumOutputs_11_24_port, B(23) => 
                           SumOutputs_11_23_port, B(22) => 
                           SumOutputs_11_22_port, B(21) => 
                           SumOutputs_11_21_port, B(20) => 
                           SumOutputs_11_20_port, B(19) => 
                           SumOutputs_11_19_port, B(18) => 
                           SumOutputs_11_18_port, B(17) => 
                           SumOutputs_11_17_port, B(16) => 
                           SumOutputs_11_16_port, B(15) => 
                           SumOutputs_11_15_port, B(14) => 
                           SumOutputs_11_14_port, B(13) => 
                           SumOutputs_11_13_port, B(12) => 
                           SumOutputs_11_12_port, B(11) => 
                           SumOutputs_11_11_port, B(10) => 
                           SumOutputs_11_10_port, B(9) => SumOutputs_11_9_port,
                           B(8) => SumOutputs_11_8_port, B(7) => 
                           SumOutputs_11_7_port, B(6) => SumOutputs_11_6_port, 
                           B(5) => SumOutputs_11_5_port, B(4) => 
                           SumOutputs_11_4_port, B(3) => SumOutputs_11_3_port, 
                           B(2) => SumOutputs_11_2_port, B(1) => 
                           SumOutputs_11_1_port, B(0) => SumOutputs_11_0_port, 
                           Ci => X_Logic0_port, S(63) => SumOutputs_12_63_port,
                           S(62) => SumOutputs_12_62_port, S(61) => 
                           SumOutputs_12_61_port, S(60) => 
                           SumOutputs_12_60_port, S(59) => 
                           SumOutputs_12_59_port, S(58) => 
                           SumOutputs_12_58_port, S(57) => 
                           SumOutputs_12_57_port, S(56) => 
                           SumOutputs_12_56_port, S(55) => 
                           SumOutputs_12_55_port, S(54) => 
                           SumOutputs_12_54_port, S(53) => 
                           SumOutputs_12_53_port, S(52) => 
                           SumOutputs_12_52_port, S(51) => 
                           SumOutputs_12_51_port, S(50) => 
                           SumOutputs_12_50_port, S(49) => 
                           SumOutputs_12_49_port, S(48) => 
                           SumOutputs_12_48_port, S(47) => 
                           SumOutputs_12_47_port, S(46) => 
                           SumOutputs_12_46_port, S(45) => 
                           SumOutputs_12_45_port, S(44) => 
                           SumOutputs_12_44_port, S(43) => 
                           SumOutputs_12_43_port, S(42) => 
                           SumOutputs_12_42_port, S(41) => 
                           SumOutputs_12_41_port, S(40) => 
                           SumOutputs_12_40_port, S(39) => 
                           SumOutputs_12_39_port, S(38) => 
                           SumOutputs_12_38_port, S(37) => 
                           SumOutputs_12_37_port, S(36) => 
                           SumOutputs_12_36_port, S(35) => 
                           SumOutputs_12_35_port, S(34) => 
                           SumOutputs_12_34_port, S(33) => 
                           SumOutputs_12_33_port, S(32) => 
                           SumOutputs_12_32_port, S(31) => 
                           SumOutputs_12_31_port, S(30) => 
                           SumOutputs_12_30_port, S(29) => 
                           SumOutputs_12_29_port, S(28) => 
                           SumOutputs_12_28_port, S(27) => 
                           SumOutputs_12_27_port, S(26) => 
                           SumOutputs_12_26_port, S(25) => 
                           SumOutputs_12_25_port, S(24) => 
                           SumOutputs_12_24_port, S(23) => 
                           SumOutputs_12_23_port, S(22) => 
                           SumOutputs_12_22_port, S(21) => 
                           SumOutputs_12_21_port, S(20) => 
                           SumOutputs_12_20_port, S(19) => 
                           SumOutputs_12_19_port, S(18) => 
                           SumOutputs_12_18_port, S(17) => 
                           SumOutputs_12_17_port, S(16) => 
                           SumOutputs_12_16_port, S(15) => 
                           SumOutputs_12_15_port, S(14) => 
                           SumOutputs_12_14_port, S(13) => 
                           SumOutputs_12_13_port, S(12) => 
                           SumOutputs_12_12_port, S(11) => 
                           SumOutputs_12_11_port, S(10) => 
                           SumOutputs_12_10_port, S(9) => SumOutputs_12_9_port,
                           S(8) => SumOutputs_12_8_port, S(7) => 
                           SumOutputs_12_7_port, S(6) => SumOutputs_12_6_port, 
                           S(5) => SumOutputs_12_5_port, S(4) => 
                           SumOutputs_12_4_port, S(3) => SumOutputs_12_3_port, 
                           S(2) => SumOutputs_12_2_port, S(1) => 
                           SumOutputs_12_1_port, S(0) => SumOutputs_12_0_port, 
                           Co => n_1139);
   SUMI_13 : RCA_NbitRca64_2 port map( A(63) => MuxOutputs_14_63_port, A(62) =>
                           MuxOutputs_14_62_port, A(61) => 
                           MuxOutputs_14_61_port, A(60) => 
                           MuxOutputs_14_60_port, A(59) => 
                           MuxOutputs_14_59_port, A(58) => 
                           MuxOutputs_14_58_port, A(57) => 
                           MuxOutputs_14_57_port, A(56) => 
                           MuxOutputs_14_56_port, A(55) => 
                           MuxOutputs_14_55_port, A(54) => 
                           MuxOutputs_14_54_port, A(53) => 
                           MuxOutputs_14_53_port, A(52) => 
                           MuxOutputs_14_52_port, A(51) => 
                           MuxOutputs_14_51_port, A(50) => 
                           MuxOutputs_14_50_port, A(49) => 
                           MuxOutputs_14_49_port, A(48) => 
                           MuxOutputs_14_48_port, A(47) => 
                           MuxOutputs_14_47_port, A(46) => 
                           MuxOutputs_14_46_port, A(45) => 
                           MuxOutputs_14_45_port, A(44) => 
                           MuxOutputs_14_44_port, A(43) => 
                           MuxOutputs_14_43_port, A(42) => 
                           MuxOutputs_14_42_port, A(41) => 
                           MuxOutputs_14_41_port, A(40) => 
                           MuxOutputs_14_40_port, A(39) => 
                           MuxOutputs_14_39_port, A(38) => 
                           MuxOutputs_14_38_port, A(37) => 
                           MuxOutputs_14_37_port, A(36) => 
                           MuxOutputs_14_36_port, A(35) => 
                           MuxOutputs_14_35_port, A(34) => 
                           MuxOutputs_14_34_port, A(33) => 
                           MuxOutputs_14_33_port, A(32) => 
                           MuxOutputs_14_32_port, A(31) => 
                           MuxOutputs_14_31_port, A(30) => 
                           MuxOutputs_14_30_port, A(29) => 
                           MuxOutputs_14_29_port, A(28) => 
                           MuxOutputs_14_28_port, A(27) => 
                           MuxOutputs_14_27_port, A(26) => 
                           MuxOutputs_14_26_port, A(25) => 
                           MuxOutputs_14_25_port, A(24) => 
                           MuxOutputs_14_24_port, A(23) => 
                           MuxOutputs_14_23_port, A(22) => 
                           MuxOutputs_14_22_port, A(21) => 
                           MuxOutputs_14_21_port, A(20) => 
                           MuxOutputs_14_20_port, A(19) => 
                           MuxOutputs_14_19_port, A(18) => 
                           MuxOutputs_14_18_port, A(17) => 
                           MuxOutputs_14_17_port, A(16) => 
                           MuxOutputs_14_16_port, A(15) => 
                           MuxOutputs_14_15_port, A(14) => 
                           MuxOutputs_14_14_port, A(13) => 
                           MuxOutputs_14_13_port, A(12) => 
                           MuxOutputs_14_12_port, A(11) => 
                           MuxOutputs_14_11_port, A(10) => 
                           MuxOutputs_14_10_port, A(9) => MuxOutputs_14_9_port,
                           A(8) => MuxOutputs_14_8_port, A(7) => 
                           MuxOutputs_14_7_port, A(6) => MuxOutputs_14_6_port, 
                           A(5) => MuxOutputs_14_5_port, A(4) => 
                           MuxOutputs_14_4_port, A(3) => MuxOutputs_14_3_port, 
                           A(2) => MuxOutputs_14_2_port, A(1) => 
                           MuxOutputs_14_1_port, A(0) => MuxOutputs_14_0_port, 
                           B(63) => SumOutputs_12_63_port, B(62) => 
                           SumOutputs_12_62_port, B(61) => 
                           SumOutputs_12_61_port, B(60) => 
                           SumOutputs_12_60_port, B(59) => 
                           SumOutputs_12_59_port, B(58) => 
                           SumOutputs_12_58_port, B(57) => 
                           SumOutputs_12_57_port, B(56) => 
                           SumOutputs_12_56_port, B(55) => 
                           SumOutputs_12_55_port, B(54) => 
                           SumOutputs_12_54_port, B(53) => 
                           SumOutputs_12_53_port, B(52) => 
                           SumOutputs_12_52_port, B(51) => 
                           SumOutputs_12_51_port, B(50) => 
                           SumOutputs_12_50_port, B(49) => 
                           SumOutputs_12_49_port, B(48) => 
                           SumOutputs_12_48_port, B(47) => 
                           SumOutputs_12_47_port, B(46) => 
                           SumOutputs_12_46_port, B(45) => 
                           SumOutputs_12_45_port, B(44) => 
                           SumOutputs_12_44_port, B(43) => 
                           SumOutputs_12_43_port, B(42) => 
                           SumOutputs_12_42_port, B(41) => 
                           SumOutputs_12_41_port, B(40) => 
                           SumOutputs_12_40_port, B(39) => 
                           SumOutputs_12_39_port, B(38) => 
                           SumOutputs_12_38_port, B(37) => 
                           SumOutputs_12_37_port, B(36) => 
                           SumOutputs_12_36_port, B(35) => 
                           SumOutputs_12_35_port, B(34) => 
                           SumOutputs_12_34_port, B(33) => 
                           SumOutputs_12_33_port, B(32) => 
                           SumOutputs_12_32_port, B(31) => 
                           SumOutputs_12_31_port, B(30) => 
                           SumOutputs_12_30_port, B(29) => 
                           SumOutputs_12_29_port, B(28) => 
                           SumOutputs_12_28_port, B(27) => 
                           SumOutputs_12_27_port, B(26) => 
                           SumOutputs_12_26_port, B(25) => 
                           SumOutputs_12_25_port, B(24) => 
                           SumOutputs_12_24_port, B(23) => 
                           SumOutputs_12_23_port, B(22) => 
                           SumOutputs_12_22_port, B(21) => 
                           SumOutputs_12_21_port, B(20) => 
                           SumOutputs_12_20_port, B(19) => 
                           SumOutputs_12_19_port, B(18) => 
                           SumOutputs_12_18_port, B(17) => 
                           SumOutputs_12_17_port, B(16) => 
                           SumOutputs_12_16_port, B(15) => 
                           SumOutputs_12_15_port, B(14) => 
                           SumOutputs_12_14_port, B(13) => 
                           SumOutputs_12_13_port, B(12) => 
                           SumOutputs_12_12_port, B(11) => 
                           SumOutputs_12_11_port, B(10) => 
                           SumOutputs_12_10_port, B(9) => SumOutputs_12_9_port,
                           B(8) => SumOutputs_12_8_port, B(7) => 
                           SumOutputs_12_7_port, B(6) => SumOutputs_12_6_port, 
                           B(5) => SumOutputs_12_5_port, B(4) => 
                           SumOutputs_12_4_port, B(3) => SumOutputs_12_3_port, 
                           B(2) => SumOutputs_12_2_port, B(1) => 
                           SumOutputs_12_1_port, B(0) => SumOutputs_12_0_port, 
                           Ci => X_Logic0_port, S(63) => SumOutputs_13_63_port,
                           S(62) => SumOutputs_13_62_port, S(61) => 
                           SumOutputs_13_61_port, S(60) => 
                           SumOutputs_13_60_port, S(59) => 
                           SumOutputs_13_59_port, S(58) => 
                           SumOutputs_13_58_port, S(57) => 
                           SumOutputs_13_57_port, S(56) => 
                           SumOutputs_13_56_port, S(55) => 
                           SumOutputs_13_55_port, S(54) => 
                           SumOutputs_13_54_port, S(53) => 
                           SumOutputs_13_53_port, S(52) => 
                           SumOutputs_13_52_port, S(51) => 
                           SumOutputs_13_51_port, S(50) => 
                           SumOutputs_13_50_port, S(49) => 
                           SumOutputs_13_49_port, S(48) => 
                           SumOutputs_13_48_port, S(47) => 
                           SumOutputs_13_47_port, S(46) => 
                           SumOutputs_13_46_port, S(45) => 
                           SumOutputs_13_45_port, S(44) => 
                           SumOutputs_13_44_port, S(43) => 
                           SumOutputs_13_43_port, S(42) => 
                           SumOutputs_13_42_port, S(41) => 
                           SumOutputs_13_41_port, S(40) => 
                           SumOutputs_13_40_port, S(39) => 
                           SumOutputs_13_39_port, S(38) => 
                           SumOutputs_13_38_port, S(37) => 
                           SumOutputs_13_37_port, S(36) => 
                           SumOutputs_13_36_port, S(35) => 
                           SumOutputs_13_35_port, S(34) => 
                           SumOutputs_13_34_port, S(33) => 
                           SumOutputs_13_33_port, S(32) => 
                           SumOutputs_13_32_port, S(31) => 
                           SumOutputs_13_31_port, S(30) => 
                           SumOutputs_13_30_port, S(29) => 
                           SumOutputs_13_29_port, S(28) => 
                           SumOutputs_13_28_port, S(27) => 
                           SumOutputs_13_27_port, S(26) => 
                           SumOutputs_13_26_port, S(25) => 
                           SumOutputs_13_25_port, S(24) => 
                           SumOutputs_13_24_port, S(23) => 
                           SumOutputs_13_23_port, S(22) => 
                           SumOutputs_13_22_port, S(21) => 
                           SumOutputs_13_21_port, S(20) => 
                           SumOutputs_13_20_port, S(19) => 
                           SumOutputs_13_19_port, S(18) => 
                           SumOutputs_13_18_port, S(17) => 
                           SumOutputs_13_17_port, S(16) => 
                           SumOutputs_13_16_port, S(15) => 
                           SumOutputs_13_15_port, S(14) => 
                           SumOutputs_13_14_port, S(13) => 
                           SumOutputs_13_13_port, S(12) => 
                           SumOutputs_13_12_port, S(11) => 
                           SumOutputs_13_11_port, S(10) => 
                           SumOutputs_13_10_port, S(9) => SumOutputs_13_9_port,
                           S(8) => SumOutputs_13_8_port, S(7) => 
                           SumOutputs_13_7_port, S(6) => SumOutputs_13_6_port, 
                           S(5) => SumOutputs_13_5_port, S(4) => 
                           SumOutputs_13_4_port, S(3) => SumOutputs_13_3_port, 
                           S(2) => SumOutputs_13_2_port, S(1) => 
                           SumOutputs_13_1_port, S(0) => SumOutputs_13_0_port, 
                           Co => n_1140);
   SUMI_14 : RCA_NbitRca64_1 port map( A(63) => MuxOutputs_15_63_port, A(62) =>
                           MuxOutputs_15_62_port, A(61) => 
                           MuxOutputs_15_61_port, A(60) => 
                           MuxOutputs_15_60_port, A(59) => 
                           MuxOutputs_15_59_port, A(58) => 
                           MuxOutputs_15_58_port, A(57) => 
                           MuxOutputs_15_57_port, A(56) => 
                           MuxOutputs_15_56_port, A(55) => 
                           MuxOutputs_15_55_port, A(54) => 
                           MuxOutputs_15_54_port, A(53) => 
                           MuxOutputs_15_53_port, A(52) => 
                           MuxOutputs_15_52_port, A(51) => 
                           MuxOutputs_15_51_port, A(50) => 
                           MuxOutputs_15_50_port, A(49) => 
                           MuxOutputs_15_49_port, A(48) => 
                           MuxOutputs_15_48_port, A(47) => 
                           MuxOutputs_15_47_port, A(46) => 
                           MuxOutputs_15_46_port, A(45) => 
                           MuxOutputs_15_45_port, A(44) => 
                           MuxOutputs_15_44_port, A(43) => 
                           MuxOutputs_15_43_port, A(42) => 
                           MuxOutputs_15_42_port, A(41) => 
                           MuxOutputs_15_41_port, A(40) => 
                           MuxOutputs_15_40_port, A(39) => 
                           MuxOutputs_15_39_port, A(38) => 
                           MuxOutputs_15_38_port, A(37) => 
                           MuxOutputs_15_37_port, A(36) => 
                           MuxOutputs_15_36_port, A(35) => 
                           MuxOutputs_15_35_port, A(34) => 
                           MuxOutputs_15_34_port, A(33) => 
                           MuxOutputs_15_33_port, A(32) => 
                           MuxOutputs_15_32_port, A(31) => 
                           MuxOutputs_15_31_port, A(30) => 
                           MuxOutputs_15_30_port, A(29) => 
                           MuxOutputs_15_29_port, A(28) => 
                           MuxOutputs_15_28_port, A(27) => 
                           MuxOutputs_15_27_port, A(26) => 
                           MuxOutputs_15_26_port, A(25) => 
                           MuxOutputs_15_25_port, A(24) => 
                           MuxOutputs_15_24_port, A(23) => 
                           MuxOutputs_15_23_port, A(22) => 
                           MuxOutputs_15_22_port, A(21) => 
                           MuxOutputs_15_21_port, A(20) => 
                           MuxOutputs_15_20_port, A(19) => 
                           MuxOutputs_15_19_port, A(18) => 
                           MuxOutputs_15_18_port, A(17) => 
                           MuxOutputs_15_17_port, A(16) => 
                           MuxOutputs_15_16_port, A(15) => 
                           MuxOutputs_15_15_port, A(14) => 
                           MuxOutputs_15_14_port, A(13) => 
                           MuxOutputs_15_13_port, A(12) => 
                           MuxOutputs_15_12_port, A(11) => 
                           MuxOutputs_15_11_port, A(10) => 
                           MuxOutputs_15_10_port, A(9) => MuxOutputs_15_9_port,
                           A(8) => MuxOutputs_15_8_port, A(7) => 
                           MuxOutputs_15_7_port, A(6) => MuxOutputs_15_6_port, 
                           A(5) => MuxOutputs_15_5_port, A(4) => 
                           MuxOutputs_15_4_port, A(3) => MuxOutputs_15_3_port, 
                           A(2) => MuxOutputs_15_2_port, A(1) => 
                           MuxOutputs_15_1_port, A(0) => MuxOutputs_15_0_port, 
                           B(63) => SumOutputs_13_63_port, B(62) => 
                           SumOutputs_13_62_port, B(61) => 
                           SumOutputs_13_61_port, B(60) => 
                           SumOutputs_13_60_port, B(59) => 
                           SumOutputs_13_59_port, B(58) => 
                           SumOutputs_13_58_port, B(57) => 
                           SumOutputs_13_57_port, B(56) => 
                           SumOutputs_13_56_port, B(55) => 
                           SumOutputs_13_55_port, B(54) => 
                           SumOutputs_13_54_port, B(53) => 
                           SumOutputs_13_53_port, B(52) => 
                           SumOutputs_13_52_port, B(51) => 
                           SumOutputs_13_51_port, B(50) => 
                           SumOutputs_13_50_port, B(49) => 
                           SumOutputs_13_49_port, B(48) => 
                           SumOutputs_13_48_port, B(47) => 
                           SumOutputs_13_47_port, B(46) => 
                           SumOutputs_13_46_port, B(45) => 
                           SumOutputs_13_45_port, B(44) => 
                           SumOutputs_13_44_port, B(43) => 
                           SumOutputs_13_43_port, B(42) => 
                           SumOutputs_13_42_port, B(41) => 
                           SumOutputs_13_41_port, B(40) => 
                           SumOutputs_13_40_port, B(39) => 
                           SumOutputs_13_39_port, B(38) => 
                           SumOutputs_13_38_port, B(37) => 
                           SumOutputs_13_37_port, B(36) => 
                           SumOutputs_13_36_port, B(35) => 
                           SumOutputs_13_35_port, B(34) => 
                           SumOutputs_13_34_port, B(33) => 
                           SumOutputs_13_33_port, B(32) => 
                           SumOutputs_13_32_port, B(31) => 
                           SumOutputs_13_31_port, B(30) => 
                           SumOutputs_13_30_port, B(29) => 
                           SumOutputs_13_29_port, B(28) => 
                           SumOutputs_13_28_port, B(27) => 
                           SumOutputs_13_27_port, B(26) => 
                           SumOutputs_13_26_port, B(25) => 
                           SumOutputs_13_25_port, B(24) => 
                           SumOutputs_13_24_port, B(23) => 
                           SumOutputs_13_23_port, B(22) => 
                           SumOutputs_13_22_port, B(21) => 
                           SumOutputs_13_21_port, B(20) => 
                           SumOutputs_13_20_port, B(19) => 
                           SumOutputs_13_19_port, B(18) => 
                           SumOutputs_13_18_port, B(17) => 
                           SumOutputs_13_17_port, B(16) => 
                           SumOutputs_13_16_port, B(15) => 
                           SumOutputs_13_15_port, B(14) => 
                           SumOutputs_13_14_port, B(13) => 
                           SumOutputs_13_13_port, B(12) => 
                           SumOutputs_13_12_port, B(11) => 
                           SumOutputs_13_11_port, B(10) => 
                           SumOutputs_13_10_port, B(9) => SumOutputs_13_9_port,
                           B(8) => SumOutputs_13_8_port, B(7) => 
                           SumOutputs_13_7_port, B(6) => SumOutputs_13_6_port, 
                           B(5) => SumOutputs_13_5_port, B(4) => 
                           SumOutputs_13_4_port, B(3) => SumOutputs_13_3_port, 
                           B(2) => SumOutputs_13_2_port, B(1) => 
                           SumOutputs_13_1_port, B(0) => SumOutputs_13_0_port, 
                           Ci => X_Logic0_port, S(63) => P(63), S(62) => P(62),
                           S(61) => P(61), S(60) => P(60), S(59) => P(59), 
                           S(58) => P(58), S(57) => P(57), S(56) => P(56), 
                           S(55) => P(55), S(54) => P(54), S(53) => P(53), 
                           S(52) => P(52), S(51) => P(51), S(50) => P(50), 
                           S(49) => P(49), S(48) => P(48), S(47) => P(47), 
                           S(46) => P(46), S(45) => P(45), S(44) => P(44), 
                           S(43) => P(43), S(42) => P(42), S(41) => P(41), 
                           S(40) => P(40), S(39) => P(39), S(38) => P(38), 
                           S(37) => P(37), S(36) => P(36), S(35) => P(35), 
                           S(34) => P(34), S(33) => P(33), S(32) => P(32), 
                           S(31) => P(31), S(30) => P(30), S(29) => P(29), 
                           S(28) => P(28), S(27) => P(27), S(26) => P(26), 
                           S(25) => P(25), S(24) => P(24), S(23) => P(23), 
                           S(22) => P(22), S(21) => P(21), S(20) => P(20), 
                           S(19) => P(19), S(18) => P(18), S(17) => P(17), 
                           S(16) => P(16), S(15) => P(15), S(14) => P(14), 
                           S(13) => P(13), S(12) => P(12), S(11) => P(11), 
                           S(10) => P(10), S(9) => P(9), S(8) => P(8), S(7) => 
                           P(7), S(6) => P(6), S(5) => P(5), S(4) => P(4), S(3)
                           => P(3), S(2) => P(2), S(1) => P(1), S(0) => P(0), 
                           Co => n_1141);
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   n9 <= '0';
   U3 : BUF_X1 port map( A => negative_inputs_1_11_port, Z => n17);
   U4 : CLKBUF_X1 port map( A => negative_inputs_1_13_port, Z => n13);
   U5 : BUF_X1 port map( A => negative_inputs_0_15_port, Z => n40);
   U6 : BUF_X1 port map( A => negative_inputs_0_20_port, Z => n32);
   U7 : BUF_X1 port map( A => negative_inputs_0_24_port, Z => n10);
   U8 : BUF_X1 port map( A => negative_inputs_0_27_port, Z => n25);
   U9 : BUF_X1 port map( A => negative_inputs_0_28_port, Z => n28);
   U10 : BUF_X1 port map( A => negative_inputs_0_30_port, Z => n22);
   U12 : BUF_X1 port map( A => negative_inputs_0_29_port, Z => n24);
   U13 : BUF_X1 port map( A => negative_inputs_0_31_port, Z => n23);
   U14 : BUF_X1 port map( A => negative_inputs_0_32_port, Z => n15);
   U15 : BUF_X1 port map( A => negative_inputs_0_39_port, Z => n151);
   U16 : BUF_X1 port map( A => negative_inputs_0_47_port, Z => n14);
   U17 : CLKBUF_X1 port map( A => negative_inputs_1_10_port, Z => n18);
   U18 : BUF_X1 port map( A => A(1), Z => n11);
   U19 : BUF_X1 port map( A => negative_inputs_1_3_port, Z => n12);
   U20 : BUF_X2 port map( A => negative_inputs_0_11_port, Z => n43);
   U21 : CLKBUF_X1 port map( A => negative_inputs_1_8_port, Z => n20);
   U22 : BUF_X2 port map( A => negative_inputs_0_17_port, Z => n16);
   U23 : CLKBUF_X1 port map( A => negative_inputs_7_28_port, Z => n115);
   U24 : INV_X2 port map( A => n30, ZN => n31);
   U25 : BUF_X1 port map( A => negative_inputs_0_10_port, Z => n46);
   U26 : CLKBUF_X1 port map( A => negative_inputs_7_25_port, Z => n109);
   U27 : BUF_X1 port map( A => negative_inputs_0_9_port, Z => n45);
   U28 : BUF_X2 port map( A => negative_inputs_0_16_port, Z => n19);
   U29 : BUF_X1 port map( A => negative_inputs_1_5_port, Z => n21);
   U30 : CLKBUF_X1 port map( A => negative_inputs_0_4_port, Z => n37);
   U31 : BUF_X1 port map( A => A(0), Z => n72);
   U32 : INV_X1 port map( A => negative_inputs_0_46_port, ZN => n26);
   U33 : INV_X1 port map( A => n26, ZN => n27);
   U34 : BUF_X2 port map( A => negative_inputs_0_19_port, Z => n29);
   U35 : INV_X1 port map( A => negative_inputs_0_45_port, ZN => n30);
   U36 : BUF_X1 port map( A => negative_inputs_7_10_port, Z => n79);
   U37 : BUF_X2 port map( A => negative_inputs_0_22_port, Z => n33);
   U38 : BUF_X1 port map( A => negative_inputs_1_6_port, Z => n34);
   U39 : BUF_X1 port map( A => negative_inputs_0_5_port, Z => n48);
   U40 : BUF_X1 port map( A => negative_inputs_1_7_port, Z => n35);
   U41 : BUF_X2 port map( A => negative_inputs_0_25_port, Z => n36);
   U42 : BUF_X2 port map( A => negative_inputs_0_3_port, Z => n71);
   U43 : CLKBUF_X1 port map( A => negative_inputs_7_11_port, Z => n81);
   U44 : BUF_X2 port map( A => negative_inputs_0_13_port, Z => n38);
   U45 : BUF_X2 port map( A => negative_inputs_0_23_port, Z => n39);
   U46 : CLKBUF_X1 port map( A => negative_inputs_7_22_port, Z => n103);
   U47 : CLKBUF_X1 port map( A => negative_inputs_7_31_port, Z => n121);
   U48 : INV_X1 port map( A => negative_inputs_1_43_port, ZN => n41);
   U49 : INV_X1 port map( A => n41, ZN => n42);
   U50 : CLKBUF_X1 port map( A => negative_inputs_7_32_port, Z => n123);
   U51 : BUF_X2 port map( A => negative_inputs_0_8_port, Z => n44);
   U52 : CLKBUF_X1 port map( A => negative_inputs_7_30_port, Z => n119);
   U53 : CLKBUF_X1 port map( A => negative_inputs_7_24_port, Z => n107);
   U54 : BUF_X2 port map( A => negative_inputs_0_14_port, Z => n47);
   U55 : CLKBUF_X1 port map( A => negative_inputs_7_13_port, Z => n85);
   U56 : CLKBUF_X1 port map( A => negative_inputs_7_15_port, Z => n89);
   U57 : CLKBUF_X1 port map( A => negative_inputs_7_18_port, Z => n95);
   U58 : CLKBUF_X1 port map( A => negative_inputs_7_16_port, Z => n91);
   U59 : CLKBUF_X1 port map( A => negative_inputs_7_14_port, Z => n87);
   U60 : CLKBUF_X1 port map( A => negative_inputs_7_12_port, Z => n83);
   U61 : CLKBUF_X1 port map( A => negative_inputs_11_48_port, Z => n148);
   U62 : CLKBUF_X1 port map( A => negative_inputs_12_48_port, Z => n146);
   U63 : CLKBUF_X1 port map( A => negative_inputs_13_48_port, Z => n144);
   U64 : CLKBUF_X1 port map( A => negative_inputs_14_48_port, Z => n142);
   U65 : CLKBUF_X1 port map( A => negative_inputs_10_48_port, Z => n150);
   U66 : CLKBUF_X1 port map( A => positive_inputs_7_7_port, Z => n154);
   U67 : BUF_X1 port map( A => positive_inputs_7_20_port, Z => n180);
   U68 : BUF_X1 port map( A => positive_inputs_7_21_port, Z => n182);
   U69 : BUF_X1 port map( A => positive_inputs_7_22_port, Z => n184);
   U70 : BUF_X1 port map( A => positive_inputs_7_23_port, Z => n186);
   U71 : BUF_X1 port map( A => positive_inputs_7_24_port, Z => n188);
   U72 : BUF_X1 port map( A => positive_inputs_7_25_port, Z => n190);
   U73 : BUF_X1 port map( A => positive_inputs_7_26_port, Z => n192);
   U74 : BUF_X1 port map( A => positive_inputs_7_27_port, Z => n194);
   U75 : BUF_X1 port map( A => positive_inputs_7_28_port, Z => n196);
   U76 : BUF_X1 port map( A => positive_inputs_7_29_port, Z => n198);
   U77 : BUF_X1 port map( A => positive_inputs_7_30_port, Z => n200);
   U78 : BUF_X1 port map( A => positive_inputs_7_31_port, Z => n202);
   U79 : BUF_X1 port map( A => positive_inputs_7_32_port, Z => n204);
   U80 : BUF_X1 port map( A => positive_inputs_7_33_port, Z => n206);
   U81 : BUF_X1 port map( A => positive_inputs_7_34_port, Z => n208);
   U82 : BUF_X1 port map( A => positive_inputs_2_38_port, Z => n49);
   U83 : BUF_X1 port map( A => positive_inputs_1_38_port, Z => n50);
   U84 : BUF_X1 port map( A => positive_inputs_7_35_port, Z => n210);
   U85 : BUF_X1 port map( A => positive_inputs_7_36_port, Z => n212);
   U86 : BUF_X1 port map( A => positive_inputs_7_37_port, Z => n214);
   U87 : BUF_X1 port map( A => positive_inputs_4_39_port, Z => n55);
   U88 : BUF_X1 port map( A => positive_inputs_5_39_port, Z => n54);
   U89 : BUF_X1 port map( A => positive_inputs_7_38_port, Z => n51);
   U90 : BUF_X1 port map( A => positive_inputs_7_39_port, Z => n52);
   U91 : BUF_X1 port map( A => positive_inputs_6_39_port, Z => n53);
   U92 : BUF_X1 port map( A => positive_inputs_2_48_port, Z => n69);
   U93 : BUF_X1 port map( A => positive_inputs_1_48_port, Z => n70);
   U94 : BUF_X1 port map( A => positive_inputs_4_48_port, Z => n68);
   U95 : BUF_X1 port map( A => positive_inputs_5_48_port, Z => n67);
   U96 : BUF_X1 port map( A => positive_inputs_7_48_port, Z => n66);
   U97 : BUF_X1 port map( A => positive_inputs_8_48_port, Z => n65);
   U98 : BUF_X1 port map( A => positive_inputs_9_48_port, Z => n64);
   U99 : BUF_X1 port map( A => positive_inputs_10_48_port, Z => n63);
   U100 : BUF_X1 port map( A => negative_inputs_16_19_port, Z => n80);
   U101 : BUF_X1 port map( A => negative_inputs_16_42_port, Z => n126);
   U102 : BUF_X1 port map( A => negative_inputs_16_41_port, Z => n124);
   U103 : BUF_X1 port map( A => negative_inputs_15_48_port, Z => n140);
   U104 : BUF_X1 port map( A => negative_inputs_16_17_port, Z => n76);
   U105 : BUF_X1 port map( A => negative_inputs_16_31_port, Z => n104);
   U106 : BUF_X1 port map( A => negative_inputs_16_29_port, Z => n100);
   U107 : BUF_X1 port map( A => negative_inputs_16_30_port, Z => n102);
   U108 : BUF_X1 port map( A => negative_inputs_16_32_port, Z => n106);
   U109 : BUF_X1 port map( A => negative_inputs_16_33_port, Z => n108);
   U110 : BUF_X1 port map( A => negative_inputs_16_35_port, Z => n112);
   U111 : BUF_X1 port map( A => negative_inputs_16_36_port, Z => n114);
   U112 : BUF_X1 port map( A => negative_inputs_16_37_port, Z => n116);
   U113 : BUF_X1 port map( A => negative_inputs_16_38_port, Z => n118);
   U114 : BUF_X1 port map( A => negative_inputs_16_39_port, Z => n120);
   U115 : BUF_X1 port map( A => negative_inputs_16_40_port, Z => n122);
   U116 : BUF_X1 port map( A => negative_inputs_16_43_port, Z => n128);
   U117 : BUF_X1 port map( A => negative_inputs_16_44_port, Z => n130);
   U118 : BUF_X1 port map( A => negative_inputs_16_46_port, Z => n134);
   U119 : BUF_X1 port map( A => negative_inputs_16_47_port, Z => n136);
   U120 : BUF_X1 port map( A => negative_inputs_16_48_port, Z => n138);
   U121 : BUF_X1 port map( A => negative_inputs_16_18_port, Z => n78);
   U122 : BUF_X1 port map( A => negative_inputs_16_26_port, Z => n94);
   U123 : BUF_X1 port map( A => negative_inputs_16_28_port, Z => n98);
   U124 : BUF_X1 port map( A => negative_inputs_16_20_port, Z => n82);
   U125 : BUF_X1 port map( A => negative_inputs_16_25_port, Z => n92);
   U126 : BUF_X1 port map( A => negative_inputs_16_23_port, Z => n88);
   U127 : BUF_X1 port map( A => negative_inputs_16_24_port, Z => n90);
   U128 : BUF_X1 port map( A => negative_inputs_16_27_port, Z => n96);
   U129 : BUF_X1 port map( A => negative_inputs_16_34_port, Z => n110);
   U130 : BUF_X1 port map( A => negative_inputs_16_45_port, Z => n132);
   U131 : BUF_X1 port map( A => negative_inputs_16_21_port, Z => n84);
   U132 : BUF_X1 port map( A => negative_inputs_16_22_port, Z => n86);
   U133 : BUF_X1 port map( A => negative_inputs_2_39_port, Z => n147);
   U134 : BUF_X1 port map( A => negative_inputs_3_39_port, Z => n145);
   U135 : BUF_X1 port map( A => negative_inputs_1_39_port, Z => n149);
   U136 : BUF_X1 port map( A => negative_inputs_4_39_port, Z => n143);
   U137 : BUF_X1 port map( A => negative_inputs_5_39_port, Z => n141);
   U138 : BUF_X1 port map( A => negative_inputs_7_8_port, Z => n75);
   U139 : BUF_X1 port map( A => negative_inputs_7_20_port, Z => n99);
   U140 : BUF_X1 port map( A => negative_inputs_7_21_port, Z => n101);
   U141 : BUF_X1 port map( A => negative_inputs_7_23_port, Z => n105);
   U142 : BUF_X1 port map( A => negative_inputs_7_26_port, Z => n111);
   U143 : BUF_X1 port map( A => negative_inputs_7_27_port, Z => n113);
   U144 : BUF_X1 port map( A => negative_inputs_7_29_port, Z => n117);
   U145 : BUF_X1 port map( A => negative_inputs_7_34_port, Z => n127);
   U146 : BUF_X1 port map( A => negative_inputs_7_33_port, Z => n125);
   U147 : BUF_X1 port map( A => negative_inputs_6_39_port, Z => n139);
   U148 : BUF_X1 port map( A => negative_inputs_7_35_port, Z => n129);
   U149 : BUF_X1 port map( A => negative_inputs_7_37_port, Z => n133);
   U150 : BUF_X1 port map( A => negative_inputs_7_38_port, Z => n135);
   U151 : BUF_X1 port map( A => negative_inputs_7_39_port, Z => n137);
   U152 : BUF_X1 port map( A => negative_inputs_7_36_port, Z => n131);
   U153 : BUF_X1 port map( A => negative_inputs_8_48_port, Z => n153);
   U154 : BUF_X1 port map( A => negative_inputs_9_48_port, Z => n152);
   U155 : BUF_X1 port map( A => negative_inputs_16_16_port, Z => n74);
   U156 : BUF_X1 port map( A => positive_inputs_16_16_port, Z => n155);
   U157 : BUF_X1 port map( A => negative_inputs_7_7_port, Z => n73);
   U158 : BUF_X1 port map( A => positive_inputs_16_17_port, Z => n157);
   U159 : BUF_X1 port map( A => positive_inputs_16_18_port, Z => n159);
   U160 : BUF_X1 port map( A => positive_inputs_16_19_port, Z => n161);
   U161 : BUF_X1 port map( A => positive_inputs_16_20_port, Z => n163);
   U162 : BUF_X1 port map( A => positive_inputs_16_21_port, Z => n165);
   U163 : BUF_X1 port map( A => positive_inputs_16_22_port, Z => n167);
   U164 : BUF_X1 port map( A => positive_inputs_16_23_port, Z => n169);
   U165 : BUF_X1 port map( A => positive_inputs_16_24_port, Z => n171);
   U166 : BUF_X1 port map( A => positive_inputs_16_25_port, Z => n173);
   U167 : BUF_X1 port map( A => positive_inputs_16_26_port, Z => n175);
   U168 : BUF_X1 port map( A => positive_inputs_16_27_port, Z => n177);
   U169 : BUF_X1 port map( A => positive_inputs_16_28_port, Z => n179);
   U170 : BUF_X1 port map( A => positive_inputs_16_29_port, Z => n181);
   U171 : BUF_X1 port map( A => positive_inputs_16_30_port, Z => n183);
   U172 : BUF_X1 port map( A => positive_inputs_16_31_port, Z => n185);
   U173 : BUF_X1 port map( A => positive_inputs_16_32_port, Z => n187);
   U174 : BUF_X1 port map( A => positive_inputs_16_33_port, Z => n189);
   U175 : BUF_X1 port map( A => positive_inputs_16_34_port, Z => n191);
   U176 : BUF_X1 port map( A => positive_inputs_16_35_port, Z => n193);
   U177 : BUF_X1 port map( A => positive_inputs_16_36_port, Z => n195);
   U178 : BUF_X1 port map( A => positive_inputs_16_37_port, Z => n197);
   U179 : BUF_X1 port map( A => positive_inputs_16_41_port, Z => n205);
   U180 : BUF_X1 port map( A => positive_inputs_16_42_port, Z => n207);
   U181 : BUF_X1 port map( A => positive_inputs_16_38_port, Z => n199);
   U182 : BUF_X1 port map( A => positive_inputs_16_39_port, Z => n201);
   U183 : BUF_X1 port map( A => positive_inputs_16_40_port, Z => n203);
   U184 : BUF_X1 port map( A => positive_inputs_11_48_port, Z => n62);
   U185 : BUF_X1 port map( A => positive_inputs_16_43_port, Z => n209);
   U186 : BUF_X1 port map( A => positive_inputs_13_48_port, Z => n60);
   U187 : BUF_X1 port map( A => positive_inputs_12_48_port, Z => n61);
   U188 : BUF_X1 port map( A => positive_inputs_16_44_port, Z => n211);
   U189 : BUF_X1 port map( A => positive_inputs_16_45_port, Z => n213);
   U190 : BUF_X1 port map( A => positive_inputs_15_48_port, Z => n58);
   U191 : BUF_X1 port map( A => positive_inputs_14_48_port, Z => n59);
   U192 : BUF_X1 port map( A => positive_inputs_16_46_port, Z => n215);
   U193 : BUF_X1 port map( A => positive_inputs_16_47_port, Z => n56);
   U194 : BUF_X1 port map( A => positive_inputs_16_48_port, Z => n57);
   U195 : BUF_X1 port map( A => positive_inputs_7_8_port, Z => n156);
   U196 : BUF_X1 port map( A => positive_inputs_7_9_port, Z => n158);
   U197 : BUF_X1 port map( A => positive_inputs_7_10_port, Z => n160);
   U198 : BUF_X1 port map( A => positive_inputs_7_11_port, Z => n162);
   U199 : BUF_X1 port map( A => positive_inputs_7_12_port, Z => n164);
   U200 : BUF_X1 port map( A => positive_inputs_7_13_port, Z => n166);
   U201 : BUF_X1 port map( A => positive_inputs_7_14_port, Z => n168);
   U202 : BUF_X1 port map( A => positive_inputs_7_15_port, Z => n170);
   U203 : BUF_X1 port map( A => positive_inputs_7_16_port, Z => n172);
   U204 : BUF_X1 port map( A => positive_inputs_7_17_port, Z => n174);
   U205 : BUF_X1 port map( A => positive_inputs_7_18_port, Z => n176);
   U206 : BUF_X1 port map( A => positive_inputs_7_19_port, Z => n178);
   U207 : CLKBUF_X1 port map( A => negative_inputs_7_17_port, Z => n93);
   U208 : CLKBUF_X1 port map( A => negative_inputs_7_9_port, Z => n77);
   U209 : CLKBUF_X1 port map( A => negative_inputs_7_19_port, Z => n97);

end SYN_STRUCTURAL;
