
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_BOOTHMUL_1 is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_BOOTHMUL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_2046 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2046;

architecture SYN_BEHAVIORAL of FA_2046 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n6, n7, n8, n9, n10 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n10);
   U1 : OAI22_X1 port map( A1 => n6, A2 => n7, B1 => n8, B2 => n9, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n6);
   U3 : INV_X1 port map( A => A, ZN => n7);
   U5 : INV_X1 port map( A => Ci, ZN => n8);
   U6 : INV_X1 port map( A => n10, ZN => n9);
   U7 : XOR2_X1 port map( A => Ci, B => n10, Z => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_2045 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2045;

architecture SYN_BEHAVIORAL of FA_2045 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n6, n7, n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n8, ZN => n7);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n8);
   U3 : AND2_X1 port map( A1 => B, A2 => A, ZN => n6);
   U4 : AOI21_X1 port map( B1 => Ci, B2 => n7, A => n6, ZN => n2);
   U5 : INV_X1 port map( A => n2, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n8, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_2044 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2044;

architecture SYN_BEHAVIORAL of FA_2044 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n6, n7, n8 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => n8);
   U2 : INV_X1 port map( A => n8, ZN => n7);
   U3 : AND2_X1 port map( A1 => B, A2 => A, ZN => n6);
   U4 : XNOR2_X1 port map( A => Ci, B => n8, ZN => S);
   U5 : AOI21_X1 port map( B1 => Ci, B2 => n7, A => n6, ZN => n2);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_2043 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2043;

architecture SYN_BEHAVIORAL of FA_2043 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n6, n7, n8 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => n8);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => n6);
   U3 : AOI21_X1 port map( B1 => n7, B2 => Ci, A => n6, ZN => n2);
   U4 : INV_X1 port map( A => n8, ZN => n7);
   U5 : XNOR2_X1 port map( A => Ci, B => n8, ZN => S);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_2042 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2042;

architecture SYN_BEHAVIORAL of FA_2042 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n6, n7, n8, n9 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => n9);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => n6);
   U3 : AOI21_X1 port map( B1 => Ci, B2 => n8, A => n6, ZN => n7);
   U4 : INV_X1 port map( A => n7, ZN => Co);
   U5 : INV_X1 port map( A => n9, ZN => n8);
   U6 : XNOR2_X1 port map( A => Ci, B => n9, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_2041 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2041;

architecture SYN_BEHAVIORAL of FA_2041 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n6, n7, n8 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => n8);
   U2 : XNOR2_X1 port map( A => Ci, B => n8, ZN => S);
   U3 : AND2_X1 port map( A1 => B, A2 => A, ZN => n6);
   U4 : AOI21_X1 port map( B1 => n7, B2 => Ci, A => n6, ZN => n2);
   U5 : INV_X1 port map( A => n8, ZN => n7);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_2040 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2040;

architecture SYN_BEHAVIORAL of FA_2040 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);
   U1 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n7, B2 => Ci, ZN => n8);
   U3 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_2039 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2039;

architecture SYN_BEHAVIORAL of FA_2039 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);
   U1 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : INV_X1 port map( A => n8, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n7, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_2038 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2038;

architecture SYN_BEHAVIORAL of FA_2038 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);
   U1 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U3 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_2037 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2037;

architecture SYN_BEHAVIORAL of FA_2037 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X2
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);
   U1 : XOR2_X2 port map( A => Ci, B => n7, Z => S);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n7, B2 => Ci, ZN => n8);
   U3 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_2036 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2036;

architecture SYN_BEHAVIORAL of FA_2036 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);
   U1 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : INV_X1 port map( A => n8, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n7, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_2035 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2035;

architecture SYN_BEHAVIORAL of FA_2035 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);
   U1 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U3 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_2034 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2034;

architecture SYN_BEHAVIORAL of FA_2034 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);
   U1 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : INV_X1 port map( A => n8, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n7, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_2033 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2033;

architecture SYN_BEHAVIORAL of FA_2033 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);
   U1 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U3 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_2032 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2032;

architecture SYN_BEHAVIORAL of FA_2032 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);
   U1 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n7, B2 => Ci, ZN => n8);
   U3 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_2031 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2031;

architecture SYN_BEHAVIORAL of FA_2031 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);
   U1 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : INV_X1 port map( A => n8, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n7, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_2030 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2030;

architecture SYN_BEHAVIORAL of FA_2030 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n6, n7, n8, n9, n11 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : OAI22_X1 port map( A1 => n6, A2 => n7, B1 => n8, B2 => n9, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n6);
   U3 : INV_X1 port map( A => A, ZN => n7);
   U5 : INV_X1 port map( A => n11, ZN => n8);
   U6 : INV_X1 port map( A => Ci, ZN => n9);
   U7 : XOR2_X1 port map( A => Ci, B => n11, Z => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_2029 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2029;

architecture SYN_BEHAVIORAL of FA_2029 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n6, n7, n8, n9, n11 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : OAI22_X1 port map( A1 => n6, A2 => n7, B1 => n8, B2 => n9, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n6);
   U3 : INV_X1 port map( A => A, ZN => n7);
   U5 : INV_X1 port map( A => n11, ZN => n8);
   U6 : INV_X1 port map( A => Ci, ZN => n9);
   U7 : XOR2_X1 port map( A => Ci, B => n11, Z => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_2028 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2028;

architecture SYN_BEHAVIORAL of FA_2028 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n6, n7, n8, n9, n11 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U2 : OAI22_X1 port map( A1 => n6, A2 => n7, B1 => n8, B2 => n9, ZN => Co);
   U3 : INV_X1 port map( A => B, ZN => n6);
   U5 : INV_X1 port map( A => A, ZN => n7);
   U6 : INV_X1 port map( A => Ci, ZN => n8);
   U7 : INV_X1 port map( A => n11, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_2027 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2027;

architecture SYN_BEHAVIORAL of FA_2027 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);
   U1 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U3 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_2026 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2026;

architecture SYN_BEHAVIORAL of FA_2026 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);
   U1 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : INV_X1 port map( A => n8, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n7, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_2025 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2025;

architecture SYN_BEHAVIORAL of FA_2025 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);
   U1 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n7, B2 => Ci, ZN => n8);
   U3 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_2024 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2024;

architecture SYN_BEHAVIORAL of FA_2024 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);
   U1 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : INV_X1 port map( A => n8, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n7, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_2023 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2023;

architecture SYN_BEHAVIORAL of FA_2023 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);
   U1 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U3 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_2022 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2022;

architecture SYN_BEHAVIORAL of FA_2022 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);
   U1 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n7, B2 => Ci, ZN => n8);
   U3 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_2021 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2021;

architecture SYN_BEHAVIORAL of FA_2021 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);
   U1 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : INV_X1 port map( A => n8, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n7, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_2020 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2020;

architecture SYN_BEHAVIORAL of FA_2020 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);
   U1 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n7, B2 => Ci, ZN => n8);
   U3 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_2019 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2019;

architecture SYN_BEHAVIORAL of FA_2019 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);
   U1 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : INV_X1 port map( A => n8, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n7, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_2018 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2018;

architecture SYN_BEHAVIORAL of FA_2018 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);
   U1 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U3 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_2017 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2017;

architecture SYN_BEHAVIORAL of FA_2017 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);
   U1 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n7, B2 => Ci, ZN => n8);
   U3 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_2016 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2016;

architecture SYN_BEHAVIORAL of FA_2016 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);
   U1 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : INV_X1 port map( A => n8, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n7, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_2015 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2015;

architecture SYN_BEHAVIORAL of FA_2015 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n7, B2 => Ci, ZN => n8);
   U2 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_2014 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2014;

architecture SYN_BEHAVIORAL of FA_2014 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);
   U1 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : INV_X1 port map( A => n8, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_2013 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2013;

architecture SYN_BEHAVIORAL of FA_2013 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n6, n8, n9 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n8);
   U1 : CLKBUF_X1 port map( A => Ci, Z => n6);
   U2 : XOR2_X1 port map( A => n6, B => n8, Z => S);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n8, ZN => n9);
   U5 : INV_X1 port map( A => n9, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_2012 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2012;

architecture SYN_BEHAVIORAL of FA_2012 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);
   U1 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : INV_X1 port map( A => n8, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n7, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_2011 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2011;

architecture SYN_BEHAVIORAL of FA_2011 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);
   U1 : INV_X1 port map( A => n8, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n7, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_2009 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2009;

architecture SYN_BEHAVIORAL of FA_2009 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);
   U1 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U3 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_2008 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2008;

architecture SYN_BEHAVIORAL of FA_2008 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);
   U1 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : INV_X1 port map( A => n8, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_2007 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2007;

architecture SYN_BEHAVIORAL of FA_2007 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n7, n8 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);
   U1 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n7, B2 => Ci, ZN => n8);
   U3 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_2005 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2005;

architecture SYN_BEHAVIORAL of FA_2005 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X2 port map( A => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => n5, ZN => n4);
   U3 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_2004 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2004;

architecture SYN_BEHAVIORAL of FA_2004 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : XNOR2_X1 port map( A => Ci, B => n5, ZN => n4);
   U2 : INV_X2 port map( A => n4, ZN => S);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_2003 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2003;

architecture SYN_BEHAVIORAL of FA_2003 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => n5, ZN => n4);
   U3 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_2002 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2002;

architecture SYN_BEHAVIORAL of FA_2002 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X2
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : XOR2_X2 port map( A => Ci, B => n5, Z => S);
   U2 : INV_X1 port map( A => n6, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_2001 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2001;

architecture SYN_BEHAVIORAL of FA_2001 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X2
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : XOR2_X2 port map( A => Ci, B => n4, Z => S);
   U2 : INV_X1 port map( A => n5, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_2000 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2000;

architecture SYN_BEHAVIORAL of FA_2000 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X2
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : XOR2_X2 port map( A => Ci, B => n4, Z => S);
   U2 : INV_X1 port map( A => n5, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1999 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1999;

architecture SYN_BEHAVIORAL of FA_1999 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1998 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1998;

architecture SYN_BEHAVIORAL of FA_1998 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X2
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : XOR2_X2 port map( A => Ci, B => n4, Z => S);
   U2 : INV_X1 port map( A => n5, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1997 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1997;

architecture SYN_BEHAVIORAL of FA_1997 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1995 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1995;

architecture SYN_BEHAVIORAL of FA_1995 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1994 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1994;

architecture SYN_BEHAVIORAL of FA_1994 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1993 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1993;

architecture SYN_BEHAVIORAL of FA_1993 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1992 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1992;

architecture SYN_BEHAVIORAL of FA_1992 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1991 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1991;

architecture SYN_BEHAVIORAL of FA_1991 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1990 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1990;

architecture SYN_BEHAVIORAL of FA_1990 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1989 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1989;

architecture SYN_BEHAVIORAL of FA_1989 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1988 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1988;

architecture SYN_BEHAVIORAL of FA_1988 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1987 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1987;

architecture SYN_BEHAVIORAL of FA_1987 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1986 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1986;

architecture SYN_BEHAVIORAL of FA_1986 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1985 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1985;

architecture SYN_BEHAVIORAL of FA_1985 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1984 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1984;

architecture SYN_BEHAVIORAL of FA_1984 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1983 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1983;

architecture SYN_BEHAVIORAL of FA_1983 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1982 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1982;

architecture SYN_BEHAVIORAL of FA_1982 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1981 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1981;

architecture SYN_BEHAVIORAL of FA_1981 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal net67860, n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => net67860, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);
   U2 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => n5, Z => net67860);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1980 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1980;

architecture SYN_BEHAVIORAL of FA_1980 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal net66847, n2, n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => net66847, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : CLKBUF_X1 port map( A => A, Z => n4);
   U2 : BUF_X1 port map( A => Ci, Z => net66847);
   U5 : AOI22_X1 port map( A1 => B, A2 => n4, B1 => Ci, B2 => n5, ZN => n2);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1979 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1979;

architecture SYN_BEHAVIORAL of FA_1979 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n8);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n5, B1 => n6, B2 => n7, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U5 : INV_X1 port map( A => A, ZN => n5);
   U6 : INV_X1 port map( A => Ci, ZN => n6);
   U7 : INV_X1 port map( A => n8, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1978 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1978;

architecture SYN_BEHAVIORAL of FA_1978 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => n4);
   U2 : AOI21_X1 port map( B1 => Ci, B2 => n6, A => n4, ZN => n2);
   U3 : INV_X1 port map( A => n2, ZN => Co);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n6);
   U5 : XNOR2_X1 port map( A => Ci, B => n5, ZN => S);
   U6 : XNOR2_X1 port map( A => A, B => B, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1977 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1977;

architecture SYN_BEHAVIORAL of FA_1977 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U2 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1976 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1976;

architecture SYN_BEHAVIORAL of FA_1976 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1975 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1975;

architecture SYN_BEHAVIORAL of FA_1975 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1974 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1974;

architecture SYN_BEHAVIORAL of FA_1974 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U1 : NAND2_X1 port map( A1 => A, A2 => n5, ZN => n6);
   U2 : NAND2_X1 port map( A1 => n4, A2 => B, ZN => n7);
   U4 : NAND2_X1 port map( A1 => n6, A2 => n7, ZN => n8);
   U5 : INV_X1 port map( A => A, ZN => n4);
   U6 : INV_X1 port map( A => B, ZN => n5);
   U7 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n8, ZN => n9);
   U8 : INV_X1 port map( A => n9, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1973 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1973;

architecture SYN_BEHAVIORAL of FA_1973 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n8);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n5, B1 => n6, B2 => n7, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U5 : INV_X1 port map( A => A, ZN => n5);
   U6 : INV_X1 port map( A => Ci, ZN => n6);
   U7 : INV_X1 port map( A => n8, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1972 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1972;

architecture SYN_BEHAVIORAL of FA_1972 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1971 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1971;

architecture SYN_BEHAVIORAL of FA_1971 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1970 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1970;

architecture SYN_BEHAVIORAL of FA_1970 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U2 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1969 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1969;

architecture SYN_BEHAVIORAL of FA_1969 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1968 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1968;

architecture SYN_BEHAVIORAL of FA_1968 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1967 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1967;

architecture SYN_BEHAVIORAL of FA_1967 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1966 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1966;

architecture SYN_BEHAVIORAL of FA_1966 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U2 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1965 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1965;

architecture SYN_BEHAVIORAL of FA_1965 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1964 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1964;

architecture SYN_BEHAVIORAL of FA_1964 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n8);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n5, B1 => n6, B2 => n7, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U5 : INV_X1 port map( A => A, ZN => n5);
   U6 : INV_X1 port map( A => Ci, ZN => n6);
   U7 : INV_X1 port map( A => n8, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1963 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1963;

architecture SYN_BEHAVIORAL of FA_1963 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n8);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n5, B1 => n6, B2 => n7, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U5 : INV_X1 port map( A => A, ZN => n5);
   U6 : INV_X1 port map( A => Ci, ZN => n6);
   U7 : INV_X1 port map( A => n8, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1962 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1962;

architecture SYN_BEHAVIORAL of FA_1962 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n8);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n5, B1 => n6, B2 => n7, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U5 : INV_X1 port map( A => A, ZN => n5);
   U6 : INV_X1 port map( A => Ci, ZN => n6);
   U7 : INV_X1 port map( A => n8, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1961 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1961;

architecture SYN_BEHAVIORAL of FA_1961 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1960 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1960;

architecture SYN_BEHAVIORAL of FA_1960 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1959 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1959;

architecture SYN_BEHAVIORAL of FA_1959 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1958 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1958;

architecture SYN_BEHAVIORAL of FA_1958 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1957 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1957;

architecture SYN_BEHAVIORAL of FA_1957 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1956 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1956;

architecture SYN_BEHAVIORAL of FA_1956 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1955 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1955;

architecture SYN_BEHAVIORAL of FA_1955 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1954 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1954;

architecture SYN_BEHAVIORAL of FA_1954 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1953 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1953;

architecture SYN_BEHAVIORAL of FA_1953 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1952 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1952;

architecture SYN_BEHAVIORAL of FA_1952 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1951 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1951;

architecture SYN_BEHAVIORAL of FA_1951 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1950 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1950;

architecture SYN_BEHAVIORAL of FA_1950 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1949 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1949;

architecture SYN_BEHAVIORAL of FA_1949 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1948 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1948;

architecture SYN_BEHAVIORAL of FA_1948 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1947 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1947;

architecture SYN_BEHAVIORAL of FA_1947 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1946 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1946;

architecture SYN_BEHAVIORAL of FA_1946 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n8);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n5, B1 => n6, B2 => n7, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U5 : INV_X1 port map( A => A, ZN => n5);
   U6 : INV_X1 port map( A => n8, ZN => n6);
   U7 : INV_X1 port map( A => Ci, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1945 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1945;

architecture SYN_BEHAVIORAL of FA_1945 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1944 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1944;

architecture SYN_BEHAVIORAL of FA_1944 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1943 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1943;

architecture SYN_BEHAVIORAL of FA_1943 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U2 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1942 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1942;

architecture SYN_BEHAVIORAL of FA_1942 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1941 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1941;

architecture SYN_BEHAVIORAL of FA_1941 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n8);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n5, B1 => n6, B2 => n7, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U5 : INV_X1 port map( A => A, ZN => n5);
   U6 : INV_X1 port map( A => n8, ZN => n6);
   U7 : INV_X1 port map( A => Ci, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1940 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1940;

architecture SYN_BEHAVIORAL of FA_1940 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1939 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1939;

architecture SYN_BEHAVIORAL of FA_1939 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1938 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1938;

architecture SYN_BEHAVIORAL of FA_1938 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1937 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1937;

architecture SYN_BEHAVIORAL of FA_1937 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1936 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1936;

architecture SYN_BEHAVIORAL of FA_1936 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1935 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1935;

architecture SYN_BEHAVIORAL of FA_1935 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1934 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1934;

architecture SYN_BEHAVIORAL of FA_1934 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1933 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1933;

architecture SYN_BEHAVIORAL of FA_1933 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1932 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1932;

architecture SYN_BEHAVIORAL of FA_1932 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1931 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1931;

architecture SYN_BEHAVIORAL of FA_1931 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1930 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1930;

architecture SYN_BEHAVIORAL of FA_1930 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1929 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1929;

architecture SYN_BEHAVIORAL of FA_1929 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1928 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1928;

architecture SYN_BEHAVIORAL of FA_1928 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1927 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1927;

architecture SYN_BEHAVIORAL of FA_1927 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1926 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1926;

architecture SYN_BEHAVIORAL of FA_1926 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1925 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1925;

architecture SYN_BEHAVIORAL of FA_1925 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1924 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1924;

architecture SYN_BEHAVIORAL of FA_1924 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1923 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1923;

architecture SYN_BEHAVIORAL of FA_1923 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1922 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1922;

architecture SYN_BEHAVIORAL of FA_1922 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1921 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1921;

architecture SYN_BEHAVIORAL of FA_1921 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1920 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1920;

architecture SYN_BEHAVIORAL of FA_1920 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1919 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1919;

architecture SYN_BEHAVIORAL of FA_1919 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1918 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1918;

architecture SYN_BEHAVIORAL of FA_1918 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1917 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1917;

architecture SYN_BEHAVIORAL of FA_1917 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1916 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1916;

architecture SYN_BEHAVIORAL of FA_1916 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1915 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1915;

architecture SYN_BEHAVIORAL of FA_1915 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n9, n10 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n9, B => n6, ZN => S);
   U2 : AOI22_X1 port map( A1 => n8, A2 => n7, B1 => n4, B2 => n5, ZN => Co);
   U3 : INV_X1 port map( A => A, ZN => n4);
   U4 : INV_X1 port map( A => B, ZN => n5);
   U5 : INV_X1 port map( A => Ci, ZN => n8);
   U6 : INV_X1 port map( A => n10, ZN => n9);
   U7 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U8 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n7);
   U9 : CLKBUF_X1 port map( A => n8, Z => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1914 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1914;

architecture SYN_BEHAVIORAL of FA_1914 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U2 : AOI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n6);
   U4 : NOR2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U5 : NOR2_X1 port map( A1 => B, A2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1913 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1913;

architecture SYN_BEHAVIORAL of FA_1913 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => Ci, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U1 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => n4, B2 => Ci, ZN => n2);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1912 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1912;

architecture SYN_BEHAVIORAL of FA_1912 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U2 : INV_X1 port map( A => n4, ZN => Co);
   U4 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);
   U5 : INV_X1 port map( A => A, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1911 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1911;

architecture SYN_BEHAVIORAL of FA_1911 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U2 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U4 : INV_X1 port map( A => A, ZN => n5);
   U5 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1910 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1910;

architecture SYN_BEHAVIORAL of FA_1910 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1909 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1909;

architecture SYN_BEHAVIORAL of FA_1909 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1908 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1908;

architecture SYN_BEHAVIORAL of FA_1908 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1907 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1907;

architecture SYN_BEHAVIORAL of FA_1907 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1906 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1906;

architecture SYN_BEHAVIORAL of FA_1906 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n9);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : OAI22_X1 port map( A1 => n5, A2 => n6, B1 => n7, B2 => n8, ZN => Co);
   U5 : INV_X1 port map( A => n4, ZN => n5);
   U6 : INV_X1 port map( A => A, ZN => n6);
   U7 : INV_X1 port map( A => Ci, ZN => n7);
   U8 : INV_X1 port map( A => n9, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1905 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1905;

architecture SYN_BEHAVIORAL of FA_1905 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n5, B => Ci, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1904 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1904;

architecture SYN_BEHAVIORAL of FA_1904 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => Ci, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1903 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1903;

architecture SYN_BEHAVIORAL of FA_1903 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1902 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1902;

architecture SYN_BEHAVIORAL of FA_1902 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1901 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1901;

architecture SYN_BEHAVIORAL of FA_1901 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1900 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1900;

architecture SYN_BEHAVIORAL of FA_1900 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1899 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1899;

architecture SYN_BEHAVIORAL of FA_1899 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => Ci, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1898 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1898;

architecture SYN_BEHAVIORAL of FA_1898 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n7, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : INV_X1 port map( A => n8, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n7);
   U7 : XNOR2_X1 port map( A => B, B => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1897 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1897;

architecture SYN_BEHAVIORAL of FA_1897 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1896 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1896;

architecture SYN_BEHAVIORAL of FA_1896 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1895 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1895;

architecture SYN_BEHAVIORAL of FA_1895 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n7, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : INV_X1 port map( A => n8, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n7);
   U7 : XNOR2_X1 port map( A => n7, B => B, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1894 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1894;

architecture SYN_BEHAVIORAL of FA_1894 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1893 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1893;

architecture SYN_BEHAVIORAL of FA_1893 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n7, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : INV_X1 port map( A => n8, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n7);
   U7 : XNOR2_X1 port map( A => n7, B => B, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1892 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1892;

architecture SYN_BEHAVIORAL of FA_1892 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1891 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1891;

architecture SYN_BEHAVIORAL of FA_1891 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1890 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1890;

architecture SYN_BEHAVIORAL of FA_1890 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1889 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1889;

architecture SYN_BEHAVIORAL of FA_1889 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1888 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1888;

architecture SYN_BEHAVIORAL of FA_1888 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1887 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1887;

architecture SYN_BEHAVIORAL of FA_1887 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1886 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1886;

architecture SYN_BEHAVIORAL of FA_1886 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1885 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1885;

architecture SYN_BEHAVIORAL of FA_1885 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1884 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1884;

architecture SYN_BEHAVIORAL of FA_1884 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1883 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1883;

architecture SYN_BEHAVIORAL of FA_1883 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1882 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1882;

architecture SYN_BEHAVIORAL of FA_1882 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1881 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1881;

architecture SYN_BEHAVIORAL of FA_1881 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1880 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1880;

architecture SYN_BEHAVIORAL of FA_1880 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1879 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1879;

architecture SYN_BEHAVIORAL of FA_1879 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U2 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1878 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1878;

architecture SYN_BEHAVIORAL of FA_1878 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1877 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1877;

architecture SYN_BEHAVIORAL of FA_1877 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1876 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1876;

architecture SYN_BEHAVIORAL of FA_1876 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n8);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n5, B1 => n6, B2 => n7, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U5 : INV_X1 port map( A => A, ZN => n5);
   U6 : INV_X1 port map( A => n8, ZN => n6);
   U7 : INV_X1 port map( A => Ci, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1875 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1875;

architecture SYN_BEHAVIORAL of FA_1875 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1874 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1874;

architecture SYN_BEHAVIORAL of FA_1874 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1873 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1873;

architecture SYN_BEHAVIORAL of FA_1873 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1872 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1872;

architecture SYN_BEHAVIORAL of FA_1872 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1871 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1871;

architecture SYN_BEHAVIORAL of FA_1871 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n7, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : INV_X1 port map( A => n8, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n7);
   U7 : XNOR2_X1 port map( A => n7, B => B, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1870 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1870;

architecture SYN_BEHAVIORAL of FA_1870 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1869 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1869;

architecture SYN_BEHAVIORAL of FA_1869 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1868 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1868;

architecture SYN_BEHAVIORAL of FA_1868 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1867 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1867;

architecture SYN_BEHAVIORAL of FA_1867 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1866 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1866;

architecture SYN_BEHAVIORAL of FA_1866 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1865 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1865;

architecture SYN_BEHAVIORAL of FA_1865 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1864 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1864;

architecture SYN_BEHAVIORAL of FA_1864 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1863 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1863;

architecture SYN_BEHAVIORAL of FA_1863 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1862 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1862;

architecture SYN_BEHAVIORAL of FA_1862 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1861 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1861;

architecture SYN_BEHAVIORAL of FA_1861 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1860 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1860;

architecture SYN_BEHAVIORAL of FA_1860 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1859 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1859;

architecture SYN_BEHAVIORAL of FA_1859 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1858 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1858;

architecture SYN_BEHAVIORAL of FA_1858 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1857 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1857;

architecture SYN_BEHAVIORAL of FA_1857 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1856 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1856;

architecture SYN_BEHAVIORAL of FA_1856 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1855 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1855;

architecture SYN_BEHAVIORAL of FA_1855 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1854 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1854;

architecture SYN_BEHAVIORAL of FA_1854 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1853 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1853;

architecture SYN_BEHAVIORAL of FA_1853 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1852 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1852;

architecture SYN_BEHAVIORAL of FA_1852 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1851 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1851;

architecture SYN_BEHAVIORAL of FA_1851 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1850 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1850;

architecture SYN_BEHAVIORAL of FA_1850 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1849 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1849;

architecture SYN_BEHAVIORAL of FA_1849 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : AOI22_X1 port map( A1 => A, A2 => n4, B1 => n6, B2 => Ci, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1848 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1848;

architecture SYN_BEHAVIORAL of FA_1848 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : CLKBUF_X1 port map( A => n7, Z => n4);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n7);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);
   U7 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1847 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1847;

architecture SYN_BEHAVIORAL of FA_1847 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U4 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1846 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1846;

architecture SYN_BEHAVIORAL of FA_1846 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1845 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1845;

architecture SYN_BEHAVIORAL of FA_1845 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => n5, B2 => Ci, ZN => n4);
   U2 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1844 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1844;

architecture SYN_BEHAVIORAL of FA_1844 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U5 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1843 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1843;

architecture SYN_BEHAVIORAL of FA_1843 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1842 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1842;

architecture SYN_BEHAVIORAL of FA_1842 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1841 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1841;

architecture SYN_BEHAVIORAL of FA_1841 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n5);
   U5 : INV_X1 port map( A => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1840 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1840;

architecture SYN_BEHAVIORAL of FA_1840 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => n6, B => B, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1839 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1839;

architecture SYN_BEHAVIORAL of FA_1839 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U2 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1838 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1838;

architecture SYN_BEHAVIORAL of FA_1838 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1837 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1837;

architecture SYN_BEHAVIORAL of FA_1837 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n7, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : INV_X1 port map( A => n8, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n7);
   U7 : XNOR2_X1 port map( A => B, B => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1836 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1836;

architecture SYN_BEHAVIORAL of FA_1836 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1835 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1835;

architecture SYN_BEHAVIORAL of FA_1835 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1834 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1834;

architecture SYN_BEHAVIORAL of FA_1834 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1833 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1833;

architecture SYN_BEHAVIORAL of FA_1833 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n7, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : INV_X1 port map( A => n8, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n7);
   U7 : XNOR2_X1 port map( A => B, B => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1832 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1832;

architecture SYN_BEHAVIORAL of FA_1832 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1831 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1831;

architecture SYN_BEHAVIORAL of FA_1831 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n7, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : INV_X1 port map( A => n8, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n7);
   U7 : XNOR2_X1 port map( A => B, B => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1830 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1830;

architecture SYN_BEHAVIORAL of FA_1830 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U3 : XOR2_X1 port map( A => B, B => n6, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1829 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1829;

architecture SYN_BEHAVIORAL of FA_1829 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n7, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : INV_X1 port map( A => n8, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n7);
   U7 : XNOR2_X1 port map( A => n7, B => B, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1828 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1828;

architecture SYN_BEHAVIORAL of FA_1828 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1827 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1827;

architecture SYN_BEHAVIORAL of FA_1827 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1826 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1826;

architecture SYN_BEHAVIORAL of FA_1826 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n7, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : INV_X1 port map( A => n8, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n7);
   U7 : XNOR2_X1 port map( A => B, B => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1825 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1825;

architecture SYN_BEHAVIORAL of FA_1825 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1824 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1824;

architecture SYN_BEHAVIORAL of FA_1824 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1823 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1823;

architecture SYN_BEHAVIORAL of FA_1823 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1822 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1822;

architecture SYN_BEHAVIORAL of FA_1822 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1821 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1821;

architecture SYN_BEHAVIORAL of FA_1821 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1820 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1820;

architecture SYN_BEHAVIORAL of FA_1820 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1819 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1819;

architecture SYN_BEHAVIORAL of FA_1819 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1818 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1818;

architecture SYN_BEHAVIORAL of FA_1818 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1817 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1817;

architecture SYN_BEHAVIORAL of FA_1817 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1816 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1816;

architecture SYN_BEHAVIORAL of FA_1816 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1815 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1815;

architecture SYN_BEHAVIORAL of FA_1815 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n2);
   U5 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1814 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1814;

architecture SYN_BEHAVIORAL of FA_1814 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n4);
   U2 : INV_X1 port map( A => n4, ZN => Co);
   U4 : INV_X1 port map( A => A, ZN => n5);
   U5 : XNOR2_X1 port map( A => n5, B => B, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1813 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1813;

architecture SYN_BEHAVIORAL of FA_1813 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1812 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1812;

architecture SYN_BEHAVIORAL of FA_1812 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n9, n10 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U1 : NAND2_X1 port map( A1 => A, A2 => n5, ZN => n6);
   U2 : NAND2_X1 port map( A1 => B, A2 => n4, ZN => n7);
   U4 : NAND2_X1 port map( A1 => n6, A2 => n7, ZN => n9);
   U5 : INV_X1 port map( A => A, ZN => n4);
   U6 : INV_X1 port map( A => B, ZN => n5);
   U7 : CLKBUF_X1 port map( A => B, Z => n8);
   U8 : INV_X1 port map( A => n10, ZN => Co);
   U9 : AOI22_X1 port map( A1 => n8, A2 => A, B1 => Ci, B2 => n9, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1811 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1811;

architecture SYN_BEHAVIORAL of FA_1811 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1810 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1810;

architecture SYN_BEHAVIORAL of FA_1810 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n7, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : INV_X1 port map( A => n8, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n7);
   U7 : XNOR2_X1 port map( A => n7, B => B, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1809 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1809;

architecture SYN_BEHAVIORAL of FA_1809 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1808 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1808;

architecture SYN_BEHAVIORAL of FA_1808 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1807 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1807;

architecture SYN_BEHAVIORAL of FA_1807 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1806 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1806;

architecture SYN_BEHAVIORAL of FA_1806 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1805 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1805;

architecture SYN_BEHAVIORAL of FA_1805 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1804 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1804;

architecture SYN_BEHAVIORAL of FA_1804 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1803 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1803;

architecture SYN_BEHAVIORAL of FA_1803 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1802 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1802;

architecture SYN_BEHAVIORAL of FA_1802 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n4);
   U2 : INV_X1 port map( A => n4, ZN => Co);
   U4 : INV_X1 port map( A => A, ZN => n5);
   U5 : XNOR2_X1 port map( A => n5, B => B, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1801 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1801;

architecture SYN_BEHAVIORAL of FA_1801 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1800 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1800;

architecture SYN_BEHAVIORAL of FA_1800 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1799 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1799;

architecture SYN_BEHAVIORAL of FA_1799 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1798 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1798;

architecture SYN_BEHAVIORAL of FA_1798 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1797 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1797;

architecture SYN_BEHAVIORAL of FA_1797 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1796 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1796;

architecture SYN_BEHAVIORAL of FA_1796 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1795 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1795;

architecture SYN_BEHAVIORAL of FA_1795 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1794 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1794;

architecture SYN_BEHAVIORAL of FA_1794 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1793 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1793;

architecture SYN_BEHAVIORAL of FA_1793 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1792 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1792;

architecture SYN_BEHAVIORAL of FA_1792 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1791 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1791;

architecture SYN_BEHAVIORAL of FA_1791 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1790 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1790;

architecture SYN_BEHAVIORAL of FA_1790 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1789 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1789;

architecture SYN_BEHAVIORAL of FA_1789 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1788 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1788;

architecture SYN_BEHAVIORAL of FA_1788 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1787 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1787;

architecture SYN_BEHAVIORAL of FA_1787 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1786 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1786;

architecture SYN_BEHAVIORAL of FA_1786 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1785 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1785;

architecture SYN_BEHAVIORAL of FA_1785 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1784 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1784;

architecture SYN_BEHAVIORAL of FA_1784 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1783 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1783;

architecture SYN_BEHAVIORAL of FA_1783 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : CLKBUF_X1 port map( A => n7, Z => n5);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n7);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n7, B2 => Ci, ZN => n8);
   U7 : INV_X1 port map( A => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1782 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1782;

architecture SYN_BEHAVIORAL of FA_1782 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n6, B2 => Ci, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1781 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1781;

architecture SYN_BEHAVIORAL of FA_1781 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n6, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n6, B2 => Ci, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1780 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1780;

architecture SYN_BEHAVIORAL of FA_1780 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : XNOR2_X1 port map( A => B, B => n6, ZN => n4);
   U4 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U5 : CLKBUF_X1 port map( A => B, Z => n5);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1779 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1779;

architecture SYN_BEHAVIORAL of FA_1779 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1778 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1778;

architecture SYN_BEHAVIORAL of FA_1778 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1777 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1777;

architecture SYN_BEHAVIORAL of FA_1777 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1776 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1776;

architecture SYN_BEHAVIORAL of FA_1776 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1775 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1775;

architecture SYN_BEHAVIORAL of FA_1775 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : INV_X1 port map( A => n2, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1774 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1774;

architecture SYN_BEHAVIORAL of FA_1774 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1773 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1773;

architecture SYN_BEHAVIORAL of FA_1773 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n8, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : INV_X1 port map( A => n7, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n8);
   U7 : XNOR2_X1 port map( A => B, B => n8, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1772 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1772;

architecture SYN_BEHAVIORAL of FA_1772 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U5 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1771 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1771;

architecture SYN_BEHAVIORAL of FA_1771 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U2 : INV_X1 port map( A => n4, ZN => Co);
   U4 : INV_X1 port map( A => A, ZN => n6);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1770 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1770;

architecture SYN_BEHAVIORAL of FA_1770 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1769 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1769;

architecture SYN_BEHAVIORAL of FA_1769 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1768 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1768;

architecture SYN_BEHAVIORAL of FA_1768 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1767 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1767;

architecture SYN_BEHAVIORAL of FA_1767 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1766 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1766;

architecture SYN_BEHAVIORAL of FA_1766 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n8, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : INV_X1 port map( A => n7, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n8);
   U7 : XNOR2_X1 port map( A => B, B => n8, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1765 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1765;

architecture SYN_BEHAVIORAL of FA_1765 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1764 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1764;

architecture SYN_BEHAVIORAL of FA_1764 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1763 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1763;

architecture SYN_BEHAVIORAL of FA_1763 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1762 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1762;

architecture SYN_BEHAVIORAL of FA_1762 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n8, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : INV_X1 port map( A => n7, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n8);
   U7 : XNOR2_X1 port map( A => B, B => n8, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1761 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1761;

architecture SYN_BEHAVIORAL of FA_1761 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U5 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1760 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1760;

architecture SYN_BEHAVIORAL of FA_1760 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1759 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1759;

architecture SYN_BEHAVIORAL of FA_1759 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n8, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : INV_X1 port map( A => n7, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n8);
   U7 : XNOR2_X1 port map( A => n8, B => B, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1758 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1758;

architecture SYN_BEHAVIORAL of FA_1758 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n8, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : INV_X1 port map( A => n7, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n8);
   U7 : XNOR2_X1 port map( A => n8, B => B, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1757 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1757;

architecture SYN_BEHAVIORAL of FA_1757 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1756 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1756;

architecture SYN_BEHAVIORAL of FA_1756 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n8, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : INV_X1 port map( A => n7, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n8);
   U7 : XNOR2_X1 port map( A => n8, B => B, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1755 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1755;

architecture SYN_BEHAVIORAL of FA_1755 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n8, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : INV_X1 port map( A => n7, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n8);
   U7 : XNOR2_X1 port map( A => B, B => n8, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1754 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1754;

architecture SYN_BEHAVIORAL of FA_1754 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1753 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1753;

architecture SYN_BEHAVIORAL of FA_1753 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1752 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1752;

architecture SYN_BEHAVIORAL of FA_1752 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1751 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1751;

architecture SYN_BEHAVIORAL of FA_1751 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U5 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1750 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1750;

architecture SYN_BEHAVIORAL of FA_1750 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1749 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1749;

architecture SYN_BEHAVIORAL of FA_1749 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n7, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : INV_X1 port map( A => n8, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n7);
   U7 : XNOR2_X1 port map( A => B, B => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1748 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1748;

architecture SYN_BEHAVIORAL of FA_1748 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => n5, B => B, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1747 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1747;

architecture SYN_BEHAVIORAL of FA_1747 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => n5, B => B, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1746 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1746;

architecture SYN_BEHAVIORAL of FA_1746 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n7, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : INV_X1 port map( A => n8, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n7);
   U7 : XNOR2_X1 port map( A => B, B => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1745 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1745;

architecture SYN_BEHAVIORAL of FA_1745 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1744 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1744;

architecture SYN_BEHAVIORAL of FA_1744 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1743 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1743;

architecture SYN_BEHAVIORAL of FA_1743 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1742 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1742;

architecture SYN_BEHAVIORAL of FA_1742 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1741 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1741;

architecture SYN_BEHAVIORAL of FA_1741 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n7, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => n8, ZN => n5);
   U5 : INV_X1 port map( A => Ci, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n7);
   U7 : XNOR2_X1 port map( A => B, B => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1740 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1740;

architecture SYN_BEHAVIORAL of FA_1740 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n4);
   U2 : INV_X1 port map( A => n4, ZN => Co);
   U4 : INV_X1 port map( A => A, ZN => n5);
   U5 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1739 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1739;

architecture SYN_BEHAVIORAL of FA_1739 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => n5, B => B, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1738 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1738;

architecture SYN_BEHAVIORAL of FA_1738 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => n5, B => B, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1737 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1737;

architecture SYN_BEHAVIORAL of FA_1737 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1736 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1736;

architecture SYN_BEHAVIORAL of FA_1736 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1735 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1735;

architecture SYN_BEHAVIORAL of FA_1735 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1734 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1734;

architecture SYN_BEHAVIORAL of FA_1734 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1733 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1733;

architecture SYN_BEHAVIORAL of FA_1733 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1732 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1732;

architecture SYN_BEHAVIORAL of FA_1732 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1731 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1731;

architecture SYN_BEHAVIORAL of FA_1731 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1730 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1730;

architecture SYN_BEHAVIORAL of FA_1730 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1729 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1729;

architecture SYN_BEHAVIORAL of FA_1729 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1728 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1728;

architecture SYN_BEHAVIORAL of FA_1728 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1727 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1727;

architecture SYN_BEHAVIORAL of FA_1727 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1726 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1726;

architecture SYN_BEHAVIORAL of FA_1726 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1725 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1725;

architecture SYN_BEHAVIORAL of FA_1725 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1724 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1724;

architecture SYN_BEHAVIORAL of FA_1724 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1723 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1723;

architecture SYN_BEHAVIORAL of FA_1723 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1722 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1722;

architecture SYN_BEHAVIORAL of FA_1722 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1721 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1721;

architecture SYN_BEHAVIORAL of FA_1721 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1720 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1720;

architecture SYN_BEHAVIORAL of FA_1720 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1719 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1719;

architecture SYN_BEHAVIORAL of FA_1719 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1718 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1718;

architecture SYN_BEHAVIORAL of FA_1718 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1717 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1717;

architecture SYN_BEHAVIORAL of FA_1717 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n6, B2 => Ci, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1716 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1716;

architecture SYN_BEHAVIORAL of FA_1716 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1715 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1715;

architecture SYN_BEHAVIORAL of FA_1715 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1714 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1714;

architecture SYN_BEHAVIORAL of FA_1714 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1713 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1713;

architecture SYN_BEHAVIORAL of FA_1713 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1712 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1712;

architecture SYN_BEHAVIORAL of FA_1712 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1711 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1711;

architecture SYN_BEHAVIORAL of FA_1711 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : OAI22_X1 port map( A1 => n5, A2 => n9, B1 => n6, B2 => n7, ZN => Co);
   U4 : INV_X1 port map( A => n4, ZN => n5);
   U5 : INV_X1 port map( A => Ci, ZN => n6);
   U6 : INV_X1 port map( A => n8, ZN => n7);
   U7 : INV_X1 port map( A => A, ZN => n9);
   U8 : XNOR2_X1 port map( A => B, B => n9, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1710 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1710;

architecture SYN_BEHAVIORAL of FA_1710 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => n6, B2 => Ci, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1709 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1709;

architecture SYN_BEHAVIORAL of FA_1709 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n6, B2 => Ci, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1708 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1708;

architecture SYN_BEHAVIORAL of FA_1708 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1707 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1707;

architecture SYN_BEHAVIORAL of FA_1707 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1706 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1706;

architecture SYN_BEHAVIORAL of FA_1706 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1705 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1705;

architecture SYN_BEHAVIORAL of FA_1705 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1704 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1704;

architecture SYN_BEHAVIORAL of FA_1704 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1703 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1703;

architecture SYN_BEHAVIORAL of FA_1703 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U1 : XOR2_X1 port map( A => B, B => n7, Z => n4);
   U2 : OAI22_X1 port map( A1 => n5, A2 => n7, B1 => n6, B2 => n4, ZN => Co);
   U4 : INV_X1 port map( A => B, ZN => n5);
   U5 : INV_X1 port map( A => Ci, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n7);
   U7 : XNOR2_X1 port map( A => B, B => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1702 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1702;

architecture SYN_BEHAVIORAL of FA_1702 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1701 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1701;

architecture SYN_BEHAVIORAL of FA_1701 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n7, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : INV_X1 port map( A => n8, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n7);
   U7 : XNOR2_X1 port map( A => B, B => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1700 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1700;

architecture SYN_BEHAVIORAL of FA_1700 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1699 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1699;

architecture SYN_BEHAVIORAL of FA_1699 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U4 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1698 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1698;

architecture SYN_BEHAVIORAL of FA_1698 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U2 : OAI22_X1 port map( A1 => n4, A2 => n7, B1 => n5, B2 => n6, ZN => Co);
   U4 : INV_X1 port map( A => B, ZN => n4);
   U5 : INV_X1 port map( A => Ci, ZN => n5);
   U6 : INV_X1 port map( A => A, ZN => n7);
   U7 : XNOR2_X1 port map( A => B, B => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1697 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1697;

architecture SYN_BEHAVIORAL of FA_1697 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U5 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1696 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1696;

architecture SYN_BEHAVIORAL of FA_1696 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1695 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1695;

architecture SYN_BEHAVIORAL of FA_1695 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n4);
   U2 : INV_X1 port map( A => n4, ZN => Co);
   U4 : INV_X1 port map( A => A, ZN => n5);
   U5 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1694 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1694;

architecture SYN_BEHAVIORAL of FA_1694 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n7, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : INV_X1 port map( A => n8, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n7);
   U7 : XNOR2_X1 port map( A => B, B => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1693 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1693;

architecture SYN_BEHAVIORAL of FA_1693 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1692 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1692;

architecture SYN_BEHAVIORAL of FA_1692 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U3 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U5 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1691 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1691;

architecture SYN_BEHAVIORAL of FA_1691 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U5 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1690 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1690;

architecture SYN_BEHAVIORAL of FA_1690 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n4);
   U2 : INV_X1 port map( A => n4, ZN => Co);
   U4 : INV_X1 port map( A => A, ZN => n5);
   U5 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1689 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1689;

architecture SYN_BEHAVIORAL of FA_1689 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1688 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1688;

architecture SYN_BEHAVIORAL of FA_1688 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1687 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1687;

architecture SYN_BEHAVIORAL of FA_1687 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U5 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1686 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1686;

architecture SYN_BEHAVIORAL of FA_1686 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1685 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1685;

architecture SYN_BEHAVIORAL of FA_1685 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n7, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : INV_X1 port map( A => n8, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n7);
   U7 : XNOR2_X1 port map( A => B, B => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1684 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1684;

architecture SYN_BEHAVIORAL of FA_1684 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1683 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1683;

architecture SYN_BEHAVIORAL of FA_1683 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1682 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1682;

architecture SYN_BEHAVIORAL of FA_1682 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n9, B => Ci, Z => S);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : OAI22_X1 port map( A1 => n5, A2 => n8, B1 => n6, B2 => n7, ZN => Co);
   U4 : INV_X1 port map( A => n4, ZN => n5);
   U5 : INV_X1 port map( A => Ci, ZN => n6);
   U6 : INV_X1 port map( A => n9, ZN => n7);
   U7 : INV_X1 port map( A => A, ZN => n8);
   U8 : XNOR2_X1 port map( A => B, B => n8, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1681 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1681;

architecture SYN_BEHAVIORAL of FA_1681 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1680 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1680;

architecture SYN_BEHAVIORAL of FA_1680 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1679 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1679;

architecture SYN_BEHAVIORAL of FA_1679 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1678 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1678;

architecture SYN_BEHAVIORAL of FA_1678 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1677 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1677;

architecture SYN_BEHAVIORAL of FA_1677 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1676 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1676;

architecture SYN_BEHAVIORAL of FA_1676 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1675 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1675;

architecture SYN_BEHAVIORAL of FA_1675 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1674 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1674;

architecture SYN_BEHAVIORAL of FA_1674 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1673 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1673;

architecture SYN_BEHAVIORAL of FA_1673 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1672 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1672;

architecture SYN_BEHAVIORAL of FA_1672 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1671 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1671;

architecture SYN_BEHAVIORAL of FA_1671 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1670 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1670;

architecture SYN_BEHAVIORAL of FA_1670 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1669 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1669;

architecture SYN_BEHAVIORAL of FA_1669 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1668 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1668;

architecture SYN_BEHAVIORAL of FA_1668 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1667 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1667;

architecture SYN_BEHAVIORAL of FA_1667 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1666 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1666;

architecture SYN_BEHAVIORAL of FA_1666 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1665 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1665;

architecture SYN_BEHAVIORAL of FA_1665 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => n6, ZN => Co);
   U2 : INV_X1 port map( A => A, ZN => n4);
   U4 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1664 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1664;

architecture SYN_BEHAVIORAL of FA_1664 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1663 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1663;

architecture SYN_BEHAVIORAL of FA_1663 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1662 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1662;

architecture SYN_BEHAVIORAL of FA_1662 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1661 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1661;

architecture SYN_BEHAVIORAL of FA_1661 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1660 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1660;

architecture SYN_BEHAVIORAL of FA_1660 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1659 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1659;

architecture SYN_BEHAVIORAL of FA_1659 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1658 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1658;

architecture SYN_BEHAVIORAL of FA_1658 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1657 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1657;

architecture SYN_BEHAVIORAL of FA_1657 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1656 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1656;

architecture SYN_BEHAVIORAL of FA_1656 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1655 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1655;

architecture SYN_BEHAVIORAL of FA_1655 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1654 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1654;

architecture SYN_BEHAVIORAL of FA_1654 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1653 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1653;

architecture SYN_BEHAVIORAL of FA_1653 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1652 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1652;

architecture SYN_BEHAVIORAL of FA_1652 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1651 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1651;

architecture SYN_BEHAVIORAL of FA_1651 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => n6, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n6, B2 => Ci, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1650 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1650;

architecture SYN_BEHAVIORAL of FA_1650 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n5, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1649 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1649;

architecture SYN_BEHAVIORAL of FA_1649 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1648 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1648;

architecture SYN_BEHAVIORAL of FA_1648 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1647 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1647;

architecture SYN_BEHAVIORAL of FA_1647 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1646 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1646;

architecture SYN_BEHAVIORAL of FA_1646 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1645 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1645;

architecture SYN_BEHAVIORAL of FA_1645 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1644 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1644;

architecture SYN_BEHAVIORAL of FA_1644 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1643 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1643;

architecture SYN_BEHAVIORAL of FA_1643 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1642 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1642;

architecture SYN_BEHAVIORAL of FA_1642 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1641 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1641;

architecture SYN_BEHAVIORAL of FA_1641 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1640 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1640;

architecture SYN_BEHAVIORAL of FA_1640 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n7, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : INV_X1 port map( A => n8, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n7);
   U7 : XNOR2_X1 port map( A => B, B => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1639 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1639;

architecture SYN_BEHAVIORAL of FA_1639 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n6, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => n6, B2 => Ci, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1638 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1638;

architecture SYN_BEHAVIORAL of FA_1638 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1637 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1637;

architecture SYN_BEHAVIORAL of FA_1637 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n9, B => Ci, Z => S);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : OAI22_X1 port map( A1 => n5, A2 => n8, B1 => n6, B2 => n7, ZN => Co);
   U4 : INV_X1 port map( A => n4, ZN => n5);
   U5 : INV_X1 port map( A => Ci, ZN => n6);
   U6 : INV_X1 port map( A => n9, ZN => n7);
   U7 : INV_X1 port map( A => A, ZN => n8);
   U8 : XNOR2_X1 port map( A => B, B => n8, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1636 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1636;

architecture SYN_BEHAVIORAL of FA_1636 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1635 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1635;

architecture SYN_BEHAVIORAL of FA_1635 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n4);
   U2 : INV_X1 port map( A => n4, ZN => Co);
   U4 : INV_X1 port map( A => A, ZN => n5);
   U5 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1634 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1634;

architecture SYN_BEHAVIORAL of FA_1634 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1633 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1633;

architecture SYN_BEHAVIORAL of FA_1633 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U5 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1632 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1632;

architecture SYN_BEHAVIORAL of FA_1632 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n7, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : INV_X1 port map( A => n8, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n7);
   U7 : XNOR2_X1 port map( A => B, B => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1631 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1631;

architecture SYN_BEHAVIORAL of FA_1631 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n7, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : INV_X1 port map( A => n8, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n7);
   U7 : XNOR2_X1 port map( A => B, B => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1630 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1630;

architecture SYN_BEHAVIORAL of FA_1630 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U4 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1629 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1629;

architecture SYN_BEHAVIORAL of FA_1629 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U4 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1628 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1628;

architecture SYN_BEHAVIORAL of FA_1628 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n7, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : INV_X1 port map( A => n8, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n7);
   U7 : XNOR2_X1 port map( A => B, B => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1627 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1627;

architecture SYN_BEHAVIORAL of FA_1627 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U5 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1626 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1626;

architecture SYN_BEHAVIORAL of FA_1626 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1625 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1625;

architecture SYN_BEHAVIORAL of FA_1625 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U4 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1624 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1624;

architecture SYN_BEHAVIORAL of FA_1624 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U4 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1623 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1623;

architecture SYN_BEHAVIORAL of FA_1623 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U5 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1622 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1622;

architecture SYN_BEHAVIORAL of FA_1622 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1621 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1621;

architecture SYN_BEHAVIORAL of FA_1621 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1620 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1620;

architecture SYN_BEHAVIORAL of FA_1620 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U4 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1619 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1619;

architecture SYN_BEHAVIORAL of FA_1619 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n4);
   U2 : INV_X1 port map( A => n4, ZN => Co);
   U4 : INV_X1 port map( A => A, ZN => n5);
   U5 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1618 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1618;

architecture SYN_BEHAVIORAL of FA_1618 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U1 : XOR2_X1 port map( A => B, B => n8, Z => n4);
   U2 : CLKBUF_X1 port map( A => B, Z => n5);
   U4 : OAI22_X1 port map( A1 => n6, A2 => n8, B1 => n7, B2 => n4, ZN => Co);
   U5 : INV_X1 port map( A => n5, ZN => n6);
   U6 : INV_X1 port map( A => Ci, ZN => n7);
   U7 : INV_X1 port map( A => A, ZN => n8);
   U8 : XNOR2_X1 port map( A => B, B => n8, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1617 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1617;

architecture SYN_BEHAVIORAL of FA_1617 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U4 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1616 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1616;

architecture SYN_BEHAVIORAL of FA_1616 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U4 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1615 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1615;

architecture SYN_BEHAVIORAL of FA_1615 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U4 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1614 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1614;

architecture SYN_BEHAVIORAL of FA_1614 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U4 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1613 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1613;

architecture SYN_BEHAVIORAL of FA_1613 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U4 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1612 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1612;

architecture SYN_BEHAVIORAL of FA_1612 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U4 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1611 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1611;

architecture SYN_BEHAVIORAL of FA_1611 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U4 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1610 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1610;

architecture SYN_BEHAVIORAL of FA_1610 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U4 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1609 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1609;

architecture SYN_BEHAVIORAL of FA_1609 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U4 : XNOR2_X1 port map( A => n4, B => B, ZN => n5);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1608 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1608;

architecture SYN_BEHAVIORAL of FA_1608 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U4 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1607 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1607;

architecture SYN_BEHAVIORAL of FA_1607 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U4 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1606 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1606;

architecture SYN_BEHAVIORAL of FA_1606 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1605 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1605;

architecture SYN_BEHAVIORAL of FA_1605 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1604 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1604;

architecture SYN_BEHAVIORAL of FA_1604 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1603 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1603;

architecture SYN_BEHAVIORAL of FA_1603 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n7, ZN => n5);
   U4 : INV_X1 port map( A => n5, ZN => Co);
   U5 : INV_X1 port map( A => A, ZN => n6);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1602 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1602;

architecture SYN_BEHAVIORAL of FA_1602 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n6, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n6, B2 => Ci, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1601 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1601;

architecture SYN_BEHAVIORAL of FA_1601 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1600 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1600;

architecture SYN_BEHAVIORAL of FA_1600 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1599 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1599;

architecture SYN_BEHAVIORAL of FA_1599 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1598 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1598;

architecture SYN_BEHAVIORAL of FA_1598 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1597 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1597;

architecture SYN_BEHAVIORAL of FA_1597 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1596 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1596;

architecture SYN_BEHAVIORAL of FA_1596 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1595 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1595;

architecture SYN_BEHAVIORAL of FA_1595 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1594 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1594;

architecture SYN_BEHAVIORAL of FA_1594 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1593 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1593;

architecture SYN_BEHAVIORAL of FA_1593 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1592 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1592;

architecture SYN_BEHAVIORAL of FA_1592 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1591 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1591;

architecture SYN_BEHAVIORAL of FA_1591 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1590 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1590;

architecture SYN_BEHAVIORAL of FA_1590 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1589 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1589;

architecture SYN_BEHAVIORAL of FA_1589 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1588 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1588;

architecture SYN_BEHAVIORAL of FA_1588 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1587 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1587;

architecture SYN_BEHAVIORAL of FA_1587 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1586 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1586;

architecture SYN_BEHAVIORAL of FA_1586 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1585 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1585;

architecture SYN_BEHAVIORAL of FA_1585 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n6, B2 => Ci, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1584 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1584;

architecture SYN_BEHAVIORAL of FA_1584 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n5, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1583 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1583;

architecture SYN_BEHAVIORAL of FA_1583 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U4 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1582 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1582;

architecture SYN_BEHAVIORAL of FA_1582 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1581 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1581;

architecture SYN_BEHAVIORAL of FA_1581 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1580 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1580;

architecture SYN_BEHAVIORAL of FA_1580 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1579 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1579;

architecture SYN_BEHAVIORAL of FA_1579 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1578 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1578;

architecture SYN_BEHAVIORAL of FA_1578 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1577 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1577;

architecture SYN_BEHAVIORAL of FA_1577 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1576 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1576;

architecture SYN_BEHAVIORAL of FA_1576 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1575 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1575;

architecture SYN_BEHAVIORAL of FA_1575 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n5);
   U5 : INV_X1 port map( A => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1574 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1574;

architecture SYN_BEHAVIORAL of FA_1574 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1573 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1573;

architecture SYN_BEHAVIORAL of FA_1573 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : OAI22_X1 port map( A1 => n5, A2 => n9, B1 => n7, B2 => n6, ZN => Co);
   U4 : INV_X1 port map( A => n4, ZN => n5);
   U5 : INV_X1 port map( A => n8, ZN => n6);
   U6 : INV_X1 port map( A => Ci, ZN => n7);
   U7 : INV_X1 port map( A => A, ZN => n9);
   U8 : XNOR2_X1 port map( A => B, B => n9, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1572 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1572;

architecture SYN_BEHAVIORAL of FA_1572 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1571 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1571;

architecture SYN_BEHAVIORAL of FA_1571 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1570 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1570;

architecture SYN_BEHAVIORAL of FA_1570 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1569 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1569;

architecture SYN_BEHAVIORAL of FA_1569 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : INV_X1 port map( A => n2, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1568 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1568;

architecture SYN_BEHAVIORAL of FA_1568 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n8, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : INV_X1 port map( A => n7, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n8);
   U7 : XNOR2_X1 port map( A => B, B => n8, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1567 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1567;

architecture SYN_BEHAVIORAL of FA_1567 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1566 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1566;

architecture SYN_BEHAVIORAL of FA_1566 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1565 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1565;

architecture SYN_BEHAVIORAL of FA_1565 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1564 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1564;

architecture SYN_BEHAVIORAL of FA_1564 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U2 : INV_X1 port map( A => n4, ZN => Co);
   U4 : INV_X1 port map( A => A, ZN => n6);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1563 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1563;

architecture SYN_BEHAVIORAL of FA_1563 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : INV_X1 port map( A => n2, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1562 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1562;

architecture SYN_BEHAVIORAL of FA_1562 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1561 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1561;

architecture SYN_BEHAVIORAL of FA_1561 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n8, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : INV_X1 port map( A => n7, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n8);
   U7 : XNOR2_X1 port map( A => B, B => n8, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1560 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1560;

architecture SYN_BEHAVIORAL of FA_1560 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n8, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : INV_X1 port map( A => n7, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n8);
   U7 : XNOR2_X1 port map( A => B, B => n8, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1559 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1559;

architecture SYN_BEHAVIORAL of FA_1559 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : INV_X1 port map( A => n2, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1558 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1558;

architecture SYN_BEHAVIORAL of FA_1558 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1557 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1557;

architecture SYN_BEHAVIORAL of FA_1557 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1556 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1556;

architecture SYN_BEHAVIORAL of FA_1556 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1555 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1555;

architecture SYN_BEHAVIORAL of FA_1555 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1554 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1554;

architecture SYN_BEHAVIORAL of FA_1554 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n8, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : INV_X1 port map( A => n7, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n8);
   U7 : XNOR2_X1 port map( A => B, B => n8, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1553 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1553;

architecture SYN_BEHAVIORAL of FA_1553 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1552 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1552;

architecture SYN_BEHAVIORAL of FA_1552 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1551 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1551;

architecture SYN_BEHAVIORAL of FA_1551 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1550 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1550;

architecture SYN_BEHAVIORAL of FA_1550 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1549 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1549;

architecture SYN_BEHAVIORAL of FA_1549 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1548 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1548;

architecture SYN_BEHAVIORAL of FA_1548 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1547 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1547;

architecture SYN_BEHAVIORAL of FA_1547 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1546 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1546;

architecture SYN_BEHAVIORAL of FA_1546 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => n6, B => B, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1545 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1545;

architecture SYN_BEHAVIORAL of FA_1545 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n8, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : INV_X1 port map( A => n7, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n8);
   U7 : XNOR2_X1 port map( A => B, B => n8, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1544 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1544;

architecture SYN_BEHAVIORAL of FA_1544 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1543 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1543;

architecture SYN_BEHAVIORAL of FA_1543 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1542 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1542;

architecture SYN_BEHAVIORAL of FA_1542 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n8, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : INV_X1 port map( A => n7, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n8);
   U7 : XNOR2_X1 port map( A => B, B => n8, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1541 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1541;

architecture SYN_BEHAVIORAL of FA_1541 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n5, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1540 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1540;

architecture SYN_BEHAVIORAL of FA_1540 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n5);
   U5 : INV_X1 port map( A => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1539 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1539;

architecture SYN_BEHAVIORAL of FA_1539 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n5);
   U5 : INV_X1 port map( A => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1538 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1538;

architecture SYN_BEHAVIORAL of FA_1538 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n6, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n6, B2 => Ci, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1537 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1537;

architecture SYN_BEHAVIORAL of FA_1537 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1536 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1536;

architecture SYN_BEHAVIORAL of FA_1536 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1535 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1535;

architecture SYN_BEHAVIORAL of FA_1535 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1534 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1534;

architecture SYN_BEHAVIORAL of FA_1534 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1533 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1533;

architecture SYN_BEHAVIORAL of FA_1533 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1532 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1532;

architecture SYN_BEHAVIORAL of FA_1532 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1531 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1531;

architecture SYN_BEHAVIORAL of FA_1531 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1530 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1530;

architecture SYN_BEHAVIORAL of FA_1530 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1529 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1529;

architecture SYN_BEHAVIORAL of FA_1529 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1528 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1528;

architecture SYN_BEHAVIORAL of FA_1528 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1527 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1527;

architecture SYN_BEHAVIORAL of FA_1527 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1526 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1526;

architecture SYN_BEHAVIORAL of FA_1526 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1525 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1525;

architecture SYN_BEHAVIORAL of FA_1525 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1524 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1524;

architecture SYN_BEHAVIORAL of FA_1524 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1523 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1523;

architecture SYN_BEHAVIORAL of FA_1523 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1522 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1522;

architecture SYN_BEHAVIORAL of FA_1522 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1521 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1521;

architecture SYN_BEHAVIORAL of FA_1521 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1520 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1520;

architecture SYN_BEHAVIORAL of FA_1520 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1519 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1519;

architecture SYN_BEHAVIORAL of FA_1519 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => n6, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n6, B2 => Ci, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1518 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1518;

architecture SYN_BEHAVIORAL of FA_1518 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : CLKBUF_X1 port map( A => Ci, Z => n4);
   U4 : CLKBUF_X1 port map( A => n8, Z => n5);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n8);
   U6 : CLKBUF_X1 port map( A => B, Z => n7);
   U7 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n8, ZN => n9);
   U8 : INV_X1 port map( A => n9, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1517 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1517;

architecture SYN_BEHAVIORAL of FA_1517 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1516 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1516;

architecture SYN_BEHAVIORAL of FA_1516 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U4 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1515 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1515;

architecture SYN_BEHAVIORAL of FA_1515 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1514 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1514;

architecture SYN_BEHAVIORAL of FA_1514 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1513 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1513;

architecture SYN_BEHAVIORAL of FA_1513 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : INV_X1 port map( A => n2, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1512 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1512;

architecture SYN_BEHAVIORAL of FA_1512 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1511 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1511;

architecture SYN_BEHAVIORAL of FA_1511 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1510 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1510;

architecture SYN_BEHAVIORAL of FA_1510 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1509 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1509;

architecture SYN_BEHAVIORAL of FA_1509 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n8, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => n7, ZN => n5);
   U5 : INV_X1 port map( A => Ci, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n8);
   U7 : XNOR2_X1 port map( A => B, B => n8, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1508 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1508;

architecture SYN_BEHAVIORAL of FA_1508 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1507 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1507;

architecture SYN_BEHAVIORAL of FA_1507 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1506 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1506;

architecture SYN_BEHAVIORAL of FA_1506 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1505 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1505;

architecture SYN_BEHAVIORAL of FA_1505 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1504 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1504;

architecture SYN_BEHAVIORAL of FA_1504 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1503 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1503;

architecture SYN_BEHAVIORAL of FA_1503 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1502 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1502;

architecture SYN_BEHAVIORAL of FA_1502 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1501 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1501;

architecture SYN_BEHAVIORAL of FA_1501 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1500 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1500;

architecture SYN_BEHAVIORAL of FA_1500 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n7, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : INV_X1 port map( A => n8, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n7);
   U7 : XNOR2_X1 port map( A => B, B => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1499 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1499;

architecture SYN_BEHAVIORAL of FA_1499 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U5 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1498 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1498;

architecture SYN_BEHAVIORAL of FA_1498 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1497 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1497;

architecture SYN_BEHAVIORAL of FA_1497 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n7, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : INV_X1 port map( A => n8, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n7);
   U7 : XNOR2_X1 port map( A => B, B => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1496 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1496;

architecture SYN_BEHAVIORAL of FA_1496 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1495 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1495;

architecture SYN_BEHAVIORAL of FA_1495 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U5 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1494 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1494;

architecture SYN_BEHAVIORAL of FA_1494 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n4);
   U2 : INV_X1 port map( A => n4, ZN => Co);
   U4 : INV_X1 port map( A => A, ZN => n5);
   U5 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1493 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1493;

architecture SYN_BEHAVIORAL of FA_1493 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n4);
   U2 : INV_X1 port map( A => n4, ZN => Co);
   U4 : INV_X1 port map( A => A, ZN => n5);
   U5 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1492 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1492;

architecture SYN_BEHAVIORAL of FA_1492 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n7, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : INV_X1 port map( A => n8, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n7);
   U7 : XNOR2_X1 port map( A => B, B => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1491 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1491;

architecture SYN_BEHAVIORAL of FA_1491 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U4 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1490 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1490;

architecture SYN_BEHAVIORAL of FA_1490 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : XNOR2_X1 port map( A => Ci, B => n7, ZN => n4);
   U3 : INV_X1 port map( A => n4, ZN => S);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n7);
   U6 : INV_X1 port map( A => n8, ZN => Co);
   U7 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1489 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1489;

architecture SYN_BEHAVIORAL of FA_1489 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1488 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1488;

architecture SYN_BEHAVIORAL of FA_1488 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1487 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1487;

architecture SYN_BEHAVIORAL of FA_1487 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1486 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1486;

architecture SYN_BEHAVIORAL of FA_1486 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1485 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1485;

architecture SYN_BEHAVIORAL of FA_1485 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U4 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1484 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1484;

architecture SYN_BEHAVIORAL of FA_1484 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n7, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : INV_X1 port map( A => n8, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n7);
   U7 : XNOR2_X1 port map( A => B, B => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1483 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1483;

architecture SYN_BEHAVIORAL of FA_1483 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n4);
   U2 : INV_X1 port map( A => n4, ZN => Co);
   U4 : INV_X1 port map( A => A, ZN => n5);
   U5 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1482 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1482;

architecture SYN_BEHAVIORAL of FA_1482 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n7, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : INV_X1 port map( A => n8, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n7);
   U7 : XNOR2_X1 port map( A => B, B => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1481 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1481;

architecture SYN_BEHAVIORAL of FA_1481 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1480 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1480;

architecture SYN_BEHAVIORAL of FA_1480 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1479 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1479;

architecture SYN_BEHAVIORAL of FA_1479 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1478 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1478;

architecture SYN_BEHAVIORAL of FA_1478 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1477 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1477;

architecture SYN_BEHAVIORAL of FA_1477 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1476 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1476;

architecture SYN_BEHAVIORAL of FA_1476 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1475 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1475;

architecture SYN_BEHAVIORAL of FA_1475 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1474 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1474;

architecture SYN_BEHAVIORAL of FA_1474 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n2);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U5 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1473 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1473;

architecture SYN_BEHAVIORAL of FA_1473 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1472 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1472;

architecture SYN_BEHAVIORAL of FA_1472 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1471 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1471;

architecture SYN_BEHAVIORAL of FA_1471 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1470 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1470;

architecture SYN_BEHAVIORAL of FA_1470 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1469 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1469;

architecture SYN_BEHAVIORAL of FA_1469 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1468 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1468;

architecture SYN_BEHAVIORAL of FA_1468 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1467 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1467;

architecture SYN_BEHAVIORAL of FA_1467 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1466 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1466;

architecture SYN_BEHAVIORAL of FA_1466 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1465 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1465;

architecture SYN_BEHAVIORAL of FA_1465 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1464 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1464;

architecture SYN_BEHAVIORAL of FA_1464 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1463 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1463;

architecture SYN_BEHAVIORAL of FA_1463 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1462 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1462;

architecture SYN_BEHAVIORAL of FA_1462 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1461 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1461;

architecture SYN_BEHAVIORAL of FA_1461 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1460 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1460;

architecture SYN_BEHAVIORAL of FA_1460 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1459 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1459;

architecture SYN_BEHAVIORAL of FA_1459 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1458 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1458;

architecture SYN_BEHAVIORAL of FA_1458 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1457 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1457;

architecture SYN_BEHAVIORAL of FA_1457 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1456 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1456;

architecture SYN_BEHAVIORAL of FA_1456 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1455 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1455;

architecture SYN_BEHAVIORAL of FA_1455 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1454 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1454;

architecture SYN_BEHAVIORAL of FA_1454 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1453 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1453;

architecture SYN_BEHAVIORAL of FA_1453 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1452 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1452;

architecture SYN_BEHAVIORAL of FA_1452 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1451 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1451;

architecture SYN_BEHAVIORAL of FA_1451 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n5, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1450 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1450;

architecture SYN_BEHAVIORAL of FA_1450 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1449 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1449;

architecture SYN_BEHAVIORAL of FA_1449 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n2);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U5 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1448 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1448;

architecture SYN_BEHAVIORAL of FA_1448 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1447 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1447;

architecture SYN_BEHAVIORAL of FA_1447 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1446 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1446;

architecture SYN_BEHAVIORAL of FA_1446 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1445 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1445;

architecture SYN_BEHAVIORAL of FA_1445 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U5 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1444 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1444;

architecture SYN_BEHAVIORAL of FA_1444 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1443 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1443;

architecture SYN_BEHAVIORAL of FA_1443 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1442 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1442;

architecture SYN_BEHAVIORAL of FA_1442 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1441 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1441;

architecture SYN_BEHAVIORAL of FA_1441 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : INV_X1 port map( A => n2, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1440 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1440;

architecture SYN_BEHAVIORAL of FA_1440 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n8, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : INV_X1 port map( A => n7, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n8);
   U7 : XNOR2_X1 port map( A => B, B => n8, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1439 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1439;

architecture SYN_BEHAVIORAL of FA_1439 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n5, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1438 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1438;

architecture SYN_BEHAVIORAL of FA_1438 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1437 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1437;

architecture SYN_BEHAVIORAL of FA_1437 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n7, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : INV_X1 port map( A => n8, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n7);
   U7 : XNOR2_X1 port map( A => B, B => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1436 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1436;

architecture SYN_BEHAVIORAL of FA_1436 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n7, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : INV_X1 port map( A => n8, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n7);
   U7 : XNOR2_X1 port map( A => B, B => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1435 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1435;

architecture SYN_BEHAVIORAL of FA_1435 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n5, ZN => n2);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1434 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1434;

architecture SYN_BEHAVIORAL of FA_1434 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => n5, B => B, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1433 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1433;

architecture SYN_BEHAVIORAL of FA_1433 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n4);
   U2 : INV_X1 port map( A => n4, ZN => Co);
   U4 : INV_X1 port map( A => A, ZN => n5);
   U5 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1432 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1432;

architecture SYN_BEHAVIORAL of FA_1432 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1431 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1431;

architecture SYN_BEHAVIORAL of FA_1431 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : XNOR2_X1 port map( A => n5, B => B, ZN => n4);
   U5 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1430 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1430;

architecture SYN_BEHAVIORAL of FA_1430 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1429 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1429;

architecture SYN_BEHAVIORAL of FA_1429 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n4);
   U2 : INV_X1 port map( A => n4, ZN => Co);
   U4 : INV_X1 port map( A => A, ZN => n5);
   U5 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1428 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1428;

architecture SYN_BEHAVIORAL of FA_1428 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1427 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1427;

architecture SYN_BEHAVIORAL of FA_1427 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1426 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1426;

architecture SYN_BEHAVIORAL of FA_1426 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n7, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : INV_X1 port map( A => n8, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n7);
   U7 : XNOR2_X1 port map( A => B, B => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1425 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1425;

architecture SYN_BEHAVIORAL of FA_1425 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1424 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1424;

architecture SYN_BEHAVIORAL of FA_1424 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1423 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1423;

architecture SYN_BEHAVIORAL of FA_1423 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1422 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1422;

architecture SYN_BEHAVIORAL of FA_1422 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1421 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1421;

architecture SYN_BEHAVIORAL of FA_1421 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U4 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1420 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1420;

architecture SYN_BEHAVIORAL of FA_1420 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n7, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : INV_X1 port map( A => n8, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n7);
   U7 : XNOR2_X1 port map( A => B, B => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1419 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1419;

architecture SYN_BEHAVIORAL of FA_1419 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n7, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : INV_X1 port map( A => n8, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n7);
   U7 : XNOR2_X1 port map( A => B, B => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1418 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1418;

architecture SYN_BEHAVIORAL of FA_1418 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1417 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1417;

architecture SYN_BEHAVIORAL of FA_1417 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1416 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1416;

architecture SYN_BEHAVIORAL of FA_1416 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1415 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1415;

architecture SYN_BEHAVIORAL of FA_1415 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1414 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1414;

architecture SYN_BEHAVIORAL of FA_1414 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1413 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1413;

architecture SYN_BEHAVIORAL of FA_1413 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1412 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1412;

architecture SYN_BEHAVIORAL of FA_1412 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1411 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1411;

architecture SYN_BEHAVIORAL of FA_1411 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n9, n10 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n8);
   U2 : NAND2_X1 port map( A1 => Ci, A2 => n5, ZN => n6);
   U3 : NAND2_X1 port map( A1 => n4, A2 => n9, ZN => n7);
   U4 : NAND2_X1 port map( A1 => n7, A2 => n6, ZN => S);
   U5 : INV_X1 port map( A => Ci, ZN => n4);
   U6 : INV_X1 port map( A => n9, ZN => n5);
   U7 : XNOR2_X1 port map( A => B, B => n8, ZN => n9);
   U8 : INV_X1 port map( A => n10, ZN => Co);
   U9 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n9, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1410 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1410;

architecture SYN_BEHAVIORAL of FA_1410 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n2);
   U5 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1409 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1409;

architecture SYN_BEHAVIORAL of FA_1409 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U1 : MUX2_X1 port map( A => n7, B => n5, S => Ci, Z => S);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U3 : XOR2_X1 port map( A => B, B => n6, Z => n5);
   U4 : INV_X1 port map( A => A, ZN => n6);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n7);
   U6 : INV_X1 port map( A => n8, ZN => Co);
   U7 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n7, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1408 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1408;

architecture SYN_BEHAVIORAL of FA_1408 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1407 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1407;

architecture SYN_BEHAVIORAL of FA_1407 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1406 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1406;

architecture SYN_BEHAVIORAL of FA_1406 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1405 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1405;

architecture SYN_BEHAVIORAL of FA_1405 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1404 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1404;

architecture SYN_BEHAVIORAL of FA_1404 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1403 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1403;

architecture SYN_BEHAVIORAL of FA_1403 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1402 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1402;

architecture SYN_BEHAVIORAL of FA_1402 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1401 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1401;

architecture SYN_BEHAVIORAL of FA_1401 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1400 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1400;

architecture SYN_BEHAVIORAL of FA_1400 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1399 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1399;

architecture SYN_BEHAVIORAL of FA_1399 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1398 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1398;

architecture SYN_BEHAVIORAL of FA_1398 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1397 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1397;

architecture SYN_BEHAVIORAL of FA_1397 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1396 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1396;

architecture SYN_BEHAVIORAL of FA_1396 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1395 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1395;

architecture SYN_BEHAVIORAL of FA_1395 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1394 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1394;

architecture SYN_BEHAVIORAL of FA_1394 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1393 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1393;

architecture SYN_BEHAVIORAL of FA_1393 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1392 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1392;

architecture SYN_BEHAVIORAL of FA_1392 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1391 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1391;

architecture SYN_BEHAVIORAL of FA_1391 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1390 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1390;

architecture SYN_BEHAVIORAL of FA_1390 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1389 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1389;

architecture SYN_BEHAVIORAL of FA_1389 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1388 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1388;

architecture SYN_BEHAVIORAL of FA_1388 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1387 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1387;

architecture SYN_BEHAVIORAL of FA_1387 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1386 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1386;

architecture SYN_BEHAVIORAL of FA_1386 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1385 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1385;

architecture SYN_BEHAVIORAL of FA_1385 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U5 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1384 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1384;

architecture SYN_BEHAVIORAL of FA_1384 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1383 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1383;

architecture SYN_BEHAVIORAL of FA_1383 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n5);
   U5 : INV_X1 port map( A => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1382 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1382;

architecture SYN_BEHAVIORAL of FA_1382 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1381 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1381;

architecture SYN_BEHAVIORAL of FA_1381 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U5 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1380 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1380;

architecture SYN_BEHAVIORAL of FA_1380 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1379 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1379;

architecture SYN_BEHAVIORAL of FA_1379 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1378 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1378;

architecture SYN_BEHAVIORAL of FA_1378 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1377 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1377;

architecture SYN_BEHAVIORAL of FA_1377 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : INV_X1 port map( A => n2, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1376 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1376;

architecture SYN_BEHAVIORAL of FA_1376 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : OAI22_X1 port map( A1 => n5, A2 => n9, B1 => n6, B2 => n7, ZN => Co);
   U4 : INV_X1 port map( A => n4, ZN => n5);
   U5 : INV_X1 port map( A => Ci, ZN => n6);
   U6 : INV_X1 port map( A => n8, ZN => n7);
   U7 : INV_X1 port map( A => A, ZN => n9);
   U8 : XNOR2_X1 port map( A => B, B => n9, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1375 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1375;

architecture SYN_BEHAVIORAL of FA_1375 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1374 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1374;

architecture SYN_BEHAVIORAL of FA_1374 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1373 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1373;

architecture SYN_BEHAVIORAL of FA_1373 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : OAI22_X1 port map( A1 => n8, A2 => n4, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : INV_X1 port map( A => n7, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n8);
   U7 : XNOR2_X1 port map( A => B, B => n8, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1372 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1372;

architecture SYN_BEHAVIORAL of FA_1372 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1371 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1371;

architecture SYN_BEHAVIORAL of FA_1371 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : INV_X1 port map( A => n2, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1370 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1370;

architecture SYN_BEHAVIORAL of FA_1370 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1369 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1369;

architecture SYN_BEHAVIORAL of FA_1369 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n8, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : INV_X1 port map( A => n7, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n8);
   U7 : XNOR2_X1 port map( A => B, B => n8, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1368 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1368;

architecture SYN_BEHAVIORAL of FA_1368 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1367 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1367;

architecture SYN_BEHAVIORAL of FA_1367 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : INV_X1 port map( A => n2, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1366 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1366;

architecture SYN_BEHAVIORAL of FA_1366 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1365 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1365;

architecture SYN_BEHAVIORAL of FA_1365 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1364 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1364;

architecture SYN_BEHAVIORAL of FA_1364 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1363 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1363;

architecture SYN_BEHAVIORAL of FA_1363 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1362 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1362;

architecture SYN_BEHAVIORAL of FA_1362 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n8, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : INV_X1 port map( A => n7, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n8);
   U7 : XNOR2_X1 port map( A => B, B => n8, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1361 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1361;

architecture SYN_BEHAVIORAL of FA_1361 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1360 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1360;

architecture SYN_BEHAVIORAL of FA_1360 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1359 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1359;

architecture SYN_BEHAVIORAL of FA_1359 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1358 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1358;

architecture SYN_BEHAVIORAL of FA_1358 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n8, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : INV_X1 port map( A => n7, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n8);
   U7 : XNOR2_X1 port map( A => B, B => n8, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1357 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1357;

architecture SYN_BEHAVIORAL of FA_1357 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1356 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1356;

architecture SYN_BEHAVIORAL of FA_1356 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n8, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : INV_X1 port map( A => n7, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n8);
   U7 : XNOR2_X1 port map( A => B, B => n8, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1355 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1355;

architecture SYN_BEHAVIORAL of FA_1355 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n5, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1354 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1354;

architecture SYN_BEHAVIORAL of FA_1354 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1353 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1353;

architecture SYN_BEHAVIORAL of FA_1353 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1352 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1352;

architecture SYN_BEHAVIORAL of FA_1352 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U2 : INV_X1 port map( A => n4, ZN => Co);
   U4 : INV_X1 port map( A => A, ZN => n6);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1351 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1351;

architecture SYN_BEHAVIORAL of FA_1351 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1350 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1350;

architecture SYN_BEHAVIORAL of FA_1350 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1349 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1349;

architecture SYN_BEHAVIORAL of FA_1349 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1348 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1348;

architecture SYN_BEHAVIORAL of FA_1348 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1347 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1347;

architecture SYN_BEHAVIORAL of FA_1347 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n6, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n5);
   U5 : INV_X1 port map( A => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1346 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1346;

architecture SYN_BEHAVIORAL of FA_1346 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U3 : MUX2_X1 port map( A => n5, B => n7, S => Ci, Z => S);
   U4 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n5, B2 => Ci, ZN => n2);
   U6 : INV_X1 port map( A => A, ZN => n6);
   U7 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1345 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1345;

architecture SYN_BEHAVIORAL of FA_1345 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => n7, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n7);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : INV_X1 port map( A => n8, ZN => Co);
   U7 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => n4, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1344 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1344;

architecture SYN_BEHAVIORAL of FA_1344 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1343 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1343;

architecture SYN_BEHAVIORAL of FA_1343 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1342 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1342;

architecture SYN_BEHAVIORAL of FA_1342 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1341 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1341;

architecture SYN_BEHAVIORAL of FA_1341 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1340 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1340;

architecture SYN_BEHAVIORAL of FA_1340 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1339 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1339;

architecture SYN_BEHAVIORAL of FA_1339 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1338 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1338;

architecture SYN_BEHAVIORAL of FA_1338 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1337 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1337;

architecture SYN_BEHAVIORAL of FA_1337 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1336 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1336;

architecture SYN_BEHAVIORAL of FA_1336 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1335 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1335;

architecture SYN_BEHAVIORAL of FA_1335 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1334 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1334;

architecture SYN_BEHAVIORAL of FA_1334 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1333 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1333;

architecture SYN_BEHAVIORAL of FA_1333 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1332 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1332;

architecture SYN_BEHAVIORAL of FA_1332 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1331 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1331;

architecture SYN_BEHAVIORAL of FA_1331 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1330 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1330;

architecture SYN_BEHAVIORAL of FA_1330 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1329 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1329;

architecture SYN_BEHAVIORAL of FA_1329 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1328 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1328;

architecture SYN_BEHAVIORAL of FA_1328 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1327 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1327;

architecture SYN_BEHAVIORAL of FA_1327 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1326 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1326;

architecture SYN_BEHAVIORAL of FA_1326 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1325 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1325;

architecture SYN_BEHAVIORAL of FA_1325 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1324 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1324;

architecture SYN_BEHAVIORAL of FA_1324 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1323 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1323;

architecture SYN_BEHAVIORAL of FA_1323 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1322 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1322;

architecture SYN_BEHAVIORAL of FA_1322 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1321 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1321;

architecture SYN_BEHAVIORAL of FA_1321 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1320 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1320;

architecture SYN_BEHAVIORAL of FA_1320 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1319 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1319;

architecture SYN_BEHAVIORAL of FA_1319 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n5, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n5);
   U4 : AOI22_X1 port map( A1 => A, A2 => B, B1 => n5, B2 => Ci, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1318 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1318;

architecture SYN_BEHAVIORAL of FA_1318 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1317 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1317;

architecture SYN_BEHAVIORAL of FA_1317 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1316 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1316;

architecture SYN_BEHAVIORAL of FA_1316 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1315 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1315;

architecture SYN_BEHAVIORAL of FA_1315 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1314 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1314;

architecture SYN_BEHAVIORAL of FA_1314 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1313 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1313;

architecture SYN_BEHAVIORAL of FA_1313 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n4);
   U2 : INV_X1 port map( A => n4, ZN => Co);
   U4 : INV_X1 port map( A => A, ZN => n5);
   U5 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1312 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1312;

architecture SYN_BEHAVIORAL of FA_1312 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n5, B => Ci, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n5, ZN => n2);
   U5 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1311 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1311;

architecture SYN_BEHAVIORAL of FA_1311 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1310 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1310;

architecture SYN_BEHAVIORAL of FA_1310 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1309 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1309;

architecture SYN_BEHAVIORAL of FA_1309 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n8, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : INV_X1 port map( A => n7, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n8);
   U7 : XNOR2_X1 port map( A => B, B => n8, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1308 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1308;

architecture SYN_BEHAVIORAL of FA_1308 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n8, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : INV_X1 port map( A => n7, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n8);
   U7 : XNOR2_X1 port map( A => B, B => n8, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1307 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1307;

architecture SYN_BEHAVIORAL of FA_1307 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U5 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1306 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1306;

architecture SYN_BEHAVIORAL of FA_1306 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U4 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1305 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1305;

architecture SYN_BEHAVIORAL of FA_1305 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U4 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1304 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1304;

architecture SYN_BEHAVIORAL of FA_1304 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U4 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1303 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1303;

architecture SYN_BEHAVIORAL of FA_1303 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U5 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1302 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1302;

architecture SYN_BEHAVIORAL of FA_1302 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n7, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : INV_X1 port map( A => n8, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n7);
   U7 : XNOR2_X1 port map( A => n7, B => B, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1301 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1301;

architecture SYN_BEHAVIORAL of FA_1301 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n5, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U4 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1300 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1300;

architecture SYN_BEHAVIORAL of FA_1300 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U4 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1299 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1299;

architecture SYN_BEHAVIORAL of FA_1299 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => n5, B => B, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1298 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1298;

architecture SYN_BEHAVIORAL of FA_1298 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U4 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1297 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1297;

architecture SYN_BEHAVIORAL of FA_1297 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1296 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1296;

architecture SYN_BEHAVIORAL of FA_1296 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1295 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1295;

architecture SYN_BEHAVIORAL of FA_1295 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n7, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : INV_X1 port map( A => n8, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n7);
   U7 : XNOR2_X1 port map( A => B, B => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1294 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1294;

architecture SYN_BEHAVIORAL of FA_1294 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1293 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1293;

architecture SYN_BEHAVIORAL of FA_1293 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U4 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1292 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1292;

architecture SYN_BEHAVIORAL of FA_1292 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n9, Z => S);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : OAI22_X1 port map( A1 => n5, A2 => n8, B1 => n6, B2 => n7, ZN => Co);
   U4 : INV_X1 port map( A => n4, ZN => n5);
   U5 : INV_X1 port map( A => Ci, ZN => n6);
   U6 : INV_X1 port map( A => n9, ZN => n7);
   U7 : INV_X1 port map( A => A, ZN => n8);
   U8 : XNOR2_X1 port map( A => B, B => n8, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1291 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1291;

architecture SYN_BEHAVIORAL of FA_1291 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1290 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1290;

architecture SYN_BEHAVIORAL of FA_1290 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1289 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1289;

architecture SYN_BEHAVIORAL of FA_1289 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1288 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1288;

architecture SYN_BEHAVIORAL of FA_1288 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1287 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1287;

architecture SYN_BEHAVIORAL of FA_1287 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1286 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1286;

architecture SYN_BEHAVIORAL of FA_1286 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n7, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : INV_X1 port map( A => n8, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n7);
   U7 : XNOR2_X1 port map( A => B, B => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1285 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1285;

architecture SYN_BEHAVIORAL of FA_1285 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1284 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1284;

architecture SYN_BEHAVIORAL of FA_1284 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1283 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1283;

architecture SYN_BEHAVIORAL of FA_1283 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n6, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n6, B2 => Ci, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1282 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1282;

architecture SYN_BEHAVIORAL of FA_1282 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n2);
   U5 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1281 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1281;

architecture SYN_BEHAVIORAL of FA_1281 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : CLKBUF_X1 port map( A => n7, Z => n5);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n7);
   U6 : INV_X1 port map( A => n8, ZN => Co);
   U7 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n5, B2 => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1280 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1280;

architecture SYN_BEHAVIORAL of FA_1280 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1279 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1279;

architecture SYN_BEHAVIORAL of FA_1279 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1278 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1278;

architecture SYN_BEHAVIORAL of FA_1278 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1277 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1277;

architecture SYN_BEHAVIORAL of FA_1277 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1276 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1276;

architecture SYN_BEHAVIORAL of FA_1276 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1275 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1275;

architecture SYN_BEHAVIORAL of FA_1275 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1274 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1274;

architecture SYN_BEHAVIORAL of FA_1274 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1273 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1273;

architecture SYN_BEHAVIORAL of FA_1273 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1272 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1272;

architecture SYN_BEHAVIORAL of FA_1272 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1271 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1271;

architecture SYN_BEHAVIORAL of FA_1271 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1270 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1270;

architecture SYN_BEHAVIORAL of FA_1270 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1269 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1269;

architecture SYN_BEHAVIORAL of FA_1269 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1268 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1268;

architecture SYN_BEHAVIORAL of FA_1268 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1267 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1267;

architecture SYN_BEHAVIORAL of FA_1267 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1266 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1266;

architecture SYN_BEHAVIORAL of FA_1266 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1265 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1265;

architecture SYN_BEHAVIORAL of FA_1265 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1264 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1264;

architecture SYN_BEHAVIORAL of FA_1264 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1263 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1263;

architecture SYN_BEHAVIORAL of FA_1263 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1262 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1262;

architecture SYN_BEHAVIORAL of FA_1262 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1261 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1261;

architecture SYN_BEHAVIORAL of FA_1261 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1260 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1260;

architecture SYN_BEHAVIORAL of FA_1260 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1259 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1259;

architecture SYN_BEHAVIORAL of FA_1259 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1258 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1258;

architecture SYN_BEHAVIORAL of FA_1258 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1257 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1257;

architecture SYN_BEHAVIORAL of FA_1257 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1256 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1256;

architecture SYN_BEHAVIORAL of FA_1256 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1255 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1255;

architecture SYN_BEHAVIORAL of FA_1255 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n6, B2 => Ci, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1254 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1254;

architecture SYN_BEHAVIORAL of FA_1254 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1253 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1253;

architecture SYN_BEHAVIORAL of FA_1253 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n5, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1252 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1252;

architecture SYN_BEHAVIORAL of FA_1252 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n5, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1251 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1251;

architecture SYN_BEHAVIORAL of FA_1251 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1250 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1250;

architecture SYN_BEHAVIORAL of FA_1250 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1249 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1249;

architecture SYN_BEHAVIORAL of FA_1249 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U5 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1248 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1248;

architecture SYN_BEHAVIORAL of FA_1248 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1247 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1247;

architecture SYN_BEHAVIORAL of FA_1247 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1246 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1246;

architecture SYN_BEHAVIORAL of FA_1246 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => n6, B => B, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1245 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1245;

architecture SYN_BEHAVIORAL of FA_1245 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1244 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1244;

architecture SYN_BEHAVIORAL of FA_1244 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U2 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1243 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1243;

architecture SYN_BEHAVIORAL of FA_1243 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : INV_X1 port map( A => n2, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1242 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1242;

architecture SYN_BEHAVIORAL of FA_1242 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U2 : INV_X1 port map( A => n4, ZN => Co);
   U4 : INV_X1 port map( A => A, ZN => n6);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1241 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1241;

architecture SYN_BEHAVIORAL of FA_1241 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => Ci, A2 => n5, ZN => n6);
   U2 : NAND2_X1 port map( A1 => n4, A2 => n11, ZN => n7);
   U3 : NAND2_X1 port map( A1 => n6, A2 => n7, ZN => S);
   U4 : INV_X1 port map( A => Ci, ZN => n4);
   U5 : INV_X1 port map( A => n11, ZN => n5);
   U6 : OAI22_X1 port map( A1 => n8, A2 => n12, B1 => n9, B2 => n10, ZN => Co);
   U7 : INV_X1 port map( A => B, ZN => n8);
   U8 : INV_X1 port map( A => Ci, ZN => n9);
   U9 : INV_X1 port map( A => n11, ZN => n10);
   U10 : INV_X1 port map( A => A, ZN => n12);
   U11 : XNOR2_X1 port map( A => B, B => n12, ZN => n11);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1240 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1240;

architecture SYN_BEHAVIORAL of FA_1240 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1239 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1239;

architecture SYN_BEHAVIORAL of FA_1239 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U4 : INV_X1 port map( A => n2, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1238 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1238;

architecture SYN_BEHAVIORAL of FA_1238 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1237 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1237;

architecture SYN_BEHAVIORAL of FA_1237 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1236 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1236;

architecture SYN_BEHAVIORAL of FA_1236 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1235 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1235;

architecture SYN_BEHAVIORAL of FA_1235 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n8, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : INV_X1 port map( A => n7, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n8);
   U7 : XNOR2_X1 port map( A => B, B => n8, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1234 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1234;

architecture SYN_BEHAVIORAL of FA_1234 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n8, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : INV_X1 port map( A => n7, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n8);
   U7 : XNOR2_X1 port map( A => B, B => n8, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1233 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1233;

architecture SYN_BEHAVIORAL of FA_1233 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1232 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1232;

architecture SYN_BEHAVIORAL of FA_1232 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U2 : INV_X1 port map( A => n4, ZN => Co);
   U4 : INV_X1 port map( A => A, ZN => n6);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1231 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1231;

architecture SYN_BEHAVIORAL of FA_1231 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n8, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : INV_X1 port map( A => n7, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n8);
   U7 : XNOR2_X1 port map( A => B, B => n8, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1230 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1230;

architecture SYN_BEHAVIORAL of FA_1230 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1229 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1229;

architecture SYN_BEHAVIORAL of FA_1229 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1228 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1228;

architecture SYN_BEHAVIORAL of FA_1228 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n8, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : INV_X1 port map( A => n7, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n8);
   U7 : XNOR2_X1 port map( A => B, B => n8, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1227 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1227;

architecture SYN_BEHAVIORAL of FA_1227 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U4 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1226 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1226;

architecture SYN_BEHAVIORAL of FA_1226 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1225 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1225;

architecture SYN_BEHAVIORAL of FA_1225 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n6);
   U4 : CLKBUF_X1 port map( A => B, Z => n5);
   U5 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1224 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1224;

architecture SYN_BEHAVIORAL of FA_1224 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1223 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1223;

architecture SYN_BEHAVIORAL of FA_1223 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n7, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : INV_X1 port map( A => n8, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n7);
   U7 : XNOR2_X1 port map( A => B, B => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1222 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1222;

architecture SYN_BEHAVIORAL of FA_1222 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1221 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1221;

architecture SYN_BEHAVIORAL of FA_1221 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => Co);
   U6 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1220 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1220;

architecture SYN_BEHAVIORAL of FA_1220 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n7);
   U6 : INV_X1 port map( A => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1219 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1219;

architecture SYN_BEHAVIORAL of FA_1219 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1218 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1218;

architecture SYN_BEHAVIORAL of FA_1218 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n7, B => Ci, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n8, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => n7, ZN => n5);
   U5 : INV_X1 port map( A => Ci, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n8);
   U7 : XNOR2_X1 port map( A => B, B => n8, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1217 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1217;

architecture SYN_BEHAVIORAL of FA_1217 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : CLKBUF_X1 port map( A => n8, Z => n4);
   U4 : CLKBUF_X1 port map( A => Ci, Z => n5);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n8);
   U7 : INV_X1 port map( A => n9, ZN => Co);
   U8 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => n4, B2 => n5, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1216 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1216;

architecture SYN_BEHAVIORAL of FA_1216 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1215 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1215;

architecture SYN_BEHAVIORAL of FA_1215 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1214 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1214;

architecture SYN_BEHAVIORAL of FA_1214 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1213 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1213;

architecture SYN_BEHAVIORAL of FA_1213 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1212 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1212;

architecture SYN_BEHAVIORAL of FA_1212 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1211 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1211;

architecture SYN_BEHAVIORAL of FA_1211 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1210 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1210;

architecture SYN_BEHAVIORAL of FA_1210 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1209 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1209;

architecture SYN_BEHAVIORAL of FA_1209 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1208 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1208;

architecture SYN_BEHAVIORAL of FA_1208 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1207 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1207;

architecture SYN_BEHAVIORAL of FA_1207 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1206 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1206;

architecture SYN_BEHAVIORAL of FA_1206 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1205 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1205;

architecture SYN_BEHAVIORAL of FA_1205 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1204 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1204;

architecture SYN_BEHAVIORAL of FA_1204 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1203 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1203;

architecture SYN_BEHAVIORAL of FA_1203 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1202 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1202;

architecture SYN_BEHAVIORAL of FA_1202 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1201 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1201;

architecture SYN_BEHAVIORAL of FA_1201 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1200 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1200;

architecture SYN_BEHAVIORAL of FA_1200 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1199 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1199;

architecture SYN_BEHAVIORAL of FA_1199 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1198 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1198;

architecture SYN_BEHAVIORAL of FA_1198 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1197 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1197;

architecture SYN_BEHAVIORAL of FA_1197 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1196 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1196;

architecture SYN_BEHAVIORAL of FA_1196 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1195 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1195;

architecture SYN_BEHAVIORAL of FA_1195 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1194 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1194;

architecture SYN_BEHAVIORAL of FA_1194 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1193 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1193;

architecture SYN_BEHAVIORAL of FA_1193 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1192 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1192;

architecture SYN_BEHAVIORAL of FA_1192 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1191 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1191;

architecture SYN_BEHAVIORAL of FA_1191 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1190 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1190;

architecture SYN_BEHAVIORAL of FA_1190 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1189 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1189;

architecture SYN_BEHAVIORAL of FA_1189 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1188 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1188;

architecture SYN_BEHAVIORAL of FA_1188 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n5, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1187 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1187;

architecture SYN_BEHAVIORAL of FA_1187 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1186 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1186;

architecture SYN_BEHAVIORAL of FA_1186 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1185 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1185;

architecture SYN_BEHAVIORAL of FA_1185 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1184 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1184;

architecture SYN_BEHAVIORAL of FA_1184 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1183 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1183;

architecture SYN_BEHAVIORAL of FA_1183 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1182 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1182;

architecture SYN_BEHAVIORAL of FA_1182 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1181 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1181;

architecture SYN_BEHAVIORAL of FA_1181 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1180 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1180;

architecture SYN_BEHAVIORAL of FA_1180 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1179 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1179;

architecture SYN_BEHAVIORAL of FA_1179 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1178 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1178;

architecture SYN_BEHAVIORAL of FA_1178 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1177 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1177;

architecture SYN_BEHAVIORAL of FA_1177 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U2 : INV_X1 port map( A => n5, ZN => Co);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1176 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1176;

architecture SYN_BEHAVIORAL of FA_1176 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1175 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1175;

architecture SYN_BEHAVIORAL of FA_1175 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U2 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1174 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1174;

architecture SYN_BEHAVIORAL of FA_1174 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n7, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : INV_X1 port map( A => n8, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n7);
   U7 : XNOR2_X1 port map( A => B, B => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1173 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1173;

architecture SYN_BEHAVIORAL of FA_1173 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1172 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1172;

architecture SYN_BEHAVIORAL of FA_1172 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n4);
   U2 : INV_X1 port map( A => n4, ZN => Co);
   U4 : INV_X1 port map( A => A, ZN => n5);
   U5 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1171 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1171;

architecture SYN_BEHAVIORAL of FA_1171 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n6, Z => S);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n6, ZN => n4);
   U2 : INV_X1 port map( A => n4, ZN => Co);
   U4 : INV_X1 port map( A => A, ZN => n5);
   U5 : XNOR2_X1 port map( A => B, B => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1170 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1170;

architecture SYN_BEHAVIORAL of FA_1170 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n7, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : INV_X1 port map( A => n8, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n7);
   U7 : XNOR2_X1 port map( A => B, B => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1169 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1169;

architecture SYN_BEHAVIORAL of FA_1169 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1168 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1168;

architecture SYN_BEHAVIORAL of FA_1168 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1167 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1167;

architecture SYN_BEHAVIORAL of FA_1167 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n5, B => n8, ZN => S);
   U2 : OAI22_X1 port map( A1 => n4, A2 => n7, B1 => n5, B2 => n6, ZN => Co);
   U3 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : INV_X1 port map( A => n8, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n7);
   U7 : XNOR2_X1 port map( A => B, B => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1166 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1166;

architecture SYN_BEHAVIORAL of FA_1166 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1165 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1165;

architecture SYN_BEHAVIORAL of FA_1165 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n7, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : INV_X1 port map( A => n8, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n7);
   U7 : XNOR2_X1 port map( A => n7, B => B, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1164 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1164;

architecture SYN_BEHAVIORAL of FA_1164 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U2 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1163 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1163;

architecture SYN_BEHAVIORAL of FA_1163 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1162 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1162;

architecture SYN_BEHAVIORAL of FA_1162 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1161 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1161;

architecture SYN_BEHAVIORAL of FA_1161 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n8, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : INV_X1 port map( A => n7, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n8);
   U7 : XNOR2_X1 port map( A => B, B => n8, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1160 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1160;

architecture SYN_BEHAVIORAL of FA_1160 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U2 : INV_X1 port map( A => n4, ZN => Co);
   U4 : INV_X1 port map( A => A, ZN => n6);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1159 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1159;

architecture SYN_BEHAVIORAL of FA_1159 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n8, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : INV_X1 port map( A => n7, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n8);
   U7 : XNOR2_X1 port map( A => B, B => n8, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1158 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1158;

architecture SYN_BEHAVIORAL of FA_1158 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U2 : INV_X1 port map( A => n4, ZN => Co);
   U4 : INV_X1 port map( A => A, ZN => n6);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1157 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1157;

architecture SYN_BEHAVIORAL of FA_1157 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n6, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n5);
   U5 : INV_X1 port map( A => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1156 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1156;

architecture SYN_BEHAVIORAL of FA_1156 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n8, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : INV_X1 port map( A => n7, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n8);
   U7 : XNOR2_X1 port map( A => B, B => n8, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1155 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1155;

architecture SYN_BEHAVIORAL of FA_1155 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n5, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1154 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1154;

architecture SYN_BEHAVIORAL of FA_1154 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => Ci, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n2);
   U5 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1153 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1153;

architecture SYN_BEHAVIORAL of FA_1153 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n6, n7, n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => Ci, ZN => n7);
   U2 : OR2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U3 : AND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : XNOR2_X1 port map( A => Ci, B => n8, ZN => S);
   U5 : NOR2_X1 port map( A1 => n8, A2 => n7, ZN => n6);
   U6 : XNOR2_X1 port map( A => B, B => A, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1152 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1152;

architecture SYN_BEHAVIORAL of FA_1152 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1151 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1151;

architecture SYN_BEHAVIORAL of FA_1151 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1150 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1150;

architecture SYN_BEHAVIORAL of FA_1150 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1149 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1149;

architecture SYN_BEHAVIORAL of FA_1149 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1148 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1148;

architecture SYN_BEHAVIORAL of FA_1148 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1147 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1147;

architecture SYN_BEHAVIORAL of FA_1147 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1146 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1146;

architecture SYN_BEHAVIORAL of FA_1146 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1145 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1145;

architecture SYN_BEHAVIORAL of FA_1145 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1144 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1144;

architecture SYN_BEHAVIORAL of FA_1144 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1143 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1143;

architecture SYN_BEHAVIORAL of FA_1143 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1142 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1142;

architecture SYN_BEHAVIORAL of FA_1142 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1141 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1141;

architecture SYN_BEHAVIORAL of FA_1141 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1140 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1140;

architecture SYN_BEHAVIORAL of FA_1140 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1139 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1139;

architecture SYN_BEHAVIORAL of FA_1139 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1138 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1138;

architecture SYN_BEHAVIORAL of FA_1138 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1137 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1137;

architecture SYN_BEHAVIORAL of FA_1137 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1136 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1136;

architecture SYN_BEHAVIORAL of FA_1136 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1135 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1135;

architecture SYN_BEHAVIORAL of FA_1135 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1134 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1134;

architecture SYN_BEHAVIORAL of FA_1134 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1133 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1133;

architecture SYN_BEHAVIORAL of FA_1133 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1132 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1132;

architecture SYN_BEHAVIORAL of FA_1132 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1131 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1131;

architecture SYN_BEHAVIORAL of FA_1131 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1130 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1130;

architecture SYN_BEHAVIORAL of FA_1130 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1129 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1129;

architecture SYN_BEHAVIORAL of FA_1129 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1128 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1128;

architecture SYN_BEHAVIORAL of FA_1128 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1127 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1127;

architecture SYN_BEHAVIORAL of FA_1127 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1126 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1126;

architecture SYN_BEHAVIORAL of FA_1126 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1125 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1125;

architecture SYN_BEHAVIORAL of FA_1125 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1124 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1124;

architecture SYN_BEHAVIORAL of FA_1124 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1123 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1123;

architecture SYN_BEHAVIORAL of FA_1123 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1122 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1122;

architecture SYN_BEHAVIORAL of FA_1122 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => Ci, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1121 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1121;

architecture SYN_BEHAVIORAL of FA_1121 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1120 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1120;

architecture SYN_BEHAVIORAL of FA_1120 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1119 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1119;

architecture SYN_BEHAVIORAL of FA_1119 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1118 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1118;

architecture SYN_BEHAVIORAL of FA_1118 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1117 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1117;

architecture SYN_BEHAVIORAL of FA_1117 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1116 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1116;

architecture SYN_BEHAVIORAL of FA_1116 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1115 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1115;

architecture SYN_BEHAVIORAL of FA_1115 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1114 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1114;

architecture SYN_BEHAVIORAL of FA_1114 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n8);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n5, B1 => n6, B2 => n7, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U5 : INV_X1 port map( A => A, ZN => n5);
   U6 : INV_X1 port map( A => n8, ZN => n6);
   U7 : INV_X1 port map( A => Ci, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1113 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1113;

architecture SYN_BEHAVIORAL of FA_1113 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1112 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1112;

architecture SYN_BEHAVIORAL of FA_1112 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1111 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1111;

architecture SYN_BEHAVIORAL of FA_1111 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U2 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1110 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1110;

architecture SYN_BEHAVIORAL of FA_1110 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n9 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => n9);
   U3 : XNOR2_X1 port map( A => Ci, B => n8, ZN => S);
   U4 : OAI22_X1 port map( A1 => n5, A2 => n6, B1 => n7, B2 => n8, ZN => Co);
   U5 : INV_X1 port map( A => B, ZN => n5);
   U6 : INV_X1 port map( A => A, ZN => n6);
   U7 : INV_X1 port map( A => Ci, ZN => n7);
   U8 : INV_X1 port map( A => n9, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1109 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1109;

architecture SYN_BEHAVIORAL of FA_1109 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1108 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1108;

architecture SYN_BEHAVIORAL of FA_1108 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1107 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1107;

architecture SYN_BEHAVIORAL of FA_1107 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1106 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1106;

architecture SYN_BEHAVIORAL of FA_1106 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1105 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1105;

architecture SYN_BEHAVIORAL of FA_1105 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n8, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : INV_X1 port map( A => n7, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n8);
   U7 : XNOR2_X1 port map( A => B, B => n8, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1104 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1104;

architecture SYN_BEHAVIORAL of FA_1104 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1103 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1103;

architecture SYN_BEHAVIORAL of FA_1103 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1102 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1102;

architecture SYN_BEHAVIORAL of FA_1102 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : OAI22_X1 port map( A1 => n5, A2 => n9, B1 => n6, B2 => n7, ZN => Co);
   U4 : INV_X1 port map( A => n4, ZN => n5);
   U5 : INV_X1 port map( A => Ci, ZN => n6);
   U6 : INV_X1 port map( A => n8, ZN => n7);
   U7 : INV_X1 port map( A => A, ZN => n9);
   U8 : XNOR2_X1 port map( A => n9, B => B, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1101 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1101;

architecture SYN_BEHAVIORAL of FA_1101 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1100 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1100;

architecture SYN_BEHAVIORAL of FA_1100 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1099 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1099;

architecture SYN_BEHAVIORAL of FA_1099 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1098 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1098;

architecture SYN_BEHAVIORAL of FA_1098 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => n6, B => B, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1097 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1097;

architecture SYN_BEHAVIORAL of FA_1097 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n8, B1 => n5, B2 => n6, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : INV_X1 port map( A => n7, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n8);
   U7 : XNOR2_X1 port map( A => B, B => n8, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1096 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1096;

architecture SYN_BEHAVIORAL of FA_1096 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n8);
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U2 : OAI22_X1 port map( A1 => n4, A2 => n5, B1 => n6, B2 => n7, ZN => Co);
   U5 : INV_X1 port map( A => B, ZN => n4);
   U6 : INV_X1 port map( A => A, ZN => n5);
   U7 : INV_X1 port map( A => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1095 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1095;

architecture SYN_BEHAVIORAL of FA_1095 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1094 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1094;

architecture SYN_BEHAVIORAL of FA_1094 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : AOI22_X1 port map( A1 => n6, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => B, B => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1093 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1093;

architecture SYN_BEHAVIORAL of FA_1093 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n8, B => n6, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : AOI22_X1 port map( A1 => n4, A2 => A, B1 => Ci, B2 => n6, ZN => n5);
   U5 : INV_X1 port map( A => n5, ZN => Co);
   U6 : CLKBUF_X1 port map( A => Ci, Z => n8);
   U7 : XNOR2_X1 port map( A => B, B => n7, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1092 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1092;

architecture SYN_BEHAVIORAL of FA_1092 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1091 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1091;

architecture SYN_BEHAVIORAL of FA_1091 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => n7, A2 => A, B1 => Ci, B2 => n5, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1090 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1090;

architecture SYN_BEHAVIORAL of FA_1090 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : XNOR2_X1 port map( A => B, B => n6, ZN => n4);
   U4 : AOI22_X1 port map( A1 => n5, A2 => A, B1 => Ci, B2 => n4, ZN => n2);
   U5 : CLKBUF_X1 port map( A => B, Z => n5);
   U6 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1089 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1089;

architecture SYN_BEHAVIORAL of FA_1089 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net69052, net71649, n4, n6, n7, n8 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n4);
   U2 : OR2_X1 port map( A1 => n8, A2 => n6, ZN => Co);
   U3 : AND2_X1 port map( A1 => A, A2 => n4, ZN => n6);
   U4 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);
   U5 : CLKBUF_X1 port map( A => Ci, Z => net71649);
   U6 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U7 : INV_X1 port map( A => net71649, ZN => net69052);
   U8 : NOR2_X1 port map( A1 => net69052, A2 => n7, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1088 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1088;

architecture SYN_BEHAVIORAL of FA_1088 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1087 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1087;

architecture SYN_BEHAVIORAL of FA_1087 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1086 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1086;

architecture SYN_BEHAVIORAL of FA_1086 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1085 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1085;

architecture SYN_BEHAVIORAL of FA_1085 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1084 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1084;

architecture SYN_BEHAVIORAL of FA_1084 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1083 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1083;

architecture SYN_BEHAVIORAL of FA_1083 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1082 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1082;

architecture SYN_BEHAVIORAL of FA_1082 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1081 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1081;

architecture SYN_BEHAVIORAL of FA_1081 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1080 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1080;

architecture SYN_BEHAVIORAL of FA_1080 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1079 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1079;

architecture SYN_BEHAVIORAL of FA_1079 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1078 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1078;

architecture SYN_BEHAVIORAL of FA_1078 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1077 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1077;

architecture SYN_BEHAVIORAL of FA_1077 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1076 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1076;

architecture SYN_BEHAVIORAL of FA_1076 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1075 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1075;

architecture SYN_BEHAVIORAL of FA_1075 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1074 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1074;

architecture SYN_BEHAVIORAL of FA_1074 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1073 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1073;

architecture SYN_BEHAVIORAL of FA_1073 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1072 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1072;

architecture SYN_BEHAVIORAL of FA_1072 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1071 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1071;

architecture SYN_BEHAVIORAL of FA_1071 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1070 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1070;

architecture SYN_BEHAVIORAL of FA_1070 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1069 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1069;

architecture SYN_BEHAVIORAL of FA_1069 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1068 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1068;

architecture SYN_BEHAVIORAL of FA_1068 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1067 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1067;

architecture SYN_BEHAVIORAL of FA_1067 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1066 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1066;

architecture SYN_BEHAVIORAL of FA_1066 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1065 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1065;

architecture SYN_BEHAVIORAL of FA_1065 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1064 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1064;

architecture SYN_BEHAVIORAL of FA_1064 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1063 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1063;

architecture SYN_BEHAVIORAL of FA_1063 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1062 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1062;

architecture SYN_BEHAVIORAL of FA_1062 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1061 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1061;

architecture SYN_BEHAVIORAL of FA_1061 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1060 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1060;

architecture SYN_BEHAVIORAL of FA_1060 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1059 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1059;

architecture SYN_BEHAVIORAL of FA_1059 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1058 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1058;

architecture SYN_BEHAVIORAL of FA_1058 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1057 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1057;

architecture SYN_BEHAVIORAL of FA_1057 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1056 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1056;

architecture SYN_BEHAVIORAL of FA_1056 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1055 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1055;

architecture SYN_BEHAVIORAL of FA_1055 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1054 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1054;

architecture SYN_BEHAVIORAL of FA_1054 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1053 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1053;

architecture SYN_BEHAVIORAL of FA_1053 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1052 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1052;

architecture SYN_BEHAVIORAL of FA_1052 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : CLKBUF_X1 port map( A => n5, Z => n4);
   U2 : INV_X1 port map( A => n6, ZN => Co);
   U5 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1051 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1051;

architecture SYN_BEHAVIORAL of FA_1051 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1050 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1050;

architecture SYN_BEHAVIORAL of FA_1050 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1049 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1049;

architecture SYN_BEHAVIORAL of FA_1049 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1048 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1048;

architecture SYN_BEHAVIORAL of FA_1048 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1047 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1047;

architecture SYN_BEHAVIORAL of FA_1047 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n8);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n5, B1 => n6, B2 => n7, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U5 : INV_X1 port map( A => A, ZN => n5);
   U6 : INV_X1 port map( A => n8, ZN => n6);
   U7 : INV_X1 port map( A => Ci, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1046 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1046;

architecture SYN_BEHAVIORAL of FA_1046 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : CLKBUF_X1 port map( A => Ci, Z => n4);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1045 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1045;

architecture SYN_BEHAVIORAL of FA_1045 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n8);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n5, B1 => n6, B2 => n7, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U5 : INV_X1 port map( A => A, ZN => n5);
   U6 : INV_X1 port map( A => n8, ZN => n6);
   U7 : INV_X1 port map( A => Ci, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1044 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1044;

architecture SYN_BEHAVIORAL of FA_1044 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1043 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1043;

architecture SYN_BEHAVIORAL of FA_1043 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1042 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1042;

architecture SYN_BEHAVIORAL of FA_1042 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U1 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U2 : INV_X1 port map( A => n5, ZN => Co);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1041 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1041;

architecture SYN_BEHAVIORAL of FA_1041 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n9 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n9);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n5, B1 => n6, B2 => n7, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U5 : INV_X1 port map( A => A, ZN => n5);
   U6 : INV_X1 port map( A => n9, ZN => n6);
   U7 : INV_X1 port map( A => Ci, ZN => n7);
   U8 : CLKBUF_X1 port map( A => n9, Z => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1040 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1040;

architecture SYN_BEHAVIORAL of FA_1040 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1039 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1039;

architecture SYN_BEHAVIORAL of FA_1039 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : CLKBUF_X1 port map( A => Ci, Z => n4);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1038 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1038;

architecture SYN_BEHAVIORAL of FA_1038 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : INV_X1 port map( A => n5, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n4, B2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1037 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1037;

architecture SYN_BEHAVIORAL of FA_1037 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n8);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n5, B1 => n6, B2 => n7, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U5 : INV_X1 port map( A => A, ZN => n5);
   U6 : INV_X1 port map( A => Ci, ZN => n6);
   U7 : INV_X1 port map( A => n8, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1036 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1036;

architecture SYN_BEHAVIORAL of FA_1036 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n4, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1035 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1035;

architecture SYN_BEHAVIORAL of FA_1035 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U2 : CLKBUF_X1 port map( A => Ci, Z => n4);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1034 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1034;

architecture SYN_BEHAVIORAL of FA_1034 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : AOI22_X1 port map( A1 => B, A2 => A, B1 => Ci, B2 => n5, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1033 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1033;

architecture SYN_BEHAVIORAL of FA_1033 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n5, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U2 : CLKBUF_X1 port map( A => Ci, Z => n4);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1032 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1032;

architecture SYN_BEHAVIORAL of FA_1032 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n6);
   U2 : CLKBUF_X1 port map( A => n5, Z => n4);
   U5 : INV_X1 port map( A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1031 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1031;

architecture SYN_BEHAVIORAL of FA_1031 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n9, n10 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n9, B => n8, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n10);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n5, B1 => n6, B2 => n7, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U5 : INV_X1 port map( A => A, ZN => n5);
   U6 : INV_X1 port map( A => n10, ZN => n6);
   U7 : INV_X1 port map( A => Ci, ZN => n7);
   U8 : CLKBUF_X1 port map( A => n10, Z => n8);
   U9 : CLKBUF_X1 port map( A => Ci, Z => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1030 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1030;

architecture SYN_BEHAVIORAL of FA_1030 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n9, n10 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n9, B => n8, Z => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n10);
   U1 : OAI22_X1 port map( A1 => n4, A2 => n5, B1 => n6, B2 => n7, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n4);
   U5 : INV_X1 port map( A => A, ZN => n5);
   U6 : INV_X1 port map( A => n10, ZN => n6);
   U7 : INV_X1 port map( A => Ci, ZN => n7);
   U8 : CLKBUF_X1 port map( A => n10, Z => n8);
   U9 : CLKBUF_X1 port map( A => Ci, Z => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1029 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1029;

architecture SYN_BEHAVIORAL of FA_1029 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net69181, n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => net69181, B => n5, Z => S);
   U1 : NOR2_X1 port map( A1 => B, A2 => A, ZN => n6);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => n4);
   U4 : NOR2_X1 port map( A1 => n4, A2 => Ci, ZN => n7);
   U5 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U6 : NOR2_X1 port map( A1 => n7, A2 => n6, ZN => Co);
   U7 : CLKBUF_X1 port map( A => Ci, Z => net69181);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1028 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1028;

architecture SYN_BEHAVIORAL of FA_1028 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n5, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n6);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : XNOR2_X1 port map( A => B, B => n6, ZN => n5);
   U6 : CLKBUF_X1 port map( A => Ci, Z => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1027 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1027;

architecture SYN_BEHAVIORAL of FA_1027 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n5, B => n7, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n8);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n6, B2 => Ci, ZN => n4);
   U4 : INV_X1 port map( A => n4, ZN => Co);
   U5 : CLKBUF_X1 port map( A => n6, Z => n5);
   U6 : XNOR2_X1 port map( A => B, B => n8, ZN => n6);
   U7 : CLKBUF_X1 port map( A => Ci, Z => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1026 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1026;

architecture SYN_BEHAVIORAL of FA_1026 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net67696, n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => net67696, B => n5, Z => S);
   U1 : OR2_X1 port map( A1 => A, A2 => B, ZN => n4);
   U2 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U4 : OAI21_X1 port map( B1 => n7, B2 => Ci, A => n4, ZN => n6);
   U5 : INV_X1 port map( A => n6, ZN => Co);
   U6 : AND2_X1 port map( A1 => A, A2 => B, ZN => n7);
   U7 : CLKBUF_X1 port map( A => Ci, Z => net67696);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1025 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1025;

architecture SYN_BEHAVIORAL of FA_1025 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net66690, net73549, net73544, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => net66690, ZN => net73544);
   U2 : OR2_X1 port map( A1 => n7, A2 => n5, ZN => Co);
   U3 : AND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : XNOR2_X1 port map( A => n6, B => Ci, ZN => S);
   U5 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U6 : CLKBUF_X1 port map( A => n6, Z => net73549);
   U7 : CLKBUF_X1 port map( A => Ci, Z => net66690);
   U8 : NOR2_X1 port map( A1 => net73549, A2 => net73544, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity MUX51_MuxNbit64_31 is

   port( zeroSignal, A_signal, A_neg, A_shifted, A_neg_shifted : in 
         std_logic_vector (63 downto 0);  Sel : in std_logic_vector (2 downto 
         0);  Y : out std_logic_vector (63 downto 0));

end MUX51_MuxNbit64_31;

architecture SYN_BEHAVIORAL_2 of MUX51_MuxNbit64_31 is

   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X4
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X8
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, 
      n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, 
      n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, 
      n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, 
      n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, 
      n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, 
      n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, 
      n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, 
      n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, 
      n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, 
      n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, 
      n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, 
      n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, 
      n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, 
      n308, n309, n310, n311, n312, n313, n314 : std_logic;

begin
   
   U1 : NOR3_X1 port map( A1 => n313, A2 => Sel(2), A3 => n314, ZN => n310);
   U2 : BUF_X1 port map( A => n165, Z => n156);
   U3 : CLKBUF_X1 port map( A => n144, Z => n164);
   U4 : NOR3_X1 port map( A1 => Sel(0), A2 => Sel(2), A3 => n314, ZN => n307);
   U5 : BUF_X1 port map( A => n179, Z => n153);
   U6 : CLKBUF_X1 port map( A => n165, Z => n157);
   U7 : BUF_X8 port map( A => n156, Z => n158);
   U8 : NOR3_X1 port map( A1 => n313, A2 => Sel(2), A3 => n314, ZN => n141);
   U9 : CLKBUF_X1 port map( A => n310, Z => n152);
   U10 : CLKBUF_X1 port map( A => n164, Z => n142);
   U11 : CLKBUF_X1 port map( A => n144, Z => n163);
   U12 : BUF_X4 port map( A => n164, Z => n162);
   U13 : BUF_X4 port map( A => n164, Z => n161);
   U14 : INV_X1 port map( A => n314, ZN => n143);
   U15 : BUF_X1 port map( A => n167, Z => n150);
   U16 : CLKBUF_X1 port map( A => n166, Z => n168);
   U17 : BUF_X1 port map( A => n178, Z => n176);
   U18 : NOR3_X1 port map( A1 => n143, A2 => Sel(2), A3 => n313, ZN => n144);
   U19 : BUF_X1 port map( A => n150, Z => n147);
   U20 : BUF_X1 port map( A => n150, Z => n149);
   U21 : BUF_X1 port map( A => n150, Z => n148);
   U22 : BUF_X1 port map( A => n151, Z => n145);
   U23 : BUF_X1 port map( A => n151, Z => n146);
   U24 : BUF_X1 port map( A => n167, Z => n151);
   U25 : BUF_X1 port map( A => n168, Z => n167);
   U26 : BUF_X1 port map( A => n177, Z => n172);
   U27 : BUF_X1 port map( A => n177, Z => n171);
   U28 : BUF_X1 port map( A => n176, Z => n174);
   U29 : BUF_X1 port map( A => n176, Z => n173);
   U30 : BUF_X1 port map( A => n177, Z => n170);
   U31 : BUF_X1 port map( A => n176, Z => n175);
   U32 : CLKBUF_X1 port map( A => n308, Z => n166);
   U33 : BUF_X1 port map( A => n178, Z => n177);
   U34 : INV_X1 port map( A => Sel(1), ZN => n314);
   U35 : BUF_X1 port map( A => n309, Z => n178);
   U36 : NOR2_X1 port map( A1 => n148, A2 => n180, ZN => n309);
   U37 : AOI22_X1 port map( A1 => A_neg(3), A2 => n307, B1 => A_signal(3), B2 
                           => n144, ZN => n248);
   U38 : AOI222_X1 port map( A1 => A_shifted(2), A2 => n154, B1 => 
                           zeroSignal(2), B2 => n171, C1 => A_neg_shifted(2), 
                           C2 => n148, ZN => n225);
   U39 : AOI222_X1 port map( A1 => A_shifted(4), A2 => n310, B1 => 
                           zeroSignal(4), B2 => n173, C1 => A_neg_shifted(4), 
                           C2 => n166, ZN => n269);
   U40 : AOI222_X1 port map( A1 => A_shifted(37), A2 => n154, B1 => 
                           zeroSignal(37), B2 => n172, C1 => A_neg_shifted(37),
                           C2 => n147, ZN => n241);
   U41 : AOI22_X1 port map( A1 => A_neg(37), A2 => n158, B1 => A_signal(37), B2
                           => n162, ZN => n242);
   U42 : NAND2_X1 port map( A1 => n304, A2 => n303, ZN => Y(7));
   U43 : NAND2_X1 port map( A1 => n244, A2 => n243, ZN => Y(38));
   U44 : AOI222_X1 port map( A1 => A_shifted(38), A2 => n155, B1 => 
                           zeroSignal(38), B2 => n172, C1 => A_neg_shifted(38),
                           C2 => n147, ZN => n243);
   U45 : AOI22_X1 port map( A1 => A_neg(38), A2 => n158, B1 => A_signal(38), B2
                           => n162, ZN => n244);
   U46 : NAND2_X1 port map( A1 => n188, A2 => n187, ZN => Y(12));
   U47 : AOI22_X1 port map( A1 => A_neg(12), A2 => n158, B1 => A_signal(12), B2
                           => n162, ZN => n188);
   U48 : NAND2_X1 port map( A1 => n312, A2 => n311, ZN => Y(9));
   U49 : NAND2_X1 port map( A1 => n292, A2 => n291, ZN => Y(5));
   U50 : NAND2_X1 port map( A1 => n186, A2 => n185, ZN => Y(11));
   U51 : NAND2_X1 port map( A1 => n190, A2 => n189, ZN => Y(13));
   U52 : AOI222_X1 port map( A1 => A_shifted(13), A2 => n155, B1 => 
                           zeroSignal(13), B2 => n170, C1 => A_neg_shifted(13),
                           C2 => n167, ZN => n189);
   U53 : AOI22_X1 port map( A1 => A_neg(13), A2 => n158, B1 => A_signal(13), B2
                           => n161, ZN => n190);
   U54 : NAND2_X1 port map( A1 => n192, A2 => n191, ZN => Y(14));
   U55 : AOI222_X1 port map( A1 => A_shifted(14), A2 => n155, B1 => 
                           zeroSignal(14), B2 => n170, C1 => A_neg_shifted(14),
                           C2 => n167, ZN => n191);
   U56 : AOI22_X1 port map( A1 => A_neg(14), A2 => n158, B1 => A_signal(14), B2
                           => n161, ZN => n192);
   U57 : NAND2_X1 port map( A1 => n194, A2 => n193, ZN => Y(15));
   U58 : AOI222_X1 port map( A1 => A_shifted(15), A2 => n155, B1 => 
                           zeroSignal(15), B2 => n170, C1 => A_neg_shifted(15),
                           C2 => n167, ZN => n193);
   U59 : AOI22_X1 port map( A1 => A_neg(15), A2 => n158, B1 => A_signal(15), B2
                           => n161, ZN => n194);
   U60 : NAND2_X1 port map( A1 => n200, A2 => n199, ZN => Y(18));
   U61 : AOI222_X1 port map( A1 => A_shifted(18), A2 => n155, B1 => 
                           zeroSignal(18), B2 => n170, C1 => A_neg_shifted(18),
                           C2 => n148, ZN => n199);
   U62 : AOI22_X1 port map( A1 => A_neg(18), A2 => n158, B1 => A_signal(18), B2
                           => n161, ZN => n200);
   U63 : NAND2_X1 port map( A1 => n198, A2 => n197, ZN => Y(17));
   U64 : AOI22_X1 port map( A1 => A_neg(17), A2 => n158, B1 => A_signal(17), B2
                           => n161, ZN => n198);
   U65 : NAND2_X1 port map( A1 => n246, A2 => n245, ZN => Y(39));
   U66 : AOI222_X1 port map( A1 => A_shifted(39), A2 => n154, B1 => 
                           zeroSignal(39), B2 => n172, C1 => A_neg_shifted(39),
                           C2 => n147, ZN => n245);
   U67 : NAND2_X1 port map( A1 => n202, A2 => n201, ZN => Y(19));
   U68 : AOI222_X1 port map( A1 => A_shifted(19), A2 => n155, B1 => 
                           zeroSignal(19), B2 => n170, C1 => A_neg_shifted(19),
                           C2 => n147, ZN => n201);
   U69 : AOI22_X1 port map( A1 => A_neg(19), A2 => n158, B1 => A_signal(19), B2
                           => n161, ZN => n202);
   U70 : NAND2_X1 port map( A1 => n196, A2 => n195, ZN => Y(16));
   U71 : AOI222_X1 port map( A1 => A_shifted(16), A2 => n155, B1 => 
                           zeroSignal(16), B2 => n170, C1 => A_neg_shifted(16),
                           C2 => n147, ZN => n195);
   U72 : NAND2_X1 port map( A1 => n288, A2 => n287, ZN => Y(58));
   U73 : AOI222_X1 port map( A1 => A_shifted(58), A2 => n155, B1 => 
                           zeroSignal(58), B2 => n174, C1 => A_neg_shifted(58),
                           C2 => n145, ZN => n287);
   U74 : AOI22_X1 port map( A1 => A_neg(58), A2 => n157, B1 => A_signal(58), B2
                           => n162, ZN => n288);
   U75 : NAND2_X1 port map( A1 => n286, A2 => n285, ZN => Y(57));
   U76 : AOI222_X1 port map( A1 => A_shifted(57), A2 => n154, B1 => 
                           zeroSignal(57), B2 => n174, C1 => A_neg_shifted(57),
                           C2 => n145, ZN => n285);
   U77 : AOI22_X1 port map( A1 => A_neg(57), A2 => n158, B1 => A_signal(57), B2
                           => n162, ZN => n286);
   U78 : NAND2_X1 port map( A1 => n208, A2 => n207, ZN => Y(21));
   U79 : AOI22_X1 port map( A1 => A_neg(21), A2 => n158, B1 => A_signal(21), B2
                           => n161, ZN => n208);
   U80 : NAND2_X1 port map( A1 => n290, A2 => n289, ZN => Y(59));
   U81 : AOI222_X1 port map( A1 => A_shifted(59), A2 => n155, B1 => 
                           zeroSignal(59), B2 => n174, C1 => A_neg_shifted(59),
                           C2 => n145, ZN => n289);
   U82 : AOI22_X1 port map( A1 => A_neg(59), A2 => n158, B1 => A_signal(59), B2
                           => n161, ZN => n290);
   U83 : NAND2_X1 port map( A1 => n294, A2 => n293, ZN => Y(60));
   U84 : AOI222_X1 port map( A1 => A_shifted(60), A2 => n154, B1 => 
                           zeroSignal(60), B2 => n174, C1 => A_neg_shifted(60),
                           C2 => n145, ZN => n293);
   U85 : AOI22_X1 port map( A1 => A_neg(60), A2 => n157, B1 => A_signal(60), B2
                           => n162, ZN => n294);
   U86 : NAND2_X1 port map( A1 => n284, A2 => n283, ZN => Y(56));
   U87 : AOI22_X1 port map( A1 => A_neg(56), A2 => n158, B1 => A_signal(56), B2
                           => n161, ZN => n284);
   U88 : NAND2_X1 port map( A1 => n210, A2 => n209, ZN => Y(22));
   U89 : AOI222_X1 port map( A1 => A_shifted(22), A2 => n155, B1 => 
                           zeroSignal(22), B2 => n171, C1 => A_neg_shifted(22),
                           C2 => n147, ZN => n209);
   U90 : AOI22_X1 port map( A1 => A_neg(22), A2 => n158, B1 => A_signal(22), B2
                           => n161, ZN => n210);
   U91 : NAND2_X1 port map( A1 => n206, A2 => n205, ZN => Y(20));
   U92 : AOI222_X1 port map( A1 => A_shifted(20), A2 => n155, B1 => 
                           zeroSignal(20), B2 => n171, C1 => A_neg_shifted(20),
                           C2 => n147, ZN => n205);
   U93 : NAND2_X1 port map( A1 => n212, A2 => n211, ZN => Y(23));
   U94 : AOI222_X1 port map( A1 => A_shifted(23), A2 => n155, B1 => 
                           zeroSignal(23), B2 => n171, C1 => A_neg_shifted(23),
                           C2 => n147, ZN => n211);
   U95 : AOI22_X1 port map( A1 => A_neg(23), A2 => n158, B1 => A_signal(23), B2
                           => n161, ZN => n212);
   U96 : NAND2_X1 port map( A1 => n298, A2 => n297, ZN => Y(62));
   U97 : AOI222_X1 port map( A1 => A_shifted(62), A2 => n154, B1 => 
                           zeroSignal(62), B2 => n174, C1 => A_neg_shifted(62),
                           C2 => n145, ZN => n297);
   U98 : AOI22_X1 port map( A1 => A_neg(62), A2 => n158, B1 => A_signal(62), B2
                           => n162, ZN => n298);
   U99 : NAND2_X1 port map( A1 => n296, A2 => n295, ZN => Y(61));
   U100 : AOI222_X1 port map( A1 => A_shifted(61), A2 => n155, B1 => 
                           zeroSignal(61), B2 => n174, C1 => A_neg_shifted(61),
                           C2 => n145, ZN => n295);
   U101 : AOI22_X1 port map( A1 => A_neg(61), A2 => n158, B1 => A_signal(61), 
                           B2 => n161, ZN => n296);
   U102 : NAND2_X1 port map( A1 => n214, A2 => n213, ZN => Y(24));
   U103 : AOI222_X1 port map( A1 => A_shifted(24), A2 => n154, B1 => 
                           zeroSignal(24), B2 => n171, C1 => A_neg_shifted(24),
                           C2 => n148, ZN => n213);
   U104 : AOI22_X1 port map( A1 => A_neg(24), A2 => n158, B1 => A_signal(24), 
                           B2 => n161, ZN => n214);
   U105 : NAND2_X1 port map( A1 => n300, A2 => n299, ZN => Y(63));
   U106 : AOI222_X1 port map( A1 => A_shifted(63), A2 => n155, B1 => 
                           zeroSignal(63), B2 => n174, C1 => A_neg_shifted(63),
                           C2 => n145, ZN => n299);
   U107 : AOI22_X1 port map( A1 => A_neg(63), A2 => n157, B1 => A_signal(63), 
                           B2 => n162, ZN => n300);
   U108 : NAND2_X1 port map( A1 => n260, A2 => n259, ZN => Y(45));
   U109 : AOI222_X1 port map( A1 => A_shifted(45), A2 => n154, B1 => 
                           zeroSignal(45), B2 => n173, C1 => A_neg_shifted(45),
                           C2 => n146, ZN => n259);
   U110 : AOI22_X1 port map( A1 => A_neg(45), A2 => n157, B1 => A_signal(45), 
                           B2 => n161, ZN => n260);
   U111 : NAND2_X1 port map( A1 => n256, A2 => n255, ZN => Y(43));
   U112 : AOI222_X1 port map( A1 => A_shifted(43), A2 => n154, B1 => 
                           zeroSignal(43), B2 => n173, C1 => A_neg_shifted(43),
                           C2 => n146, ZN => n255);
   U113 : AOI22_X1 port map( A1 => A_neg(43), A2 => n157, B1 => A_signal(43), 
                           B2 => n161, ZN => n256);
   U114 : NAND2_X1 port map( A1 => n216, A2 => n215, ZN => Y(25));
   U115 : AOI222_X1 port map( A1 => A_shifted(25), A2 => n155, B1 => 
                           zeroSignal(25), B2 => n171, C1 => A_neg_shifted(25),
                           C2 => n148, ZN => n215);
   U116 : AOI22_X1 port map( A1 => A_neg(25), A2 => n158, B1 => A_signal(25), 
                           B2 => n161, ZN => n216);
   U117 : NAND2_X1 port map( A1 => n220, A2 => n219, ZN => Y(27));
   U118 : AOI22_X1 port map( A1 => A_neg(27), A2 => n158, B1 => A_signal(27), 
                           B2 => n161, ZN => n220);
   U119 : NAND2_X1 port map( A1 => n276, A2 => n275, ZN => Y(52));
   U120 : AOI222_X1 port map( A1 => A_shifted(52), A2 => n155, B1 => 
                           zeroSignal(52), B2 => n173, C1 => A_neg_shifted(52),
                           C2 => n146, ZN => n275);
   U121 : NAND2_X1 port map( A1 => n262, A2 => n261, ZN => Y(46));
   U122 : AOI222_X1 port map( A1 => A_shifted(46), A2 => n155, B1 => 
                           zeroSignal(46), B2 => n173, C1 => A_neg_shifted(46),
                           C2 => n146, ZN => n261);
   U123 : NAND2_X1 port map( A1 => n218, A2 => n217, ZN => Y(26));
   U124 : AOI222_X1 port map( A1 => A_shifted(26), A2 => n154, B1 => 
                           zeroSignal(26), B2 => n171, C1 => A_neg_shifted(26),
                           C2 => n148, ZN => n217);
   U125 : NAND2_X1 port map( A1 => n268, A2 => n267, ZN => Y(49));
   U126 : NAND2_X1 port map( A1 => n222, A2 => n221, ZN => Y(28));
   U127 : AOI222_X1 port map( A1 => A_shifted(28), A2 => n154, B1 => 
                           zeroSignal(28), B2 => n171, C1 => A_neg_shifted(28),
                           C2 => n148, ZN => n221);
   U128 : AOI22_X1 port map( A1 => A_neg(28), A2 => n157, B1 => A_signal(28), 
                           B2 => n162, ZN => n222);
   U129 : NAND2_X1 port map( A1 => n224, A2 => n223, ZN => Y(29));
   U130 : AOI222_X1 port map( A1 => A_shifted(29), A2 => n155, B1 => 
                           zeroSignal(29), B2 => n171, C1 => A_neg_shifted(29),
                           C2 => n148, ZN => n223);
   U131 : AOI22_X1 port map( A1 => A_neg(29), A2 => n158, B1 => A_signal(29), 
                           B2 => n162, ZN => n224);
   U132 : NAND2_X1 port map( A1 => n238, A2 => n237, ZN => Y(35));
   U133 : AOI222_X1 port map( A1 => A_shifted(35), A2 => n154, B1 => 
                           zeroSignal(35), B2 => n172, C1 => A_neg_shifted(35),
                           C2 => n147, ZN => n237);
   U134 : AOI22_X1 port map( A1 => A_neg(35), A2 => n158, B1 => A_signal(35), 
                           B2 => n162, ZN => n238);
   U135 : NAND2_X1 port map( A1 => n258, A2 => n257, ZN => Y(44));
   U136 : AOI22_X1 port map( A1 => A_neg(44), A2 => n157, B1 => A_signal(44), 
                           B2 => n162, ZN => n258);
   U137 : AOI222_X1 port map( A1 => A_shifted(44), A2 => n155, B1 => 
                           zeroSignal(44), B2 => n173, C1 => A_neg_shifted(44),
                           C2 => n146, ZN => n257);
   U138 : NAND2_X1 port map( A1 => n266, A2 => n265, ZN => Y(48));
   U139 : AOI222_X1 port map( A1 => A_shifted(48), A2 => n154, B1 => 
                           zeroSignal(48), B2 => n173, C1 => A_neg_shifted(48),
                           C2 => n146, ZN => n265);
   U140 : NAND2_X1 port map( A1 => n228, A2 => n227, ZN => Y(30));
   U141 : AOI222_X1 port map( A1 => A_shifted(30), A2 => n154, B1 => 
                           zeroSignal(30), B2 => n171, C1 => A_neg_shifted(30),
                           C2 => n148, ZN => n227);
   U142 : AOI22_X1 port map( A1 => A_neg(30), A2 => n157, B1 => A_signal(30), 
                           B2 => n161, ZN => n228);
   U143 : NAND2_X1 port map( A1 => n272, A2 => n271, ZN => Y(50));
   U144 : NAND2_X1 port map( A1 => n282, A2 => n281, ZN => Y(55));
   U145 : AOI222_X1 port map( A1 => A_shifted(55), A2 => n154, B1 => 
                           zeroSignal(55), B2 => n174, C1 => A_neg_shifted(55),
                           C2 => n145, ZN => n281);
   U146 : NAND2_X1 port map( A1 => n230, A2 => n229, ZN => Y(31));
   U147 : AOI222_X1 port map( A1 => A_shifted(31), A2 => n155, B1 => 
                           zeroSignal(31), B2 => n172, C1 => A_neg_shifted(31),
                           C2 => n148, ZN => n229);
   U148 : AOI22_X1 port map( A1 => A_neg(31), A2 => n158, B1 => A_signal(31), 
                           B2 => n162, ZN => n230);
   U149 : NAND2_X1 port map( A1 => n278, A2 => n277, ZN => Y(53));
   U150 : AOI22_X1 port map( A1 => A_neg(53), A2 => n157, B1 => A_signal(53), 
                           B2 => n161, ZN => n278);
   U151 : NAND2_X1 port map( A1 => n232, A2 => n231, ZN => Y(32));
   U152 : AOI222_X1 port map( A1 => A_shifted(32), A2 => n154, B1 => 
                           zeroSignal(32), B2 => n172, C1 => A_neg_shifted(32),
                           C2 => n148, ZN => n231);
   U153 : AOI22_X1 port map( A1 => A_neg(32), A2 => n157, B1 => A_signal(32), 
                           B2 => n162, ZN => n232);
   U154 : NAND2_X1 port map( A1 => n234, A2 => n233, ZN => Y(33));
   U155 : AOI222_X1 port map( A1 => A_shifted(33), A2 => n155, B1 => 
                           zeroSignal(33), B2 => n172, C1 => A_neg_shifted(33),
                           C2 => n148, ZN => n233);
   U156 : AOI22_X1 port map( A1 => A_neg(33), A2 => n158, B1 => A_signal(33), 
                           B2 => n161, ZN => n234);
   U157 : NAND2_X1 port map( A1 => n264, A2 => n263, ZN => Y(47));
   U158 : AOI22_X1 port map( A1 => A_neg(47), A2 => n157, B1 => A_signal(47), 
                           B2 => n162, ZN => n264);
   U159 : NAND2_X1 port map( A1 => n280, A2 => n279, ZN => Y(54));
   U160 : AOI222_X1 port map( A1 => A_shifted(54), A2 => n155, B1 => 
                           zeroSignal(54), B2 => n174, C1 => A_neg_shifted(54),
                           C2 => n145, ZN => n279);
   U161 : AOI22_X1 port map( A1 => A_neg(54), A2 => n158, B1 => A_signal(54), 
                           B2 => n162, ZN => n280);
   U162 : NAND2_X1 port map( A1 => n236, A2 => n235, ZN => Y(34));
   U163 : AOI222_X1 port map( A1 => A_shifted(34), A2 => n155, B1 => 
                           zeroSignal(34), B2 => n172, C1 => A_neg_shifted(34),
                           C2 => n145, ZN => n235);
   U164 : AOI22_X1 port map( A1 => A_neg(34), A2 => n157, B1 => A_signal(34), 
                           B2 => n162, ZN => n236);
   U165 : NAND2_X1 port map( A1 => n274, A2 => n273, ZN => Y(51));
   U166 : AOI22_X1 port map( A1 => A_neg(51), A2 => n158, B1 => A_signal(51), 
                           B2 => n162, ZN => n274);
   U167 : NAND2_X1 port map( A1 => n240, A2 => n239, ZN => Y(36));
   U168 : AOI22_X1 port map( A1 => A_neg(36), A2 => n157, B1 => A_signal(36), 
                           B2 => n161, ZN => n240);
   U169 : AOI222_X1 port map( A1 => A_shifted(36), A2 => n155, B1 => 
                           zeroSignal(36), B2 => n172, C1 => A_neg_shifted(36),
                           C2 => n147, ZN => n239);
   U170 : NAND2_X1 port map( A1 => n250, A2 => n249, ZN => Y(40));
   U171 : AOI22_X1 port map( A1 => A_neg(40), A2 => n158, B1 => A_signal(40), 
                           B2 => n161, ZN => n250);
   U172 : NAND2_X1 port map( A1 => n252, A2 => n251, ZN => Y(41));
   U173 : AOI222_X1 port map( A1 => A_shifted(41), A2 => n154, B1 => 
                           zeroSignal(41), B2 => n172, C1 => A_neg_shifted(41),
                           C2 => n146, ZN => n251);
   U174 : AOI22_X1 port map( A1 => A_neg(41), A2 => n157, B1 => A_signal(41), 
                           B2 => n162, ZN => n252);
   U175 : NAND2_X1 port map( A1 => n254, A2 => n253, ZN => Y(42));
   U176 : AOI222_X1 port map( A1 => A_shifted(42), A2 => n155, B1 => 
                           zeroSignal(42), B2 => n173, C1 => A_neg_shifted(42),
                           C2 => n147, ZN => n253);
   U177 : AOI22_X1 port map( A1 => A_neg(42), A2 => n158, B1 => A_signal(42), 
                           B2 => n162, ZN => n254);
   U178 : NAND2_X1 port map( A1 => n182, A2 => n181, ZN => Y(0));
   U179 : AOI22_X1 port map( A1 => A_neg(0), A2 => n157, B1 => A_signal(0), B2 
                           => n161, ZN => n182);
   U180 : AOI222_X1 port map( A1 => A_shifted(0), A2 => n155, B1 => 
                           zeroSignal(0), B2 => n170, C1 => A_neg_shifted(0), 
                           C2 => n145, ZN => n181);
   U181 : NAND2_X1 port map( A1 => n204, A2 => n203, ZN => Y(1));
   U182 : AOI22_X1 port map( A1 => A_neg(1), A2 => n158, B1 => A_signal(1), B2 
                           => n162, ZN => n204);
   U183 : AOI222_X1 port map( A1 => A_shifted(1), A2 => n154, B1 => 
                           zeroSignal(1), B2 => n170, C1 => A_neg_shifted(1), 
                           C2 => n147, ZN => n203);
   U184 : AOI222_X1 port map( A1 => A_shifted(11), A2 => n155, B1 => 
                           zeroSignal(11), B2 => n170, C1 => A_neg_shifted(11),
                           C2 => n167, ZN => n185);
   U185 : AOI22_X1 port map( A1 => A_neg(10), A2 => n158, B1 => A_signal(10), 
                           B2 => n142, ZN => n184);
   U186 : AOI222_X1 port map( A1 => A_shifted(53), A2 => n154, B1 => 
                           zeroSignal(53), B2 => n174, C1 => A_neg_shifted(53),
                           C2 => n146, ZN => n277);
   U187 : AOI22_X1 port map( A1 => A_neg(52), A2 => n158, B1 => A_signal(52), 
                           B2 => n162, ZN => n276);
   U188 : NAND2_X1 port map( A1 => n306, A2 => n305, ZN => Y(8));
   U189 : AOI222_X1 port map( A1 => A_shifted(56), A2 => n155, B1 => 
                           zeroSignal(56), B2 => n174, C1 => A_neg_shifted(56),
                           C2 => n145, ZN => n283);
   U190 : AOI22_X1 port map( A1 => A_neg(55), A2 => n157, B1 => A_signal(55), 
                           B2 => n162, ZN => n282);
   U191 : AOI222_X1 port map( A1 => A_shifted(51), A2 => n155, B1 => 
                           zeroSignal(51), B2 => n173, C1 => A_neg_shifted(51),
                           C2 => n146, ZN => n273);
   U192 : AOI22_X1 port map( A1 => A_neg(50), A2 => n157, B1 => A_signal(50), 
                           B2 => n161, ZN => n272);
   U193 : AOI222_X1 port map( A1 => A_shifted(49), A2 => n155, B1 => 
                           zeroSignal(49), B2 => n173, C1 => A_neg_shifted(49),
                           C2 => n146, ZN => n267);
   U194 : AOI22_X1 port map( A1 => A_neg(48), A2 => n158, B1 => A_signal(48), 
                           B2 => n161, ZN => n266);
   U195 : AOI222_X1 port map( A1 => A_shifted(10), A2 => n155, B1 => 
                           zeroSignal(10), B2 => n170, C1 => A_neg_shifted(10),
                           C2 => n168, ZN => n183);
   U196 : AOI222_X1 port map( A1 => A_shifted(50), A2 => n154, B1 => 
                           zeroSignal(50), B2 => n173, C1 => A_neg_shifted(50),
                           C2 => n146, ZN => n271);
   U197 : AOI22_X1 port map( A1 => A_neg(49), A2 => n158, B1 => A_signal(49), 
                           B2 => n162, ZN => n268);
   U198 : AOI222_X1 port map( A1 => A_shifted(47), A2 => n155, B1 => 
                           zeroSignal(47), B2 => n173, C1 => A_neg_shifted(47),
                           C2 => n146, ZN => n263);
   U199 : AOI22_X1 port map( A1 => A_neg(46), A2 => n158, B1 => A_signal(46), 
                           B2 => n162, ZN => n262);
   U200 : NAND2_X1 port map( A1 => n226, A2 => n225, ZN => Y(2));
   U201 : NAND2_X1 port map( A1 => n184, A2 => n183, ZN => Y(10));
   U202 : AOI22_X1 port map( A1 => A_neg(2), A2 => n307, B1 => A_signal(2), B2 
                           => n144, ZN => n226);
   U203 : NAND2_X1 port map( A1 => n270, A2 => n269, ZN => Y(4));
   U204 : BUF_X4 port map( A => n152, Z => n154);
   U205 : BUF_X4 port map( A => n153, Z => n155);
   U206 : BUF_X1 port map( A => n310, Z => n179);
   U207 : INV_X1 port map( A => Sel(0), ZN => n313);
   U208 : BUF_X1 port map( A => n307, Z => n165);
   U209 : CLKBUF_X1 port map( A => n166, Z => n159);
   U210 : CLKBUF_X1 port map( A => n166, Z => n160);
   U211 : CLKBUF_X1 port map( A => n166, Z => n169);
   U212 : AOI222_X1 port map( A1 => A_shifted(12), A2 => n155, B1 => 
                           zeroSignal(12), B2 => n170, C1 => A_neg_shifted(12),
                           C2 => n167, ZN => n187);
   U213 : AOI22_X1 port map( A1 => A_neg(11), A2 => n158, B1 => A_signal(11), 
                           B2 => n162, ZN => n186);
   U214 : AOI21_X1 port map( B1 => n313, B2 => n314, A => Sel(2), ZN => n180);
   U215 : AND3_X1 port map( A1 => n313, A2 => n314, A3 => Sel(2), ZN => n308);
   U216 : AOI22_X1 port map( A1 => A_neg(9), A2 => n158, B1 => A_signal(9), B2 
                           => n142, ZN => n312);
   U217 : NAND2_X1 port map( A1 => n242, A2 => n241, ZN => Y(37));
   U218 : AOI222_X1 port map( A1 => A_shifted(9), A2 => n154, B1 => 
                           zeroSignal(9), B2 => n175, C1 => A_neg_shifted(9), 
                           C2 => n168, ZN => n311);
   U219 : AOI22_X1 port map( A1 => A_neg(8), A2 => n158, B1 => A_signal(8), B2 
                           => n142, ZN => n306);
   U220 : NAND2_X1 port map( A1 => n302, A2 => n301, ZN => Y(6));
   U221 : AOI222_X1 port map( A1 => A_shifted(6), A2 => n179, B1 => 
                           zeroSignal(6), B2 => n175, C1 => A_neg_shifted(6), 
                           C2 => n160, ZN => n301);
   U222 : AOI22_X1 port map( A1 => A_neg(5), A2 => n165, B1 => A_signal(5), B2 
                           => n164, ZN => n292);
   U223 : AOI22_X1 port map( A1 => A_neg(39), A2 => n157, B1 => A_signal(39), 
                           B2 => n162, ZN => n246);
   U224 : AOI222_X1 port map( A1 => A_shifted(40), A2 => n154, B1 => 
                           zeroSignal(40), B2 => n172, C1 => A_neg_shifted(40),
                           C2 => n149, ZN => n249);
   U225 : AOI222_X1 port map( A1 => A_shifted(27), A2 => n155, B1 => 
                           zeroSignal(27), B2 => n171, C1 => A_neg_shifted(27),
                           C2 => n149, ZN => n219);
   U226 : AOI22_X1 port map( A1 => A_neg(26), A2 => n158, B1 => A_signal(26), 
                           B2 => n161, ZN => n218);
   U227 : AOI222_X1 port map( A1 => A_shifted(21), A2 => n155, B1 => 
                           zeroSignal(21), B2 => n171, C1 => A_neg_shifted(21),
                           C2 => n149, ZN => n207);
   U228 : AOI22_X1 port map( A1 => A_neg(20), A2 => n158, B1 => A_signal(20), 
                           B2 => n161, ZN => n206);
   U229 : AOI222_X1 port map( A1 => A_shifted(17), A2 => n155, B1 => 
                           zeroSignal(17), B2 => n170, C1 => A_neg_shifted(17),
                           C2 => n149, ZN => n197);
   U230 : AOI22_X1 port map( A1 => A_neg(16), A2 => n158, B1 => A_signal(16), 
                           B2 => n161, ZN => n196);
   U231 : AOI222_X1 port map( A1 => A_shifted(5), A2 => n152, B1 => 
                           zeroSignal(5), B2 => n174, C1 => A_neg_shifted(5), 
                           C2 => n159, ZN => n291);
   U232 : AOI22_X1 port map( A1 => A_neg(4), A2 => n165, B1 => A_signal(4), B2 
                           => n163, ZN => n270);
   U233 : AOI222_X1 port map( A1 => A_shifted(3), A2 => n141, B1 => 
                           zeroSignal(3), B2 => n172, C1 => A_neg_shifted(3), 
                           C2 => n308, ZN => n247);
   U234 : NAND2_X1 port map( A1 => n248, A2 => n247, ZN => Y(3));
   U235 : AOI22_X1 port map( A1 => A_neg(7), A2 => n157, B1 => A_signal(7), B2 
                           => n142, ZN => n304);
   U236 : AOI222_X1 port map( A1 => A_shifted(8), A2 => n153, B1 => 
                           zeroSignal(8), B2 => n175, C1 => A_neg_shifted(8), 
                           C2 => n168, ZN => n305);
   U237 : AOI22_X1 port map( A1 => A_neg(6), A2 => n156, B1 => A_signal(6), B2 
                           => n142, ZN => n302);
   U238 : AOI222_X1 port map( A1 => A_shifted(7), A2 => n153, B1 => 
                           zeroSignal(7), B2 => n175, C1 => A_neg_shifted(7), 
                           C2 => n169, ZN => n303);

end SYN_BEHAVIORAL_2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity MUX51_MuxNbit64_30 is

   port( zeroSignal, A_signal, A_neg, A_shifted, A_neg_shifted : in 
         std_logic_vector (63 downto 0);  Sel : in std_logic_vector (2 downto 
         0);  Y : out std_logic_vector (63 downto 0));

end MUX51_MuxNbit64_30;

architecture SYN_BEHAVIORAL_2 of MUX51_MuxNbit64_30 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, 
      n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, 
      n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, 
      n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, 
      n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, 
      n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, 
      n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, 
      n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, 
      n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, 
      n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, 
      n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, 
      n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, 
      n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, 
      n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, 
      n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319 : 
      std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n196, A2 => n195, ZN => Y(13));
   U2 : CLKBUF_X1 port map( A => n167, Z => n162);
   U3 : CLKBUF_X1 port map( A => n183, Z => n180);
   U4 : CLKBUF_X1 port map( A => n167, Z => n161);
   U5 : CLKBUF_X1 port map( A => n185, Z => n184);
   U6 : CLKBUF_X1 port map( A => n151, Z => n150);
   U7 : CLKBUF_X1 port map( A => n141, Z => n166);
   U8 : CLKBUF_X1 port map( A => n142, Z => n159);
   U9 : BUF_X1 port map( A => n141, Z => n167);
   U10 : BUF_X1 port map( A => n142, Z => n158);
   U11 : BUF_X1 port map( A => n185, Z => n183);
   U12 : BUF_X1 port map( A => n151, Z => n149);
   U13 : BUF_X1 port map( A => n176, Z => n175);
   U14 : AND3_X1 port map( A1 => n318, A2 => n319, A3 => Sel(2), ZN => n141);
   U15 : NOR3_X1 port map( A1 => Sel(0), A2 => Sel(2), A3 => n319, ZN => n142);
   U16 : BUF_X1 port map( A => n315, Z => n185);
   U17 : BUF_X1 port map( A => n313, Z => n151);
   U18 : BUF_X1 port map( A => n167, Z => n160);
   U19 : BUF_X1 port map( A => n149, Z => n147);
   U20 : BUF_X1 port map( A => n183, Z => n181);
   U21 : BUF_X1 port map( A => n149, Z => n146);
   U22 : BUF_X1 port map( A => n183, Z => n182);
   U23 : BUF_X1 port map( A => n149, Z => n148);
   U24 : BUF_X1 port map( A => n158, Z => n156);
   U25 : BUF_X1 port map( A => n158, Z => n155);
   U26 : BUF_X1 port map( A => n158, Z => n157);
   U27 : BUF_X1 port map( A => n184, Z => n177);
   U28 : BUF_X1 port map( A => n150, Z => n143);
   U29 : BUF_X1 port map( A => n166, Z => n165);
   U30 : BUF_X1 port map( A => n159, Z => n152);
   U31 : BUF_X1 port map( A => n166, Z => n164);
   U32 : BUF_X1 port map( A => n150, Z => n144);
   U33 : BUF_X1 port map( A => n184, Z => n178);
   U34 : BUF_X1 port map( A => n159, Z => n153);
   U35 : BUF_X1 port map( A => n166, Z => n163);
   U36 : BUF_X1 port map( A => n150, Z => n145);
   U37 : BUF_X1 port map( A => n184, Z => n179);
   U38 : BUF_X1 port map( A => n159, Z => n154);
   U39 : BUF_X1 port map( A => n174, Z => n172);
   U40 : BUF_X1 port map( A => n175, Z => n168);
   U41 : BUF_X1 port map( A => n175, Z => n169);
   U42 : BUF_X1 port map( A => n175, Z => n170);
   U43 : BUF_X1 port map( A => n174, Z => n171);
   U44 : BUF_X1 port map( A => n174, Z => n173);
   U45 : BUF_X1 port map( A => n176, Z => n174);
   U46 : INV_X1 port map( A => Sel(0), ZN => n318);
   U47 : BUF_X1 port map( A => n314, Z => n176);
   U48 : NOR2_X1 port map( A1 => n165, A2 => n186, ZN => n314);
   U49 : AOI222_X1 port map( A1 => A_shifted(4), A2 => n180, B1 => 
                           zeroSignal(4), B2 => n171, C1 => A_neg_shifted(4), 
                           C2 => n161, ZN => n275);
   U50 : NAND2_X1 port map( A1 => n308, A2 => n307, ZN => Y(6));
   U51 : AOI222_X1 port map( A1 => A_shifted(6), A2 => n182, B1 => 
                           zeroSignal(6), B2 => n173, C1 => A_neg_shifted(6), 
                           C2 => n160, ZN => n307);
   U52 : AOI222_X1 port map( A1 => A_shifted(7), A2 => n182, B1 => 
                           zeroSignal(7), B2 => n173, C1 => A_neg_shifted(7), 
                           C2 => n160, ZN => n309);
   U53 : AOI222_X1 port map( A1 => A_shifted(8), A2 => n182, B1 => 
                           zeroSignal(8), B2 => n173, C1 => A_neg_shifted(8), 
                           C2 => n160, ZN => n311);
   U54 : NAND2_X1 port map( A1 => n200, A2 => n199, ZN => Y(15));
   U55 : AOI22_X1 port map( A1 => A_neg(15), A2 => n152, B1 => A_signal(15), B2
                           => n143, ZN => n200);
   U56 : AOI222_X1 port map( A1 => A_shifted(15), A2 => n177, B1 => 
                           zeroSignal(15), B2 => n168, C1 => A_neg_shifted(15),
                           C2 => n164, ZN => n199);
   U57 : NAND2_X1 port map( A1 => n202, A2 => n201, ZN => Y(16));
   U58 : AOI22_X1 port map( A1 => A_neg(16), A2 => n152, B1 => A_signal(16), B2
                           => n143, ZN => n202);
   U59 : AOI222_X1 port map( A1 => A_shifted(16), A2 => n177, B1 => 
                           zeroSignal(16), B2 => n168, C1 => A_neg_shifted(16),
                           C2 => n164, ZN => n201);
   U60 : NAND2_X1 port map( A1 => n204, A2 => n203, ZN => Y(17));
   U61 : AOI22_X1 port map( A1 => A_neg(17), A2 => n152, B1 => A_signal(17), B2
                           => n143, ZN => n204);
   U62 : AOI222_X1 port map( A1 => A_shifted(17), A2 => n177, B1 => 
                           zeroSignal(17), B2 => n168, C1 => A_neg_shifted(17),
                           C2 => n164, ZN => n203);
   U63 : NAND2_X1 port map( A1 => n206, A2 => n205, ZN => Y(18));
   U64 : AOI222_X1 port map( A1 => A_shifted(18), A2 => n177, B1 => 
                           zeroSignal(18), B2 => n168, C1 => A_neg_shifted(18),
                           C2 => n164, ZN => n205);
   U65 : NAND2_X1 port map( A1 => n212, A2 => n211, ZN => Y(20));
   U66 : AOI22_X1 port map( A1 => A_neg(20), A2 => n153, B1 => A_signal(20), B2
                           => n144, ZN => n212);
   U67 : AOI222_X1 port map( A1 => A_shifted(20), A2 => n178, B1 => 
                           zeroSignal(20), B2 => n169, C1 => A_neg_shifted(20),
                           C2 => n164, ZN => n211);
   U68 : NAND2_X1 port map( A1 => n214, A2 => n213, ZN => Y(21));
   U69 : AOI22_X1 port map( A1 => A_neg(21), A2 => n153, B1 => A_signal(21), B2
                           => n144, ZN => n214);
   U70 : AOI222_X1 port map( A1 => A_shifted(21), A2 => n178, B1 => 
                           zeroSignal(21), B2 => n169, C1 => A_neg_shifted(21),
                           C2 => n164, ZN => n213);
   U71 : NAND2_X1 port map( A1 => n317, A2 => n316, ZN => Y(9));
   U72 : AOI222_X1 port map( A1 => A_shifted(9), A2 => n182, B1 => 
                           zeroSignal(9), B2 => n173, C1 => A_neg_shifted(9), 
                           C2 => n160, ZN => n316);
   U73 : NAND2_X1 port map( A1 => n216, A2 => n215, ZN => Y(22));
   U74 : AOI222_X1 port map( A1 => A_shifted(22), A2 => n178, B1 => 
                           zeroSignal(22), B2 => n169, C1 => A_neg_shifted(22),
                           C2 => n164, ZN => n215);
   U75 : NAND2_X1 port map( A1 => n220, A2 => n219, ZN => Y(24));
   U76 : AOI22_X1 port map( A1 => A_neg(24), A2 => n153, B1 => A_signal(24), B2
                           => n144, ZN => n220);
   U77 : AOI222_X1 port map( A1 => A_shifted(24), A2 => n178, B1 => 
                           zeroSignal(24), B2 => n169, C1 => A_neg_shifted(24),
                           C2 => n163, ZN => n219);
   U78 : NAND2_X1 port map( A1 => n248, A2 => n247, ZN => Y(37));
   U79 : AOI222_X1 port map( A1 => A_shifted(37), A2 => n179, B1 => 
                           zeroSignal(37), B2 => n170, C1 => A_neg_shifted(37),
                           C2 => n162, ZN => n247);
   U80 : AOI22_X1 port map( A1 => A_neg(37), A2 => n154, B1 => A_signal(37), B2
                           => n145, ZN => n248);
   U81 : NAND2_X1 port map( A1 => n222, A2 => n221, ZN => Y(25));
   U82 : AOI22_X1 port map( A1 => A_neg(25), A2 => n153, B1 => A_signal(25), B2
                           => n144, ZN => n222);
   U83 : AOI222_X1 port map( A1 => A_shifted(25), A2 => n178, B1 => 
                           zeroSignal(25), B2 => n169, C1 => A_neg_shifted(25),
                           C2 => n163, ZN => n221);
   U84 : NAND2_X1 port map( A1 => n224, A2 => n223, ZN => Y(26));
   U85 : AOI22_X1 port map( A1 => A_neg(26), A2 => n153, B1 => A_signal(26), B2
                           => n144, ZN => n224);
   U86 : AOI222_X1 port map( A1 => A_shifted(26), A2 => n178, B1 => 
                           zeroSignal(26), B2 => n169, C1 => A_neg_shifted(26),
                           C2 => n163, ZN => n223);
   U87 : NAND2_X1 port map( A1 => n226, A2 => n225, ZN => Y(27));
   U88 : AOI22_X1 port map( A1 => A_neg(27), A2 => n153, B1 => A_signal(27), B2
                           => n144, ZN => n226);
   U89 : AOI222_X1 port map( A1 => A_shifted(27), A2 => n178, B1 => 
                           zeroSignal(27), B2 => n169, C1 => A_neg_shifted(27),
                           C2 => n163, ZN => n225);
   U90 : NAND2_X1 port map( A1 => n228, A2 => n227, ZN => Y(28));
   U91 : AOI222_X1 port map( A1 => A_shifted(28), A2 => n178, B1 => 
                           zeroSignal(28), B2 => n169, C1 => A_neg_shifted(28),
                           C2 => n163, ZN => n227);
   U92 : NAND2_X1 port map( A1 => n234, A2 => n233, ZN => Y(30));
   U93 : AOI22_X1 port map( A1 => A_neg(30), A2 => n153, B1 => A_signal(30), B2
                           => n144, ZN => n234);
   U94 : AOI222_X1 port map( A1 => A_shifted(30), A2 => n178, B1 => 
                           zeroSignal(30), B2 => n169, C1 => A_neg_shifted(30),
                           C2 => n163, ZN => n233);
   U95 : NAND2_X1 port map( A1 => n236, A2 => n235, ZN => Y(31));
   U96 : AOI22_X1 port map( A1 => A_neg(31), A2 => n154, B1 => A_signal(31), B2
                           => n145, ZN => n236);
   U97 : AOI222_X1 port map( A1 => A_shifted(31), A2 => n179, B1 => 
                           zeroSignal(31), B2 => n170, C1 => A_neg_shifted(31),
                           C2 => n163, ZN => n235);
   U98 : NAND2_X1 port map( A1 => n238, A2 => n237, ZN => Y(32));
   U99 : AOI22_X1 port map( A1 => A_neg(32), A2 => n154, B1 => A_signal(32), B2
                           => n145, ZN => n238);
   U100 : AOI222_X1 port map( A1 => A_shifted(32), A2 => n179, B1 => 
                           zeroSignal(32), B2 => n170, C1 => A_neg_shifted(32),
                           C2 => n163, ZN => n237);
   U101 : NAND2_X1 port map( A1 => n190, A2 => n189, ZN => Y(10));
   U102 : AOI222_X1 port map( A1 => A_shifted(10), A2 => n177, B1 => 
                           zeroSignal(10), B2 => n168, C1 => A_neg_shifted(10),
                           C2 => n165, ZN => n189);
   U103 : NAND2_X1 port map( A1 => n240, A2 => n239, ZN => Y(33));
   U104 : AOI22_X1 port map( A1 => A_neg(33), A2 => n154, B1 => A_signal(33), 
                           B2 => n145, ZN => n240);
   U105 : AOI222_X1 port map( A1 => A_shifted(33), A2 => n179, B1 => 
                           zeroSignal(33), B2 => n170, C1 => A_neg_shifted(33),
                           C2 => n163, ZN => n239);
   U106 : NAND2_X1 port map( A1 => n242, A2 => n241, ZN => Y(34));
   U107 : AOI22_X1 port map( A1 => A_neg(34), A2 => n154, B1 => A_signal(34), 
                           B2 => n145, ZN => n242);
   U108 : AOI222_X1 port map( A1 => A_shifted(34), A2 => n179, B1 => 
                           zeroSignal(34), B2 => n170, C1 => A_neg_shifted(34),
                           C2 => n163, ZN => n241);
   U109 : NAND2_X1 port map( A1 => n192, A2 => n191, ZN => Y(11));
   U110 : AOI222_X1 port map( A1 => A_shifted(11), A2 => n177, B1 => 
                           zeroSignal(11), B2 => n168, C1 => A_neg_shifted(11),
                           C2 => n165, ZN => n191);
   U111 : NAND2_X1 port map( A1 => n194, A2 => n193, ZN => Y(12));
   U112 : AOI222_X1 port map( A1 => A_shifted(12), A2 => n177, B1 => 
                           zeroSignal(12), B2 => n168, C1 => A_neg_shifted(12),
                           C2 => n165, ZN => n193);
   U113 : NAND2_X1 port map( A1 => n244, A2 => n243, ZN => Y(35));
   U114 : AOI22_X1 port map( A1 => A_neg(35), A2 => n154, B1 => A_signal(35), 
                           B2 => n145, ZN => n244);
   U115 : AOI222_X1 port map( A1 => A_shifted(35), A2 => n179, B1 => 
                           zeroSignal(35), B2 => n170, C1 => A_neg_shifted(35),
                           C2 => n162, ZN => n243);
   U116 : NAND2_X1 port map( A1 => n250, A2 => n249, ZN => Y(38));
   U117 : AOI22_X1 port map( A1 => A_neg(38), A2 => n154, B1 => A_signal(38), 
                           B2 => n145, ZN => n250);
   U118 : AOI222_X1 port map( A1 => A_shifted(38), A2 => n179, B1 => 
                           zeroSignal(38), B2 => n170, C1 => A_neg_shifted(38),
                           C2 => n162, ZN => n249);
   U119 : NAND2_X1 port map( A1 => n246, A2 => n245, ZN => Y(36));
   U120 : AOI22_X1 port map( A1 => A_neg(36), A2 => n154, B1 => A_signal(36), 
                           B2 => n145, ZN => n246);
   U121 : AOI222_X1 port map( A1 => A_shifted(36), A2 => n179, B1 => 
                           zeroSignal(36), B2 => n170, C1 => A_neg_shifted(36),
                           C2 => n162, ZN => n245);
   U122 : AOI222_X1 port map( A1 => A_shifted(13), A2 => n177, B1 => 
                           zeroSignal(13), B2 => n168, C1 => A_neg_shifted(13),
                           C2 => n164, ZN => n195);
   U123 : NAND2_X1 port map( A1 => n252, A2 => n251, ZN => Y(39));
   U124 : AOI222_X1 port map( A1 => A_shifted(39), A2 => n179, B1 => 
                           zeroSignal(39), B2 => n170, C1 => A_neg_shifted(39),
                           C2 => n162, ZN => n251);
   U125 : AOI22_X1 port map( A1 => A_neg(39), A2 => n154, B1 => A_signal(39), 
                           B2 => n145, ZN => n252);
   U126 : NAND2_X1 port map( A1 => n198, A2 => n197, ZN => Y(14));
   U127 : AOI22_X1 port map( A1 => A_neg(14), A2 => n152, B1 => A_signal(14), 
                           B2 => n143, ZN => n198);
   U128 : AOI222_X1 port map( A1 => A_shifted(14), A2 => n177, B1 => 
                           zeroSignal(14), B2 => n168, C1 => A_neg_shifted(14),
                           C2 => n164, ZN => n197);
   U129 : NAND2_X1 port map( A1 => n208, A2 => n207, ZN => Y(19));
   U130 : AOI22_X1 port map( A1 => A_neg(19), A2 => n152, B1 => A_signal(19), 
                           B2 => n143, ZN => n208);
   U131 : AOI222_X1 port map( A1 => A_shifted(19), A2 => n177, B1 => 
                           zeroSignal(19), B2 => n168, C1 => A_neg_shifted(19),
                           C2 => n164, ZN => n207);
   U132 : NAND2_X1 port map( A1 => n256, A2 => n255, ZN => Y(40));
   U133 : AOI222_X1 port map( A1 => A_shifted(40), A2 => n179, B1 => 
                           zeroSignal(40), B2 => n170, C1 => A_neg_shifted(40),
                           C2 => n162, ZN => n255);
   U134 : AOI22_X1 port map( A1 => A_neg(40), A2 => n154, B1 => A_signal(40), 
                           B2 => n145, ZN => n256);
   U135 : NAND2_X1 port map( A1 => n218, A2 => n217, ZN => Y(23));
   U136 : AOI22_X1 port map( A1 => A_neg(23), A2 => n153, B1 => A_signal(23), 
                           B2 => n144, ZN => n218);
   U137 : AOI222_X1 port map( A1 => A_shifted(23), A2 => n178, B1 => 
                           zeroSignal(23), B2 => n169, C1 => A_neg_shifted(23),
                           C2 => n164, ZN => n217);
   U138 : NAND2_X1 port map( A1 => n258, A2 => n257, ZN => Y(41));
   U139 : AOI22_X1 port map( A1 => A_neg(41), A2 => n154, B1 => A_signal(41), 
                           B2 => n145, ZN => n258);
   U140 : AOI222_X1 port map( A1 => A_shifted(41), A2 => n179, B1 => 
                           zeroSignal(41), B2 => n170, C1 => A_neg_shifted(41),
                           C2 => n162, ZN => n257);
   U141 : NAND2_X1 port map( A1 => n300, A2 => n299, ZN => Y(60));
   U142 : AOI222_X1 port map( A1 => A_shifted(60), A2 => n181, B1 => 
                           zeroSignal(60), B2 => n172, C1 => A_neg_shifted(60),
                           C2 => n160, ZN => n299);
   U143 : AOI22_X1 port map( A1 => A_neg(60), A2 => n156, B1 => A_signal(60), 
                           B2 => n147, ZN => n300);
   U144 : NAND2_X1 port map( A1 => n294, A2 => n293, ZN => Y(58));
   U145 : AOI22_X1 port map( A1 => A_neg(58), A2 => n156, B1 => A_signal(58), 
                           B2 => n147, ZN => n294);
   U146 : NAND2_X1 port map( A1 => n296, A2 => n295, ZN => Y(59));
   U147 : AOI222_X1 port map( A1 => A_shifted(59), A2 => n181, B1 => 
                           zeroSignal(59), B2 => n172, C1 => A_neg_shifted(59),
                           C2 => n160, ZN => n295);
   U148 : AOI22_X1 port map( A1 => A_neg(59), A2 => n156, B1 => A_signal(59), 
                           B2 => n147, ZN => n296);
   U149 : NAND2_X1 port map( A1 => n302, A2 => n301, ZN => Y(61));
   U150 : AOI222_X1 port map( A1 => A_shifted(61), A2 => n181, B1 => 
                           zeroSignal(61), B2 => n172, C1 => A_neg_shifted(61),
                           C2 => n160, ZN => n301);
   U151 : AOI22_X1 port map( A1 => A_neg(61), A2 => n156, B1 => A_signal(61), 
                           B2 => n147, ZN => n302);
   U152 : NAND2_X1 port map( A1 => n304, A2 => n303, ZN => Y(62));
   U153 : AOI222_X1 port map( A1 => A_shifted(62), A2 => n181, B1 => 
                           zeroSignal(62), B2 => n172, C1 => A_neg_shifted(62),
                           C2 => n160, ZN => n303);
   U154 : AOI22_X1 port map( A1 => A_neg(62), A2 => n156, B1 => A_signal(62), 
                           B2 => n147, ZN => n304);
   U155 : NAND2_X1 port map( A1 => n266, A2 => n265, ZN => Y(45));
   U156 : AOI222_X1 port map( A1 => A_shifted(45), A2 => n180, B1 => 
                           zeroSignal(45), B2 => n171, C1 => A_neg_shifted(45),
                           C2 => n162, ZN => n265);
   U157 : AOI22_X1 port map( A1 => A_neg(45), A2 => n155, B1 => A_signal(45), 
                           B2 => n146, ZN => n266);
   U158 : NAND2_X1 port map( A1 => n306, A2 => n305, ZN => Y(63));
   U159 : AOI222_X1 port map( A1 => A_shifted(63), A2 => n181, B1 => 
                           zeroSignal(63), B2 => n172, C1 => A_neg_shifted(63),
                           C2 => n160, ZN => n305);
   U160 : AOI22_X1 port map( A1 => A_neg(63), A2 => n156, B1 => A_signal(63), 
                           B2 => n147, ZN => n306);
   U161 : NAND2_X1 port map( A1 => n230, A2 => n229, ZN => Y(29));
   U162 : AOI22_X1 port map( A1 => A_neg(29), A2 => n153, B1 => A_signal(29), 
                           B2 => n144, ZN => n230);
   U163 : AOI222_X1 port map( A1 => A_shifted(29), A2 => n178, B1 => 
                           zeroSignal(29), B2 => n169, C1 => A_neg_shifted(29),
                           C2 => n163, ZN => n229);
   U164 : NAND2_X1 port map( A1 => n282, A2 => n281, ZN => Y(52));
   U165 : NAND2_X1 port map( A1 => n272, A2 => n271, ZN => Y(48));
   U166 : AOI222_X1 port map( A1 => A_shifted(48), A2 => n180, B1 => 
                           zeroSignal(48), B2 => n171, C1 => A_neg_shifted(48),
                           C2 => n161, ZN => n271);
   U167 : NAND2_X1 port map( A1 => n270, A2 => n269, ZN => Y(47));
   U168 : AOI222_X1 port map( A1 => A_shifted(47), A2 => n180, B1 => 
                           zeroSignal(47), B2 => n171, C1 => A_neg_shifted(47),
                           C2 => n161, ZN => n269);
   U169 : AOI22_X1 port map( A1 => A_neg(47), A2 => n155, B1 => A_signal(47), 
                           B2 => n146, ZN => n270);
   U170 : NAND2_X1 port map( A1 => n280, A2 => n279, ZN => Y(51));
   U171 : NAND2_X1 port map( A1 => n278, A2 => n277, ZN => Y(50));
   U172 : AOI222_X1 port map( A1 => A_shifted(50), A2 => n180, B1 => 
                           zeroSignal(50), B2 => n171, C1 => A_neg_shifted(50),
                           C2 => n161, ZN => n277);
   U173 : NAND2_X1 port map( A1 => n274, A2 => n273, ZN => Y(49));
   U174 : AOI22_X1 port map( A1 => A_neg(49), A2 => n155, B1 => A_signal(49), 
                           B2 => n146, ZN => n274);
   U175 : NAND2_X1 port map( A1 => n286, A2 => n285, ZN => Y(54));
   U176 : AOI222_X1 port map( A1 => A_shifted(54), A2 => n181, B1 => 
                           zeroSignal(54), B2 => n172, C1 => A_neg_shifted(54),
                           C2 => n161, ZN => n285);
   U177 : NAND2_X1 port map( A1 => n268, A2 => n267, ZN => Y(46));
   U178 : AOI22_X1 port map( A1 => A_neg(46), A2 => n155, B1 => A_signal(46), 
                           B2 => n146, ZN => n268);
   U179 : AOI222_X1 port map( A1 => A_shifted(46), A2 => n180, B1 => 
                           zeroSignal(46), B2 => n171, C1 => A_neg_shifted(46),
                           C2 => n161, ZN => n267);
   U180 : NAND2_X1 port map( A1 => n284, A2 => n283, ZN => Y(53));
   U181 : AOI22_X1 port map( A1 => A_neg(53), A2 => n156, B1 => A_signal(53), 
                           B2 => n147, ZN => n284);
   U182 : NAND2_X1 port map( A1 => n292, A2 => n291, ZN => Y(57));
   U183 : AOI222_X1 port map( A1 => A_shifted(57), A2 => n181, B1 => 
                           zeroSignal(57), B2 => n172, C1 => A_neg_shifted(57),
                           C2 => n160, ZN => n291);
   U184 : NAND2_X1 port map( A1 => n288, A2 => n287, ZN => Y(55));
   U185 : AOI22_X1 port map( A1 => A_neg(55), A2 => n156, B1 => A_signal(55), 
                           B2 => n147, ZN => n288);
   U186 : NAND2_X1 port map( A1 => n290, A2 => n289, ZN => Y(56));
   U187 : AOI222_X1 port map( A1 => A_shifted(56), A2 => n181, B1 => 
                           zeroSignal(56), B2 => n172, C1 => A_neg_shifted(56),
                           C2 => n161, ZN => n289);
   U188 : AOI22_X1 port map( A1 => A_neg(56), A2 => n156, B1 => A_signal(56), 
                           B2 => n147, ZN => n290);
   U189 : NAND2_X1 port map( A1 => n260, A2 => n259, ZN => Y(42));
   U190 : AOI22_X1 port map( A1 => A_neg(42), A2 => n155, B1 => A_signal(42), 
                           B2 => n146, ZN => n260);
   U191 : AOI222_X1 port map( A1 => A_shifted(42), A2 => n180, B1 => 
                           zeroSignal(42), B2 => n171, C1 => A_neg_shifted(42),
                           C2 => n162, ZN => n259);
   U192 : NAND2_X1 port map( A1 => n262, A2 => n261, ZN => Y(43));
   U193 : AOI222_X1 port map( A1 => A_shifted(43), A2 => n180, B1 => 
                           zeroSignal(43), B2 => n171, C1 => A_neg_shifted(43),
                           C2 => n162, ZN => n261);
   U194 : AOI22_X1 port map( A1 => A_neg(43), A2 => n155, B1 => A_signal(43), 
                           B2 => n146, ZN => n262);
   U195 : NAND2_X1 port map( A1 => n264, A2 => n263, ZN => Y(44));
   U196 : AOI222_X1 port map( A1 => A_shifted(44), A2 => n180, B1 => 
                           zeroSignal(44), B2 => n171, C1 => A_neg_shifted(44),
                           C2 => n162, ZN => n263);
   U197 : AOI22_X1 port map( A1 => A_neg(44), A2 => n155, B1 => A_signal(44), 
                           B2 => n146, ZN => n264);
   U198 : NAND2_X1 port map( A1 => n188, A2 => n187, ZN => Y(0));
   U199 : AOI22_X1 port map( A1 => A_neg(0), A2 => n152, B1 => A_signal(0), B2 
                           => n143, ZN => n188);
   U200 : AOI222_X1 port map( A1 => A_shifted(0), A2 => n177, B1 => 
                           zeroSignal(0), B2 => n168, C1 => A_neg_shifted(0), 
                           C2 => n165, ZN => n187);
   U201 : NAND2_X1 port map( A1 => n210, A2 => n209, ZN => Y(1));
   U202 : AOI22_X1 port map( A1 => A_neg(1), A2 => n152, B1 => A_signal(1), B2 
                           => n143, ZN => n210);
   U203 : AOI222_X1 port map( A1 => A_shifted(1), A2 => n177, B1 => 
                           zeroSignal(1), B2 => n168, C1 => A_neg_shifted(1), 
                           C2 => n164, ZN => n209);
   U204 : NAND2_X1 port map( A1 => n232, A2 => n231, ZN => Y(2));
   U205 : AOI22_X1 port map( A1 => A_neg(2), A2 => n153, B1 => A_signal(2), B2 
                           => n144, ZN => n232);
   U206 : AOI222_X1 port map( A1 => A_shifted(2), A2 => n178, B1 => 
                           zeroSignal(2), B2 => n169, C1 => A_neg_shifted(2), 
                           C2 => n163, ZN => n231);
   U207 : NAND2_X1 port map( A1 => n254, A2 => n253, ZN => Y(3));
   U208 : AOI22_X1 port map( A1 => A_neg(3), A2 => n154, B1 => A_signal(3), B2 
                           => n145, ZN => n254);
   U209 : AOI222_X1 port map( A1 => A_shifted(3), A2 => n179, B1 => 
                           zeroSignal(3), B2 => n170, C1 => A_neg_shifted(3), 
                           C2 => n162, ZN => n253);
   U210 : AOI22_X1 port map( A1 => A_neg(12), A2 => n152, B1 => A_signal(12), 
                           B2 => n143, ZN => n194);
   U211 : AOI222_X1 port map( A1 => A_shifted(55), A2 => n181, B1 => 
                           zeroSignal(55), B2 => n172, C1 => A_neg_shifted(55),
                           C2 => n161, ZN => n287);
   U212 : AOI22_X1 port map( A1 => A_neg(54), A2 => n156, B1 => A_signal(54), 
                           B2 => n147, ZN => n286);
   U213 : AOI222_X1 port map( A1 => A_shifted(58), A2 => n181, B1 => 
                           zeroSignal(58), B2 => n172, C1 => A_neg_shifted(58),
                           C2 => n160, ZN => n293);
   U214 : AOI22_X1 port map( A1 => A_neg(57), A2 => n156, B1 => A_signal(57), 
                           B2 => n147, ZN => n292);
   U215 : AOI222_X1 port map( A1 => A_shifted(53), A2 => n181, B1 => 
                           zeroSignal(53), B2 => n172, C1 => A_neg_shifted(53),
                           C2 => n161, ZN => n283);
   U216 : AOI22_X1 port map( A1 => A_neg(52), A2 => n155, B1 => A_signal(52), 
                           B2 => n146, ZN => n282);
   U217 : AOI222_X1 port map( A1 => A_shifted(51), A2 => n180, B1 => 
                           zeroSignal(51), B2 => n171, C1 => A_neg_shifted(51),
                           C2 => n161, ZN => n279);
   U218 : AOI22_X1 port map( A1 => A_neg(50), A2 => n155, B1 => A_signal(50), 
                           B2 => n146, ZN => n278);
   U219 : AOI22_X1 port map( A1 => A_neg(11), A2 => n152, B1 => A_signal(11), 
                           B2 => n143, ZN => n192);
   U220 : AOI222_X1 port map( A1 => A_shifted(52), A2 => n180, B1 => 
                           zeroSignal(52), B2 => n171, C1 => A_neg_shifted(52),
                           C2 => n161, ZN => n281);
   U221 : AOI22_X1 port map( A1 => A_neg(51), A2 => n155, B1 => A_signal(51), 
                           B2 => n146, ZN => n280);
   U222 : AOI222_X1 port map( A1 => A_shifted(49), A2 => n180, B1 => 
                           zeroSignal(49), B2 => n171, C1 => A_neg_shifted(49),
                           C2 => n161, ZN => n273);
   U223 : AOI22_X1 port map( A1 => A_neg(48), A2 => n155, B1 => A_signal(48), 
                           B2 => n146, ZN => n272);
   U224 : NAND2_X1 port map( A1 => n276, A2 => n275, ZN => Y(4));
   U225 : AOI22_X1 port map( A1 => A_neg(4), A2 => n155, B1 => A_signal(4), B2 
                           => n146, ZN => n276);
   U226 : NOR3_X1 port map( A1 => n318, A2 => Sel(2), A3 => n319, ZN => n315);
   U227 : NOR3_X1 port map( A1 => Sel(1), A2 => Sel(2), A3 => n318, ZN => n313)
                           ;
   U228 : AOI21_X1 port map( B1 => n318, B2 => n319, A => Sel(2), ZN => n186);
   U229 : NAND2_X1 port map( A1 => n298, A2 => n297, ZN => Y(5));
   U230 : AOI22_X1 port map( A1 => A_neg(5), A2 => n156, B1 => A_signal(5), B2 
                           => n147, ZN => n298);
   U231 : AOI222_X1 port map( A1 => A_shifted(5), A2 => n181, B1 => 
                           zeroSignal(5), B2 => n172, C1 => A_neg_shifted(5), 
                           C2 => n160, ZN => n297);
   U232 : INV_X1 port map( A => Sel(1), ZN => n319);
   U233 : AOI22_X1 port map( A1 => A_neg(13), A2 => n152, B1 => A_signal(13), 
                           B2 => n143, ZN => n196);
   U234 : NAND2_X1 port map( A1 => n312, A2 => n311, ZN => Y(8));
   U235 : NAND2_X1 port map( A1 => n310, A2 => n309, ZN => Y(7));
   U236 : AOI22_X1 port map( A1 => A_neg(10), A2 => n152, B1 => A_signal(10), 
                           B2 => n143, ZN => n190);
   U237 : AOI22_X1 port map( A1 => A_neg(7), A2 => n157, B1 => A_signal(7), B2 
                           => n148, ZN => n310);
   U238 : AOI22_X1 port map( A1 => A_neg(28), A2 => n153, B1 => A_signal(28), 
                           B2 => n144, ZN => n228);
   U239 : AOI22_X1 port map( A1 => A_neg(22), A2 => n153, B1 => A_signal(22), 
                           B2 => n144, ZN => n216);
   U240 : AOI22_X1 port map( A1 => A_neg(18), A2 => n152, B1 => A_signal(18), 
                           B2 => n143, ZN => n206);
   U241 : AOI22_X1 port map( A1 => A_neg(6), A2 => n157, B1 => A_signal(6), B2 
                           => n148, ZN => n308);
   U242 : AOI22_X1 port map( A1 => A_neg(9), A2 => n157, B1 => A_signal(9), B2 
                           => n148, ZN => n317);
   U243 : AOI22_X1 port map( A1 => A_neg(8), A2 => n157, B1 => A_signal(8), B2 
                           => n148, ZN => n312);

end SYN_BEHAVIORAL_2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity MUX51_MuxNbit64_29 is

   port( zeroSignal, A_signal, A_neg, A_shifted, A_neg_shifted : in 
         std_logic_vector (63 downto 0);  Sel : in std_logic_vector (2 downto 
         0);  Y : out std_logic_vector (63 downto 0));

end MUX51_MuxNbit64_29;

architecture SYN_BEHAVIORAL_2 of MUX51_MuxNbit64_29 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, 
      n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, 
      n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, 
      n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, 
      n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, 
      n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, 
      n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, 
      n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, 
      n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, 
      n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, 
      n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, 
      n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, 
      n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, 
      n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, 
      n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319 : 
      std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n264, A2 => n263, ZN => Y(44));
   U2 : CLKBUF_X1 port map( A => n167, Z => n161);
   U3 : CLKBUF_X1 port map( A => n141, Z => n166);
   U4 : BUF_X1 port map( A => n141, Z => n167);
   U5 : BUF_X1 port map( A => n142, Z => n149);
   U6 : BUF_X1 port map( A => n185, Z => n183);
   U7 : BUF_X1 port map( A => n159, Z => n157);
   U8 : BUF_X1 port map( A => n142, Z => n150);
   U9 : BUF_X1 port map( A => n185, Z => n184);
   U10 : BUF_X1 port map( A => n159, Z => n158);
   U11 : BUF_X1 port map( A => n176, Z => n175);
   U12 : BUF_X1 port map( A => n176, Z => n174);
   U13 : AND3_X1 port map( A1 => n318, A2 => n319, A3 => Sel(2), ZN => n141);
   U14 : NOR3_X1 port map( A1 => Sel(1), A2 => Sel(2), A3 => n318, ZN => n142);
   U15 : BUF_X1 port map( A => n315, Z => n185);
   U16 : BUF_X1 port map( A => n313, Z => n159);
   U17 : BUF_X1 port map( A => n157, Z => n156);
   U18 : BUF_X1 port map( A => n183, Z => n182);
   U19 : BUF_X1 port map( A => n149, Z => n148);
   U20 : BUF_X1 port map( A => n167, Z => n160);
   U21 : BUF_X1 port map( A => n184, Z => n177);
   U22 : BUF_X1 port map( A => n158, Z => n151);
   U23 : BUF_X1 port map( A => n150, Z => n143);
   U24 : BUF_X1 port map( A => n166, Z => n165);
   U25 : BUF_X1 port map( A => n166, Z => n164);
   U26 : BUF_X1 port map( A => n184, Z => n178);
   U27 : BUF_X1 port map( A => n158, Z => n152);
   U28 : BUF_X1 port map( A => n150, Z => n144);
   U29 : BUF_X1 port map( A => n166, Z => n163);
   U30 : BUF_X1 port map( A => n184, Z => n179);
   U31 : BUF_X1 port map( A => n158, Z => n153);
   U32 : BUF_X1 port map( A => n150, Z => n145);
   U33 : BUF_X1 port map( A => n167, Z => n162);
   U34 : BUF_X1 port map( A => n183, Z => n180);
   U35 : BUF_X1 port map( A => n157, Z => n154);
   U36 : BUF_X1 port map( A => n149, Z => n146);
   U37 : BUF_X1 port map( A => n183, Z => n181);
   U38 : BUF_X1 port map( A => n157, Z => n155);
   U39 : BUF_X1 port map( A => n149, Z => n147);
   U40 : BUF_X1 port map( A => n175, Z => n168);
   U41 : BUF_X1 port map( A => n175, Z => n169);
   U42 : BUF_X1 port map( A => n175, Z => n170);
   U43 : BUF_X1 port map( A => n174, Z => n171);
   U44 : BUF_X1 port map( A => n174, Z => n172);
   U45 : BUF_X1 port map( A => n174, Z => n173);
   U46 : INV_X1 port map( A => Sel(1), ZN => n319);
   U47 : NOR3_X1 port map( A1 => Sel(0), A2 => Sel(2), A3 => n319, ZN => n313);
   U48 : NOR3_X1 port map( A1 => n318, A2 => Sel(2), A3 => n319, ZN => n315);
   U49 : INV_X1 port map( A => Sel(0), ZN => n318);
   U50 : BUF_X1 port map( A => n314, Z => n176);
   U51 : NOR2_X1 port map( A1 => n165, A2 => n186, ZN => n314);
   U52 : AOI21_X1 port map( B1 => n318, B2 => n319, A => Sel(2), ZN => n186);
   U53 : AOI22_X1 port map( A1 => A_neg(7), A2 => n156, B1 => A_signal(7), B2 
                           => n148, ZN => n310);
   U54 : AOI222_X1 port map( A1 => A_shifted(6), A2 => n182, B1 => 
                           zeroSignal(6), B2 => n173, C1 => A_neg_shifted(6), 
                           C2 => n160, ZN => n307);
   U55 : NAND2_X1 port map( A1 => n312, A2 => n311, ZN => Y(8));
   U56 : AOI22_X1 port map( A1 => A_neg(8), A2 => n156, B1 => A_signal(8), B2 
                           => n148, ZN => n312);
   U57 : AOI222_X1 port map( A1 => A_shifted(8), A2 => n182, B1 => 
                           zeroSignal(8), B2 => n173, C1 => A_neg_shifted(8), 
                           C2 => n160, ZN => n311);
   U58 : NAND2_X1 port map( A1 => n317, A2 => n316, ZN => Y(9));
   U59 : AOI22_X1 port map( A1 => A_neg(9), A2 => n156, B1 => A_signal(9), B2 
                           => n148, ZN => n317);
   U60 : AOI222_X1 port map( A1 => A_shifted(9), A2 => n182, B1 => 
                           zeroSignal(9), B2 => n173, C1 => A_neg_shifted(9), 
                           C2 => n160, ZN => n316);
   U61 : NAND2_X1 port map( A1 => n190, A2 => n189, ZN => Y(10));
   U62 : AOI22_X1 port map( A1 => A_neg(10), A2 => n151, B1 => A_signal(10), B2
                           => n143, ZN => n190);
   U63 : AOI222_X1 port map( A1 => A_shifted(10), A2 => n177, B1 => 
                           zeroSignal(10), B2 => n168, C1 => A_neg_shifted(10),
                           C2 => n165, ZN => n189);
   U64 : NAND2_X1 port map( A1 => n192, A2 => n191, ZN => Y(11));
   U65 : AOI22_X1 port map( A1 => A_neg(11), A2 => n151, B1 => A_signal(11), B2
                           => n143, ZN => n192);
   U66 : AOI222_X1 port map( A1 => A_shifted(11), A2 => n177, B1 => 
                           zeroSignal(11), B2 => n168, C1 => A_neg_shifted(11),
                           C2 => n165, ZN => n191);
   U67 : NAND2_X1 port map( A1 => n194, A2 => n193, ZN => Y(12));
   U68 : AOI22_X1 port map( A1 => A_neg(12), A2 => n151, B1 => A_signal(12), B2
                           => n143, ZN => n194);
   U69 : AOI222_X1 port map( A1 => A_shifted(12), A2 => n177, B1 => 
                           zeroSignal(12), B2 => n168, C1 => A_neg_shifted(12),
                           C2 => n165, ZN => n193);
   U70 : NAND2_X1 port map( A1 => n196, A2 => n195, ZN => Y(13));
   U71 : AOI22_X1 port map( A1 => A_neg(13), A2 => n151, B1 => A_signal(13), B2
                           => n143, ZN => n196);
   U72 : AOI222_X1 port map( A1 => A_shifted(13), A2 => n177, B1 => 
                           zeroSignal(13), B2 => n168, C1 => A_neg_shifted(13),
                           C2 => n164, ZN => n195);
   U73 : NAND2_X1 port map( A1 => n206, A2 => n205, ZN => Y(18));
   U74 : AOI222_X1 port map( A1 => A_shifted(18), A2 => n177, B1 => 
                           zeroSignal(18), B2 => n168, C1 => A_neg_shifted(18),
                           C2 => n164, ZN => n205);
   U75 : AOI22_X1 port map( A1 => A_neg(18), A2 => n151, B1 => A_signal(18), B2
                           => n143, ZN => n206);
   U76 : NAND2_X1 port map( A1 => n204, A2 => n203, ZN => Y(17));
   U77 : AOI222_X1 port map( A1 => A_shifted(17), A2 => n177, B1 => 
                           zeroSignal(17), B2 => n168, C1 => A_neg_shifted(17),
                           C2 => n164, ZN => n203);
   U78 : AOI22_X1 port map( A1 => A_neg(17), A2 => n151, B1 => A_signal(17), B2
                           => n143, ZN => n204);
   U79 : NAND2_X1 port map( A1 => n208, A2 => n207, ZN => Y(19));
   U80 : AOI222_X1 port map( A1 => A_shifted(19), A2 => n177, B1 => 
                           zeroSignal(19), B2 => n168, C1 => A_neg_shifted(19),
                           C2 => n164, ZN => n207);
   U81 : AOI22_X1 port map( A1 => A_neg(19), A2 => n151, B1 => A_signal(19), B2
                           => n143, ZN => n208);
   U82 : NAND2_X1 port map( A1 => n202, A2 => n201, ZN => Y(16));
   U83 : AOI222_X1 port map( A1 => A_shifted(16), A2 => n177, B1 => 
                           zeroSignal(16), B2 => n168, C1 => A_neg_shifted(16),
                           C2 => n164, ZN => n201);
   U84 : AOI22_X1 port map( A1 => A_neg(16), A2 => n151, B1 => A_signal(16), B2
                           => n143, ZN => n202);
   U85 : NAND2_X1 port map( A1 => n216, A2 => n215, ZN => Y(22));
   U86 : AOI222_X1 port map( A1 => A_shifted(22), A2 => n178, B1 => 
                           zeroSignal(22), B2 => n169, C1 => A_neg_shifted(22),
                           C2 => n164, ZN => n215);
   U87 : AOI22_X1 port map( A1 => A_neg(22), A2 => n152, B1 => A_signal(22), B2
                           => n144, ZN => n216);
   U88 : NAND2_X1 port map( A1 => n214, A2 => n213, ZN => Y(21));
   U89 : AOI222_X1 port map( A1 => A_shifted(21), A2 => n178, B1 => 
                           zeroSignal(21), B2 => n169, C1 => A_neg_shifted(21),
                           C2 => n164, ZN => n213);
   U90 : AOI22_X1 port map( A1 => A_neg(21), A2 => n152, B1 => A_signal(21), B2
                           => n144, ZN => n214);
   U91 : NAND2_X1 port map( A1 => n218, A2 => n217, ZN => Y(23));
   U92 : AOI222_X1 port map( A1 => A_shifted(23), A2 => n178, B1 => 
                           zeroSignal(23), B2 => n169, C1 => A_neg_shifted(23),
                           C2 => n164, ZN => n217);
   U93 : AOI22_X1 port map( A1 => A_neg(23), A2 => n152, B1 => A_signal(23), B2
                           => n144, ZN => n218);
   U94 : NAND2_X1 port map( A1 => n226, A2 => n225, ZN => Y(27));
   U95 : AOI222_X1 port map( A1 => A_shifted(27), A2 => n178, B1 => 
                           zeroSignal(27), B2 => n169, C1 => A_neg_shifted(27),
                           C2 => n163, ZN => n225);
   U96 : AOI22_X1 port map( A1 => A_neg(27), A2 => n152, B1 => A_signal(27), B2
                           => n144, ZN => n226);
   U97 : NAND2_X1 port map( A1 => n212, A2 => n211, ZN => Y(20));
   U98 : AOI22_X1 port map( A1 => A_neg(20), A2 => n152, B1 => A_signal(20), B2
                           => n144, ZN => n212);
   U99 : AOI222_X1 port map( A1 => A_shifted(20), A2 => n178, B1 => 
                           zeroSignal(20), B2 => n169, C1 => A_neg_shifted(20),
                           C2 => n164, ZN => n211);
   U100 : NAND2_X1 port map( A1 => n222, A2 => n221, ZN => Y(25));
   U101 : AOI222_X1 port map( A1 => A_shifted(25), A2 => n178, B1 => 
                           zeroSignal(25), B2 => n169, C1 => A_neg_shifted(25),
                           C2 => n163, ZN => n221);
   U102 : AOI22_X1 port map( A1 => A_neg(25), A2 => n152, B1 => A_signal(25), 
                           B2 => n144, ZN => n222);
   U103 : NAND2_X1 port map( A1 => n224, A2 => n223, ZN => Y(26));
   U104 : AOI222_X1 port map( A1 => A_shifted(26), A2 => n178, B1 => 
                           zeroSignal(26), B2 => n169, C1 => A_neg_shifted(26),
                           C2 => n163, ZN => n223);
   U105 : AOI22_X1 port map( A1 => A_neg(26), A2 => n152, B1 => A_signal(26), 
                           B2 => n144, ZN => n224);
   U106 : NAND2_X1 port map( A1 => n228, A2 => n227, ZN => Y(28));
   U107 : AOI222_X1 port map( A1 => A_shifted(28), A2 => n178, B1 => 
                           zeroSignal(28), B2 => n169, C1 => A_neg_shifted(28),
                           C2 => n163, ZN => n227);
   U108 : AOI22_X1 port map( A1 => A_neg(28), A2 => n152, B1 => A_signal(28), 
                           B2 => n144, ZN => n228);
   U109 : NAND2_X1 port map( A1 => n220, A2 => n219, ZN => Y(24));
   U110 : AOI22_X1 port map( A1 => A_neg(24), A2 => n152, B1 => A_signal(24), 
                           B2 => n144, ZN => n220);
   U111 : AOI222_X1 port map( A1 => A_shifted(24), A2 => n178, B1 => 
                           zeroSignal(24), B2 => n169, C1 => A_neg_shifted(24),
                           C2 => n163, ZN => n219);
   U112 : NAND2_X1 port map( A1 => n198, A2 => n197, ZN => Y(14));
   U113 : AOI22_X1 port map( A1 => A_neg(14), A2 => n151, B1 => A_signal(14), 
                           B2 => n143, ZN => n198);
   U114 : AOI222_X1 port map( A1 => A_shifted(14), A2 => n177, B1 => 
                           zeroSignal(14), B2 => n168, C1 => A_neg_shifted(14),
                           C2 => n164, ZN => n197);
   U115 : NAND2_X1 port map( A1 => n230, A2 => n229, ZN => Y(29));
   U116 : AOI222_X1 port map( A1 => A_shifted(29), A2 => n178, B1 => 
                           zeroSignal(29), B2 => n169, C1 => A_neg_shifted(29),
                           C2 => n163, ZN => n229);
   U117 : AOI22_X1 port map( A1 => A_neg(29), A2 => n152, B1 => A_signal(29), 
                           B2 => n144, ZN => n230);
   U118 : NAND2_X1 port map( A1 => n236, A2 => n235, ZN => Y(31));
   U119 : AOI222_X1 port map( A1 => A_shifted(31), A2 => n179, B1 => 
                           zeroSignal(31), B2 => n170, C1 => A_neg_shifted(31),
                           C2 => n163, ZN => n235);
   U120 : AOI22_X1 port map( A1 => A_neg(31), A2 => n153, B1 => A_signal(31), 
                           B2 => n145, ZN => n236);
   U121 : NAND2_X1 port map( A1 => n240, A2 => n239, ZN => Y(33));
   U122 : AOI222_X1 port map( A1 => A_shifted(33), A2 => n179, B1 => 
                           zeroSignal(33), B2 => n170, C1 => A_neg_shifted(33),
                           C2 => n163, ZN => n239);
   U123 : AOI22_X1 port map( A1 => A_neg(33), A2 => n153, B1 => A_signal(33), 
                           B2 => n145, ZN => n240);
   U124 : NAND2_X1 port map( A1 => n238, A2 => n237, ZN => Y(32));
   U125 : AOI222_X1 port map( A1 => A_shifted(32), A2 => n179, B1 => 
                           zeroSignal(32), B2 => n170, C1 => A_neg_shifted(32),
                           C2 => n163, ZN => n237);
   U126 : AOI22_X1 port map( A1 => A_neg(32), A2 => n153, B1 => A_signal(32), 
                           B2 => n145, ZN => n238);
   U127 : NAND2_X1 port map( A1 => n252, A2 => n251, ZN => Y(39));
   U128 : AOI222_X1 port map( A1 => A_shifted(39), A2 => n179, B1 => 
                           zeroSignal(39), B2 => n170, C1 => A_neg_shifted(39),
                           C2 => n162, ZN => n251);
   U129 : AOI22_X1 port map( A1 => A_neg(39), A2 => n153, B1 => A_signal(39), 
                           B2 => n145, ZN => n252);
   U130 : NAND2_X1 port map( A1 => n244, A2 => n243, ZN => Y(35));
   U131 : AOI222_X1 port map( A1 => A_shifted(35), A2 => n179, B1 => 
                           zeroSignal(35), B2 => n170, C1 => A_neg_shifted(35),
                           C2 => n162, ZN => n243);
   U132 : AOI22_X1 port map( A1 => A_neg(35), A2 => n153, B1 => A_signal(35), 
                           B2 => n145, ZN => n244);
   U133 : NAND2_X1 port map( A1 => n248, A2 => n247, ZN => Y(37));
   U134 : AOI222_X1 port map( A1 => A_shifted(37), A2 => n179, B1 => 
                           zeroSignal(37), B2 => n170, C1 => A_neg_shifted(37),
                           C2 => n162, ZN => n247);
   U135 : AOI22_X1 port map( A1 => A_neg(37), A2 => n153, B1 => A_signal(37), 
                           B2 => n145, ZN => n248);
   U136 : NAND2_X1 port map( A1 => n234, A2 => n233, ZN => Y(30));
   U137 : AOI22_X1 port map( A1 => A_neg(30), A2 => n152, B1 => A_signal(30), 
                           B2 => n144, ZN => n234);
   U138 : AOI222_X1 port map( A1 => A_shifted(30), A2 => n178, B1 => 
                           zeroSignal(30), B2 => n169, C1 => A_neg_shifted(30),
                           C2 => n163, ZN => n233);
   U139 : NAND2_X1 port map( A1 => n242, A2 => n241, ZN => Y(34));
   U140 : AOI222_X1 port map( A1 => A_shifted(34), A2 => n179, B1 => 
                           zeroSignal(34), B2 => n170, C1 => A_neg_shifted(34),
                           C2 => n163, ZN => n241);
   U141 : AOI22_X1 port map( A1 => A_neg(34), A2 => n153, B1 => A_signal(34), 
                           B2 => n145, ZN => n242);
   U142 : NAND2_X1 port map( A1 => n246, A2 => n245, ZN => Y(36));
   U143 : AOI222_X1 port map( A1 => A_shifted(36), A2 => n179, B1 => 
                           zeroSignal(36), B2 => n170, C1 => A_neg_shifted(36),
                           C2 => n162, ZN => n245);
   U144 : AOI22_X1 port map( A1 => A_neg(36), A2 => n153, B1 => A_signal(36), 
                           B2 => n145, ZN => n246);
   U145 : NAND2_X1 port map( A1 => n200, A2 => n199, ZN => Y(15));
   U146 : AOI22_X1 port map( A1 => A_neg(15), A2 => n151, B1 => A_signal(15), 
                           B2 => n143, ZN => n200);
   U147 : AOI222_X1 port map( A1 => A_shifted(15), A2 => n177, B1 => 
                           zeroSignal(15), B2 => n168, C1 => A_neg_shifted(15),
                           C2 => n164, ZN => n199);
   U148 : NAND2_X1 port map( A1 => n250, A2 => n249, ZN => Y(38));
   U149 : AOI222_X1 port map( A1 => A_shifted(38), A2 => n179, B1 => 
                           zeroSignal(38), B2 => n170, C1 => A_neg_shifted(38),
                           C2 => n162, ZN => n249);
   U150 : AOI22_X1 port map( A1 => A_neg(38), A2 => n153, B1 => A_signal(38), 
                           B2 => n145, ZN => n250);
   U151 : NAND2_X1 port map( A1 => n256, A2 => n255, ZN => Y(40));
   U152 : AOI22_X1 port map( A1 => A_neg(40), A2 => n153, B1 => A_signal(40), 
                           B2 => n145, ZN => n256);
   U153 : AOI222_X1 port map( A1 => A_shifted(40), A2 => n179, B1 => 
                           zeroSignal(40), B2 => n170, C1 => A_neg_shifted(40),
                           C2 => n162, ZN => n255);
   U154 : NAND2_X1 port map( A1 => n258, A2 => n257, ZN => Y(41));
   U155 : AOI222_X1 port map( A1 => A_shifted(41), A2 => n179, B1 => 
                           zeroSignal(41), B2 => n170, C1 => A_neg_shifted(41),
                           C2 => n162, ZN => n257);
   U156 : AOI22_X1 port map( A1 => A_neg(41), A2 => n153, B1 => A_signal(41), 
                           B2 => n145, ZN => n258);
   U157 : NAND2_X1 port map( A1 => n270, A2 => n269, ZN => Y(47));
   U158 : AOI22_X1 port map( A1 => A_neg(47), A2 => n154, B1 => A_signal(47), 
                           B2 => n146, ZN => n270);
   U159 : AOI222_X1 port map( A1 => A_shifted(47), A2 => n180, B1 => 
                           zeroSignal(47), B2 => n171, C1 => A_neg_shifted(47),
                           C2 => n161, ZN => n269);
   U160 : NAND2_X1 port map( A1 => n260, A2 => n259, ZN => Y(42));
   U161 : AOI222_X1 port map( A1 => A_shifted(42), A2 => n180, B1 => 
                           zeroSignal(42), B2 => n171, C1 => A_neg_shifted(42),
                           C2 => n162, ZN => n259);
   U162 : AOI22_X1 port map( A1 => A_neg(42), A2 => n154, B1 => A_signal(42), 
                           B2 => n146, ZN => n260);
   U163 : NAND2_X1 port map( A1 => n262, A2 => n261, ZN => Y(43));
   U164 : AOI22_X1 port map( A1 => A_neg(43), A2 => n154, B1 => A_signal(43), 
                           B2 => n146, ZN => n262);
   U165 : AOI222_X1 port map( A1 => A_shifted(43), A2 => n180, B1 => 
                           zeroSignal(43), B2 => n171, C1 => A_neg_shifted(43),
                           C2 => n162, ZN => n261);
   U166 : NAND2_X1 port map( A1 => n300, A2 => n299, ZN => Y(60));
   U167 : AOI22_X1 port map( A1 => A_neg(60), A2 => n155, B1 => A_signal(60), 
                           B2 => n147, ZN => n300);
   U168 : NAND2_X1 port map( A1 => n304, A2 => n303, ZN => Y(62));
   U169 : AOI222_X1 port map( A1 => A_shifted(62), A2 => n181, B1 => 
                           zeroSignal(62), B2 => n172, C1 => A_neg_shifted(62),
                           C2 => n160, ZN => n303);
   U170 : AOI22_X1 port map( A1 => A_neg(62), A2 => n155, B1 => A_signal(62), 
                           B2 => n147, ZN => n304);
   U171 : NAND2_X1 port map( A1 => n302, A2 => n301, ZN => Y(61));
   U172 : AOI222_X1 port map( A1 => A_shifted(61), A2 => n181, B1 => 
                           zeroSignal(61), B2 => n172, C1 => A_neg_shifted(61),
                           C2 => n160, ZN => n301);
   U173 : AOI22_X1 port map( A1 => A_neg(61), A2 => n155, B1 => A_signal(61), 
                           B2 => n147, ZN => n302);
   U174 : NAND2_X1 port map( A1 => n306, A2 => n305, ZN => Y(63));
   U175 : AOI222_X1 port map( A1 => A_shifted(63), A2 => n181, B1 => 
                           zeroSignal(63), B2 => n172, C1 => A_neg_shifted(63),
                           C2 => n160, ZN => n305);
   U176 : AOI22_X1 port map( A1 => A_neg(63), A2 => n155, B1 => A_signal(63), 
                           B2 => n147, ZN => n306);
   U177 : NAND2_X1 port map( A1 => n284, A2 => n283, ZN => Y(53));
   U178 : NAND2_X1 port map( A1 => n274, A2 => n273, ZN => Y(49));
   U179 : AOI222_X1 port map( A1 => A_shifted(49), A2 => n180, B1 => 
                           zeroSignal(49), B2 => n171, C1 => A_neg_shifted(49),
                           C2 => n161, ZN => n273);
   U180 : AOI22_X1 port map( A1 => A_neg(49), A2 => n154, B1 => A_signal(49), 
                           B2 => n146, ZN => n274);
   U181 : NAND2_X1 port map( A1 => n282, A2 => n281, ZN => Y(52));
   U182 : AOI222_X1 port map( A1 => A_shifted(52), A2 => n180, B1 => 
                           zeroSignal(52), B2 => n171, C1 => A_neg_shifted(52),
                           C2 => n161, ZN => n281);
   U183 : NAND2_X1 port map( A1 => n278, A2 => n277, ZN => Y(50));
   U184 : AOI222_X1 port map( A1 => A_shifted(50), A2 => n180, B1 => 
                           zeroSignal(50), B2 => n171, C1 => A_neg_shifted(50),
                           C2 => n161, ZN => n277);
   U185 : NAND2_X1 port map( A1 => n296, A2 => n295, ZN => Y(59));
   U186 : AOI222_X1 port map( A1 => A_shifted(59), A2 => n181, B1 => 
                           zeroSignal(59), B2 => n172, C1 => A_neg_shifted(59),
                           C2 => n160, ZN => n295);
   U187 : NAND2_X1 port map( A1 => n286, A2 => n285, ZN => Y(54));
   U188 : NAND2_X1 port map( A1 => n290, A2 => n289, ZN => Y(56));
   U189 : AOI222_X1 port map( A1 => A_shifted(56), A2 => n181, B1 => 
                           zeroSignal(56), B2 => n172, C1 => A_neg_shifted(56),
                           C2 => n161, ZN => n289);
   U190 : NAND2_X1 port map( A1 => n280, A2 => n279, ZN => Y(51));
   U191 : AOI22_X1 port map( A1 => A_neg(51), A2 => n154, B1 => A_signal(51), 
                           B2 => n146, ZN => n280);
   U192 : NAND2_X1 port map( A1 => n272, A2 => n271, ZN => Y(48));
   U193 : AOI22_X1 port map( A1 => A_neg(48), A2 => n154, B1 => A_signal(48), 
                           B2 => n146, ZN => n272);
   U194 : AOI222_X1 port map( A1 => A_shifted(48), A2 => n180, B1 => 
                           zeroSignal(48), B2 => n171, C1 => A_neg_shifted(48),
                           C2 => n161, ZN => n271);
   U195 : NAND2_X1 port map( A1 => n294, A2 => n293, ZN => Y(58));
   U196 : AOI222_X1 port map( A1 => A_shifted(58), A2 => n181, B1 => 
                           zeroSignal(58), B2 => n172, C1 => A_neg_shifted(58),
                           C2 => n160, ZN => n293);
   U197 : AOI22_X1 port map( A1 => A_neg(58), A2 => n155, B1 => A_signal(58), 
                           B2 => n147, ZN => n294);
   U198 : NAND2_X1 port map( A1 => n292, A2 => n291, ZN => Y(57));
   U199 : AOI22_X1 port map( A1 => A_neg(57), A2 => n155, B1 => A_signal(57), 
                           B2 => n147, ZN => n292);
   U200 : NAND2_X1 port map( A1 => n288, A2 => n287, ZN => Y(55));
   U201 : AOI22_X1 port map( A1 => A_neg(55), A2 => n155, B1 => A_signal(55), 
                           B2 => n147, ZN => n288);
   U202 : AOI22_X1 port map( A1 => A_neg(44), A2 => n154, B1 => A_signal(44), 
                           B2 => n146, ZN => n264);
   U203 : AOI222_X1 port map( A1 => A_shifted(44), A2 => n180, B1 => 
                           zeroSignal(44), B2 => n171, C1 => A_neg_shifted(44),
                           C2 => n162, ZN => n263);
   U204 : NAND2_X1 port map( A1 => n266, A2 => n265, ZN => Y(45));
   U205 : AOI222_X1 port map( A1 => A_shifted(45), A2 => n180, B1 => 
                           zeroSignal(45), B2 => n171, C1 => A_neg_shifted(45),
                           C2 => n162, ZN => n265);
   U206 : AOI22_X1 port map( A1 => A_neg(45), A2 => n154, B1 => A_signal(45), 
                           B2 => n146, ZN => n266);
   U207 : NAND2_X1 port map( A1 => n268, A2 => n267, ZN => Y(46));
   U208 : AOI222_X1 port map( A1 => A_shifted(46), A2 => n180, B1 => 
                           zeroSignal(46), B2 => n171, C1 => A_neg_shifted(46),
                           C2 => n161, ZN => n267);
   U209 : AOI22_X1 port map( A1 => A_neg(46), A2 => n154, B1 => A_signal(46), 
                           B2 => n146, ZN => n268);
   U210 : NAND2_X1 port map( A1 => n188, A2 => n187, ZN => Y(0));
   U211 : AOI22_X1 port map( A1 => A_neg(0), A2 => n151, B1 => A_signal(0), B2 
                           => n143, ZN => n188);
   U212 : AOI222_X1 port map( A1 => A_shifted(0), A2 => n177, B1 => 
                           zeroSignal(0), B2 => n168, C1 => A_neg_shifted(0), 
                           C2 => n165, ZN => n187);
   U213 : NAND2_X1 port map( A1 => n210, A2 => n209, ZN => Y(1));
   U214 : AOI22_X1 port map( A1 => A_neg(1), A2 => n151, B1 => A_signal(1), B2 
                           => n143, ZN => n210);
   U215 : AOI222_X1 port map( A1 => A_shifted(1), A2 => n177, B1 => 
                           zeroSignal(1), B2 => n168, C1 => A_neg_shifted(1), 
                           C2 => n164, ZN => n209);
   U216 : NAND2_X1 port map( A1 => n232, A2 => n231, ZN => Y(2));
   U217 : AOI22_X1 port map( A1 => A_neg(2), A2 => n152, B1 => A_signal(2), B2 
                           => n144, ZN => n232);
   U218 : AOI222_X1 port map( A1 => A_shifted(2), A2 => n178, B1 => 
                           zeroSignal(2), B2 => n169, C1 => A_neg_shifted(2), 
                           C2 => n163, ZN => n231);
   U219 : NAND2_X1 port map( A1 => n254, A2 => n253, ZN => Y(3));
   U220 : AOI22_X1 port map( A1 => A_neg(3), A2 => n153, B1 => A_signal(3), B2 
                           => n145, ZN => n254);
   U221 : AOI222_X1 port map( A1 => A_shifted(3), A2 => n179, B1 => 
                           zeroSignal(3), B2 => n170, C1 => A_neg_shifted(3), 
                           C2 => n162, ZN => n253);
   U222 : NAND2_X1 port map( A1 => n276, A2 => n275, ZN => Y(4));
   U223 : AOI22_X1 port map( A1 => A_neg(4), A2 => n154, B1 => A_signal(4), B2 
                           => n146, ZN => n276);
   U224 : AOI222_X1 port map( A1 => A_shifted(4), A2 => n180, B1 => 
                           zeroSignal(4), B2 => n171, C1 => A_neg_shifted(4), 
                           C2 => n161, ZN => n275);
   U225 : NAND2_X1 port map( A1 => n298, A2 => n297, ZN => Y(5));
   U226 : AOI22_X1 port map( A1 => A_neg(5), A2 => n155, B1 => A_signal(5), B2 
                           => n147, ZN => n298);
   U227 : AOI222_X1 port map( A1 => A_shifted(5), A2 => n181, B1 => 
                           zeroSignal(5), B2 => n172, C1 => A_neg_shifted(5), 
                           C2 => n160, ZN => n297);
   U228 : AOI222_X1 port map( A1 => A_shifted(57), A2 => n181, B1 => 
                           zeroSignal(57), B2 => n172, C1 => A_neg_shifted(57),
                           C2 => n160, ZN => n291);
   U229 : AOI22_X1 port map( A1 => A_neg(56), A2 => n155, B1 => A_signal(56), 
                           B2 => n147, ZN => n290);
   U230 : AOI222_X1 port map( A1 => A_shifted(60), A2 => n181, B1 => 
                           zeroSignal(60), B2 => n172, C1 => A_neg_shifted(60),
                           C2 => n160, ZN => n299);
   U231 : AOI22_X1 port map( A1 => A_neg(59), A2 => n155, B1 => A_signal(59), 
                           B2 => n147, ZN => n296);
   U232 : AOI222_X1 port map( A1 => A_shifted(55), A2 => n181, B1 => 
                           zeroSignal(55), B2 => n172, C1 => A_neg_shifted(55),
                           C2 => n161, ZN => n287);
   U233 : AOI22_X1 port map( A1 => A_neg(54), A2 => n155, B1 => A_signal(54), 
                           B2 => n147, ZN => n286);
   U234 : AOI222_X1 port map( A1 => A_shifted(53), A2 => n181, B1 => 
                           zeroSignal(53), B2 => n172, C1 => A_neg_shifted(53),
                           C2 => n161, ZN => n283);
   U235 : AOI22_X1 port map( A1 => A_neg(52), A2 => n154, B1 => A_signal(52), 
                           B2 => n146, ZN => n282);
   U236 : AOI222_X1 port map( A1 => A_shifted(54), A2 => n181, B1 => 
                           zeroSignal(54), B2 => n172, C1 => A_neg_shifted(54),
                           C2 => n161, ZN => n285);
   U237 : AOI22_X1 port map( A1 => A_neg(53), A2 => n155, B1 => A_signal(53), 
                           B2 => n147, ZN => n284);
   U238 : AOI222_X1 port map( A1 => A_shifted(51), A2 => n180, B1 => 
                           zeroSignal(51), B2 => n171, C1 => A_neg_shifted(51),
                           C2 => n161, ZN => n279);
   U239 : AOI22_X1 port map( A1 => A_neg(50), A2 => n154, B1 => A_signal(50), 
                           B2 => n146, ZN => n278);
   U240 : AOI222_X1 port map( A1 => A_shifted(7), A2 => n182, B1 => 
                           zeroSignal(7), B2 => n173, C1 => A_neg_shifted(7), 
                           C2 => n160, ZN => n309);
   U241 : AOI22_X1 port map( A1 => A_neg(6), A2 => n156, B1 => A_signal(6), B2 
                           => n148, ZN => n308);
   U242 : NAND2_X1 port map( A1 => n310, A2 => n309, ZN => Y(7));
   U243 : NAND2_X1 port map( A1 => n308, A2 => n307, ZN => Y(6));

end SYN_BEHAVIORAL_2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity MUX51_MuxNbit64_28 is

   port( zeroSignal, A_signal, A_neg, A_shifted, A_neg_shifted : in 
         std_logic_vector (63 downto 0);  Sel : in std_logic_vector (2 downto 
         0);  Y : out std_logic_vector (63 downto 0));

end MUX51_MuxNbit64_28;

architecture SYN_BEHAVIORAL_2 of MUX51_MuxNbit64_28 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, 
      n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, 
      n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, 
      n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, 
      n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, 
      n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, 
      n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, 
      n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, 
      n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, 
      n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, 
      n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, 
      n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, 
      n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, 
      n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, 
      n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318 : 
      std_logic;

begin
   
   U1 : BUF_X1 port map( A => n141, Z => n168);
   U2 : BUF_X1 port map( A => n142, Z => n184);
   U3 : BUF_X1 port map( A => n143, Z => n150);
   U4 : BUF_X1 port map( A => n160, Z => n158);
   U5 : BUF_X1 port map( A => n142, Z => n185);
   U6 : BUF_X1 port map( A => n143, Z => n151);
   U7 : BUF_X1 port map( A => n141, Z => n167);
   U8 : BUF_X1 port map( A => n160, Z => n159);
   U9 : BUF_X1 port map( A => n177, Z => n176);
   U10 : BUF_X1 port map( A => n177, Z => n175);
   U11 : AND3_X1 port map( A1 => n317, A2 => n318, A3 => Sel(2), ZN => n141);
   U12 : NOR3_X1 port map( A1 => n317, A2 => Sel(2), A3 => n318, ZN => n142);
   U13 : NOR3_X1 port map( A1 => Sel(1), A2 => Sel(2), A3 => n317, ZN => n143);
   U14 : BUF_X1 port map( A => n313, Z => n160);
   U15 : BUF_X1 port map( A => n158, Z => n157);
   U16 : BUF_X1 port map( A => n184, Z => n183);
   U17 : BUF_X1 port map( A => n150, Z => n149);
   U18 : BUF_X1 port map( A => n185, Z => n178);
   U19 : BUF_X1 port map( A => n159, Z => n152);
   U20 : BUF_X1 port map( A => n168, Z => n161);
   U21 : BUF_X1 port map( A => n151, Z => n144);
   U22 : BUF_X1 port map( A => n167, Z => n166);
   U23 : BUF_X1 port map( A => n167, Z => n165);
   U24 : BUF_X1 port map( A => n185, Z => n179);
   U25 : BUF_X1 port map( A => n159, Z => n153);
   U26 : BUF_X1 port map( A => n151, Z => n145);
   U27 : BUF_X1 port map( A => n167, Z => n164);
   U28 : BUF_X1 port map( A => n185, Z => n180);
   U29 : BUF_X1 port map( A => n159, Z => n154);
   U30 : BUF_X1 port map( A => n151, Z => n146);
   U31 : BUF_X1 port map( A => n168, Z => n163);
   U32 : BUF_X1 port map( A => n184, Z => n181);
   U33 : BUF_X1 port map( A => n158, Z => n155);
   U34 : BUF_X1 port map( A => n150, Z => n147);
   U35 : BUF_X1 port map( A => n168, Z => n162);
   U36 : BUF_X1 port map( A => n158, Z => n156);
   U37 : BUF_X1 port map( A => n184, Z => n182);
   U38 : BUF_X1 port map( A => n150, Z => n148);
   U39 : BUF_X1 port map( A => n176, Z => n169);
   U40 : BUF_X1 port map( A => n176, Z => n170);
   U41 : BUF_X1 port map( A => n176, Z => n171);
   U42 : BUF_X1 port map( A => n175, Z => n172);
   U43 : BUF_X1 port map( A => n175, Z => n173);
   U44 : BUF_X1 port map( A => n175, Z => n174);
   U45 : INV_X1 port map( A => Sel(1), ZN => n318);
   U46 : NOR3_X1 port map( A1 => Sel(0), A2 => Sel(2), A3 => n318, ZN => n313);
   U47 : INV_X1 port map( A => Sel(0), ZN => n317);
   U48 : BUF_X1 port map( A => n314, Z => n177);
   U49 : NOR2_X1 port map( A1 => n166, A2 => n186, ZN => n314);
   U50 : AOI21_X1 port map( B1 => n317, B2 => n318, A => Sel(2), ZN => n186);
   U51 : AOI22_X1 port map( A1 => A_neg(9), A2 => n157, B1 => A_signal(9), B2 
                           => n149, ZN => n316);
   U52 : AOI222_X1 port map( A1 => A_shifted(8), A2 => n183, B1 => 
                           zeroSignal(8), B2 => n174, C1 => A_neg_shifted(8), 
                           C2 => n161, ZN => n311);
   U53 : NAND2_X1 port map( A1 => n190, A2 => n189, ZN => Y(10));
   U54 : AOI22_X1 port map( A1 => A_neg(10), A2 => n152, B1 => A_signal(10), B2
                           => n144, ZN => n190);
   U55 : AOI222_X1 port map( A1 => A_shifted(10), A2 => n178, B1 => 
                           zeroSignal(10), B2 => n169, C1 => A_neg_shifted(10),
                           C2 => n166, ZN => n189);
   U56 : NAND2_X1 port map( A1 => n192, A2 => n191, ZN => Y(11));
   U57 : AOI22_X1 port map( A1 => A_neg(11), A2 => n152, B1 => A_signal(11), B2
                           => n144, ZN => n192);
   U58 : AOI222_X1 port map( A1 => A_shifted(11), A2 => n178, B1 => 
                           zeroSignal(11), B2 => n169, C1 => A_neg_shifted(11),
                           C2 => n166, ZN => n191);
   U59 : NAND2_X1 port map( A1 => n194, A2 => n193, ZN => Y(12));
   U60 : AOI22_X1 port map( A1 => A_neg(12), A2 => n152, B1 => A_signal(12), B2
                           => n144, ZN => n194);
   U61 : AOI222_X1 port map( A1 => A_shifted(12), A2 => n178, B1 => 
                           zeroSignal(12), B2 => n169, C1 => A_neg_shifted(12),
                           C2 => n166, ZN => n193);
   U62 : NAND2_X1 port map( A1 => n196, A2 => n195, ZN => Y(13));
   U63 : AOI22_X1 port map( A1 => A_neg(13), A2 => n152, B1 => A_signal(13), B2
                           => n144, ZN => n196);
   U64 : AOI222_X1 port map( A1 => A_shifted(13), A2 => n178, B1 => 
                           zeroSignal(13), B2 => n169, C1 => A_neg_shifted(13),
                           C2 => n165, ZN => n195);
   U65 : NAND2_X1 port map( A1 => n198, A2 => n197, ZN => Y(14));
   U66 : AOI22_X1 port map( A1 => A_neg(14), A2 => n152, B1 => A_signal(14), B2
                           => n144, ZN => n198);
   U67 : AOI222_X1 port map( A1 => A_shifted(14), A2 => n178, B1 => 
                           zeroSignal(14), B2 => n169, C1 => A_neg_shifted(14),
                           C2 => n165, ZN => n197);
   U68 : NAND2_X1 port map( A1 => n206, A2 => n205, ZN => Y(18));
   U69 : AOI222_X1 port map( A1 => A_shifted(18), A2 => n178, B1 => 
                           zeroSignal(18), B2 => n169, C1 => A_neg_shifted(18),
                           C2 => n165, ZN => n205);
   U70 : AOI22_X1 port map( A1 => A_neg(18), A2 => n152, B1 => A_signal(18), B2
                           => n144, ZN => n206);
   U71 : NAND2_X1 port map( A1 => n200, A2 => n199, ZN => Y(15));
   U72 : AOI22_X1 port map( A1 => A_neg(15), A2 => n152, B1 => A_signal(15), B2
                           => n144, ZN => n200);
   U73 : AOI222_X1 port map( A1 => A_shifted(15), A2 => n178, B1 => 
                           zeroSignal(15), B2 => n169, C1 => A_neg_shifted(15),
                           C2 => n165, ZN => n199);
   U74 : NAND2_X1 port map( A1 => n208, A2 => n207, ZN => Y(19));
   U75 : AOI222_X1 port map( A1 => A_shifted(19), A2 => n178, B1 => 
                           zeroSignal(19), B2 => n169, C1 => A_neg_shifted(19),
                           C2 => n165, ZN => n207);
   U76 : AOI22_X1 port map( A1 => A_neg(19), A2 => n152, B1 => A_signal(19), B2
                           => n144, ZN => n208);
   U77 : NAND2_X1 port map( A1 => n212, A2 => n211, ZN => Y(20));
   U78 : AOI222_X1 port map( A1 => A_shifted(20), A2 => n179, B1 => 
                           zeroSignal(20), B2 => n170, C1 => A_neg_shifted(20),
                           C2 => n165, ZN => n211);
   U79 : AOI22_X1 port map( A1 => A_neg(20), A2 => n153, B1 => A_signal(20), B2
                           => n145, ZN => n212);
   U80 : NAND2_X1 port map( A1 => n214, A2 => n213, ZN => Y(21));
   U81 : AOI222_X1 port map( A1 => A_shifted(21), A2 => n179, B1 => 
                           zeroSignal(21), B2 => n170, C1 => A_neg_shifted(21),
                           C2 => n165, ZN => n213);
   U82 : AOI22_X1 port map( A1 => A_neg(21), A2 => n153, B1 => A_signal(21), B2
                           => n145, ZN => n214);
   U83 : NAND2_X1 port map( A1 => n220, A2 => n219, ZN => Y(24));
   U84 : AOI222_X1 port map( A1 => A_shifted(24), A2 => n179, B1 => 
                           zeroSignal(24), B2 => n170, C1 => A_neg_shifted(24),
                           C2 => n164, ZN => n219);
   U85 : AOI22_X1 port map( A1 => A_neg(24), A2 => n153, B1 => A_signal(24), B2
                           => n145, ZN => n220);
   U86 : NAND2_X1 port map( A1 => n218, A2 => n217, ZN => Y(23));
   U87 : AOI222_X1 port map( A1 => A_shifted(23), A2 => n179, B1 => 
                           zeroSignal(23), B2 => n170, C1 => A_neg_shifted(23),
                           C2 => n165, ZN => n217);
   U88 : AOI22_X1 port map( A1 => A_neg(23), A2 => n153, B1 => A_signal(23), B2
                           => n145, ZN => n218);
   U89 : NAND2_X1 port map( A1 => n222, A2 => n221, ZN => Y(25));
   U90 : AOI222_X1 port map( A1 => A_shifted(25), A2 => n179, B1 => 
                           zeroSignal(25), B2 => n170, C1 => A_neg_shifted(25),
                           C2 => n164, ZN => n221);
   U91 : AOI22_X1 port map( A1 => A_neg(25), A2 => n153, B1 => A_signal(25), B2
                           => n145, ZN => n222);
   U92 : NAND2_X1 port map( A1 => n216, A2 => n215, ZN => Y(22));
   U93 : AOI22_X1 port map( A1 => A_neg(22), A2 => n153, B1 => A_signal(22), B2
                           => n145, ZN => n216);
   U94 : AOI222_X1 port map( A1 => A_shifted(22), A2 => n179, B1 => 
                           zeroSignal(22), B2 => n170, C1 => A_neg_shifted(22),
                           C2 => n165, ZN => n215);
   U95 : NAND2_X1 port map( A1 => n226, A2 => n225, ZN => Y(27));
   U96 : AOI222_X1 port map( A1 => A_shifted(27), A2 => n179, B1 => 
                           zeroSignal(27), B2 => n170, C1 => A_neg_shifted(27),
                           C2 => n164, ZN => n225);
   U97 : AOI22_X1 port map( A1 => A_neg(27), A2 => n153, B1 => A_signal(27), B2
                           => n145, ZN => n226);
   U98 : NAND2_X1 port map( A1 => n230, A2 => n229, ZN => Y(29));
   U99 : AOI222_X1 port map( A1 => A_shifted(29), A2 => n179, B1 => 
                           zeroSignal(29), B2 => n170, C1 => A_neg_shifted(29),
                           C2 => n164, ZN => n229);
   U100 : AOI22_X1 port map( A1 => A_neg(29), A2 => n153, B1 => A_signal(29), 
                           B2 => n145, ZN => n230);
   U101 : NAND2_X1 port map( A1 => n228, A2 => n227, ZN => Y(28));
   U102 : AOI222_X1 port map( A1 => A_shifted(28), A2 => n179, B1 => 
                           zeroSignal(28), B2 => n170, C1 => A_neg_shifted(28),
                           C2 => n164, ZN => n227);
   U103 : AOI22_X1 port map( A1 => A_neg(28), A2 => n153, B1 => A_signal(28), 
                           B2 => n145, ZN => n228);
   U104 : NAND2_X1 port map( A1 => n202, A2 => n201, ZN => Y(16));
   U105 : AOI22_X1 port map( A1 => A_neg(16), A2 => n152, B1 => A_signal(16), 
                           B2 => n144, ZN => n202);
   U106 : AOI222_X1 port map( A1 => A_shifted(16), A2 => n178, B1 => 
                           zeroSignal(16), B2 => n169, C1 => A_neg_shifted(16),
                           C2 => n165, ZN => n201);
   U107 : NAND2_X1 port map( A1 => n224, A2 => n223, ZN => Y(26));
   U108 : AOI22_X1 port map( A1 => A_neg(26), A2 => n153, B1 => A_signal(26), 
                           B2 => n145, ZN => n224);
   U109 : AOI222_X1 port map( A1 => A_shifted(26), A2 => n179, B1 => 
                           zeroSignal(26), B2 => n170, C1 => A_neg_shifted(26),
                           C2 => n164, ZN => n223);
   U110 : NAND2_X1 port map( A1 => n234, A2 => n233, ZN => Y(30));
   U111 : AOI222_X1 port map( A1 => A_shifted(30), A2 => n179, B1 => 
                           zeroSignal(30), B2 => n170, C1 => A_neg_shifted(30),
                           C2 => n164, ZN => n233);
   U112 : AOI22_X1 port map( A1 => A_neg(30), A2 => n153, B1 => A_signal(30), 
                           B2 => n145, ZN => n234);
   U113 : NAND2_X1 port map( A1 => n236, A2 => n235, ZN => Y(31));
   U114 : AOI222_X1 port map( A1 => A_shifted(31), A2 => n180, B1 => 
                           zeroSignal(31), B2 => n171, C1 => A_neg_shifted(31),
                           C2 => n164, ZN => n235);
   U115 : AOI22_X1 port map( A1 => A_neg(31), A2 => n154, B1 => A_signal(31), 
                           B2 => n146, ZN => n236);
   U116 : NAND2_X1 port map( A1 => n244, A2 => n243, ZN => Y(35));
   U117 : AOI222_X1 port map( A1 => A_shifted(35), A2 => n180, B1 => 
                           zeroSignal(35), B2 => n171, C1 => A_neg_shifted(35),
                           C2 => n163, ZN => n243);
   U118 : AOI22_X1 port map( A1 => A_neg(35), A2 => n154, B1 => A_signal(35), 
                           B2 => n146, ZN => n244);
   U119 : NAND2_X1 port map( A1 => n240, A2 => n239, ZN => Y(33));
   U120 : AOI222_X1 port map( A1 => A_shifted(33), A2 => n180, B1 => 
                           zeroSignal(33), B2 => n171, C1 => A_neg_shifted(33),
                           C2 => n164, ZN => n239);
   U121 : AOI22_X1 port map( A1 => A_neg(33), A2 => n154, B1 => A_signal(33), 
                           B2 => n146, ZN => n240);
   U122 : NAND2_X1 port map( A1 => n242, A2 => n241, ZN => Y(34));
   U123 : AOI222_X1 port map( A1 => A_shifted(34), A2 => n180, B1 => 
                           zeroSignal(34), B2 => n171, C1 => A_neg_shifted(34),
                           C2 => n164, ZN => n241);
   U124 : AOI22_X1 port map( A1 => A_neg(34), A2 => n154, B1 => A_signal(34), 
                           B2 => n146, ZN => n242);
   U125 : NAND2_X1 port map( A1 => n248, A2 => n247, ZN => Y(37));
   U126 : AOI222_X1 port map( A1 => A_shifted(37), A2 => n180, B1 => 
                           zeroSignal(37), B2 => n171, C1 => A_neg_shifted(37),
                           C2 => n163, ZN => n247);
   U127 : AOI22_X1 port map( A1 => A_neg(37), A2 => n154, B1 => A_signal(37), 
                           B2 => n146, ZN => n248);
   U128 : NAND2_X1 port map( A1 => n246, A2 => n245, ZN => Y(36));
   U129 : AOI222_X1 port map( A1 => A_shifted(36), A2 => n180, B1 => 
                           zeroSignal(36), B2 => n171, C1 => A_neg_shifted(36),
                           C2 => n163, ZN => n245);
   U130 : AOI22_X1 port map( A1 => A_neg(36), A2 => n154, B1 => A_signal(36), 
                           B2 => n146, ZN => n246);
   U131 : NAND2_X1 port map( A1 => n238, A2 => n237, ZN => Y(32));
   U132 : AOI22_X1 port map( A1 => A_neg(32), A2 => n154, B1 => A_signal(32), 
                           B2 => n146, ZN => n238);
   U133 : AOI222_X1 port map( A1 => A_shifted(32), A2 => n180, B1 => 
                           zeroSignal(32), B2 => n171, C1 => A_neg_shifted(32),
                           C2 => n164, ZN => n237);
   U134 : NAND2_X1 port map( A1 => n252, A2 => n251, ZN => Y(39));
   U135 : AOI222_X1 port map( A1 => A_shifted(39), A2 => n180, B1 => 
                           zeroSignal(39), B2 => n171, C1 => A_neg_shifted(39),
                           C2 => n163, ZN => n251);
   U136 : AOI22_X1 port map( A1 => A_neg(39), A2 => n154, B1 => A_signal(39), 
                           B2 => n146, ZN => n252);
   U137 : NAND2_X1 port map( A1 => n258, A2 => n257, ZN => Y(41));
   U138 : AOI222_X1 port map( A1 => A_shifted(41), A2 => n180, B1 => 
                           zeroSignal(41), B2 => n171, C1 => A_neg_shifted(41),
                           C2 => n163, ZN => n257);
   U139 : AOI22_X1 port map( A1 => A_neg(41), A2 => n154, B1 => A_signal(41), 
                           B2 => n146, ZN => n258);
   U140 : NAND2_X1 port map( A1 => n204, A2 => n203, ZN => Y(17));
   U141 : AOI22_X1 port map( A1 => A_neg(17), A2 => n152, B1 => A_signal(17), 
                           B2 => n144, ZN => n204);
   U142 : AOI222_X1 port map( A1 => A_shifted(17), A2 => n178, B1 => 
                           zeroSignal(17), B2 => n169, C1 => A_neg_shifted(17),
                           C2 => n165, ZN => n203);
   U143 : NAND2_X1 port map( A1 => n250, A2 => n249, ZN => Y(38));
   U144 : AOI222_X1 port map( A1 => A_shifted(38), A2 => n180, B1 => 
                           zeroSignal(38), B2 => n171, C1 => A_neg_shifted(38),
                           C2 => n163, ZN => n249);
   U145 : AOI22_X1 port map( A1 => A_neg(38), A2 => n154, B1 => A_signal(38), 
                           B2 => n146, ZN => n250);
   U146 : NAND2_X1 port map( A1 => n256, A2 => n255, ZN => Y(40));
   U147 : AOI222_X1 port map( A1 => A_shifted(40), A2 => n180, B1 => 
                           zeroSignal(40), B2 => n171, C1 => A_neg_shifted(40),
                           C2 => n163, ZN => n255);
   U148 : AOI22_X1 port map( A1 => A_neg(40), A2 => n154, B1 => A_signal(40), 
                           B2 => n146, ZN => n256);
   U149 : NAND2_X1 port map( A1 => n270, A2 => n269, ZN => Y(47));
   U150 : AOI222_X1 port map( A1 => A_shifted(47), A2 => n181, B1 => 
                           zeroSignal(47), B2 => n172, C1 => A_neg_shifted(47),
                           C2 => n162, ZN => n269);
   U151 : AOI22_X1 port map( A1 => A_neg(47), A2 => n155, B1 => A_signal(47), 
                           B2 => n147, ZN => n270);
   U152 : NAND2_X1 port map( A1 => n272, A2 => n271, ZN => Y(48));
   U153 : AOI222_X1 port map( A1 => A_shifted(48), A2 => n181, B1 => 
                           zeroSignal(48), B2 => n172, C1 => A_neg_shifted(48),
                           C2 => n162, ZN => n271);
   U154 : AOI22_X1 port map( A1 => A_neg(48), A2 => n155, B1 => A_signal(48), 
                           B2 => n147, ZN => n272);
   U155 : NAND2_X1 port map( A1 => n260, A2 => n259, ZN => Y(42));
   U156 : AOI22_X1 port map( A1 => A_neg(42), A2 => n155, B1 => A_signal(42), 
                           B2 => n147, ZN => n260);
   U157 : AOI222_X1 port map( A1 => A_shifted(42), A2 => n181, B1 => 
                           zeroSignal(42), B2 => n172, C1 => A_neg_shifted(42),
                           C2 => n163, ZN => n259);
   U158 : NAND2_X1 port map( A1 => n274, A2 => n273, ZN => Y(49));
   U159 : AOI22_X1 port map( A1 => A_neg(49), A2 => n155, B1 => A_signal(49), 
                           B2 => n147, ZN => n274);
   U160 : AOI222_X1 port map( A1 => A_shifted(49), A2 => n181, B1 => 
                           zeroSignal(49), B2 => n172, C1 => A_neg_shifted(49),
                           C2 => n162, ZN => n273);
   U161 : NAND2_X1 port map( A1 => n262, A2 => n261, ZN => Y(43));
   U162 : AOI222_X1 port map( A1 => A_shifted(43), A2 => n181, B1 => 
                           zeroSignal(43), B2 => n172, C1 => A_neg_shifted(43),
                           C2 => n163, ZN => n261);
   U163 : AOI22_X1 port map( A1 => A_neg(43), A2 => n155, B1 => A_signal(43), 
                           B2 => n147, ZN => n262);
   U164 : NAND2_X1 port map( A1 => n264, A2 => n263, ZN => Y(44));
   U165 : AOI222_X1 port map( A1 => A_shifted(44), A2 => n181, B1 => 
                           zeroSignal(44), B2 => n172, C1 => A_neg_shifted(44),
                           C2 => n163, ZN => n263);
   U166 : AOI22_X1 port map( A1 => A_neg(44), A2 => n155, B1 => A_signal(44), 
                           B2 => n147, ZN => n264);
   U167 : NAND2_X1 port map( A1 => n304, A2 => n303, ZN => Y(62));
   U168 : AOI22_X1 port map( A1 => A_neg(62), A2 => n156, B1 => A_signal(62), 
                           B2 => n148, ZN => n304);
   U169 : NAND2_X1 port map( A1 => n306, A2 => n305, ZN => Y(63));
   U170 : AOI222_X1 port map( A1 => A_shifted(63), A2 => n182, B1 => 
                           zeroSignal(63), B2 => n173, C1 => A_neg_shifted(63),
                           C2 => n161, ZN => n305);
   U171 : AOI22_X1 port map( A1 => A_neg(63), A2 => n156, B1 => A_signal(63), 
                           B2 => n148, ZN => n306);
   U172 : NAND2_X1 port map( A1 => n266, A2 => n265, ZN => Y(45));
   U173 : AOI22_X1 port map( A1 => A_neg(45), A2 => n155, B1 => A_signal(45), 
                           B2 => n147, ZN => n266);
   U174 : AOI222_X1 port map( A1 => A_shifted(45), A2 => n181, B1 => 
                           zeroSignal(45), B2 => n172, C1 => A_neg_shifted(45),
                           C2 => n163, ZN => n265);
   U175 : NAND2_X1 port map( A1 => n282, A2 => n281, ZN => Y(52));
   U176 : AOI222_X1 port map( A1 => A_shifted(52), A2 => n181, B1 => 
                           zeroSignal(52), B2 => n172, C1 => A_neg_shifted(52),
                           C2 => n162, ZN => n281);
   U177 : NAND2_X1 port map( A1 => n284, A2 => n283, ZN => Y(53));
   U178 : AOI22_X1 port map( A1 => A_neg(53), A2 => n156, B1 => A_signal(53), 
                           B2 => n148, ZN => n284);
   U179 : NAND2_X1 port map( A1 => n280, A2 => n279, ZN => Y(51));
   U180 : AOI222_X1 port map( A1 => A_shifted(51), A2 => n181, B1 => 
                           zeroSignal(51), B2 => n172, C1 => A_neg_shifted(51),
                           C2 => n162, ZN => n279);
   U181 : AOI22_X1 port map( A1 => A_neg(51), A2 => n155, B1 => A_signal(51), 
                           B2 => n147, ZN => n280);
   U182 : NAND2_X1 port map( A1 => n302, A2 => n301, ZN => Y(61));
   U183 : AOI222_X1 port map( A1 => A_shifted(61), A2 => n182, B1 => 
                           zeroSignal(61), B2 => n173, C1 => A_neg_shifted(61),
                           C2 => n161, ZN => n301);
   U184 : NAND2_X1 port map( A1 => n286, A2 => n285, ZN => Y(54));
   U185 : AOI222_X1 port map( A1 => A_shifted(54), A2 => n182, B1 => 
                           zeroSignal(54), B2 => n173, C1 => A_neg_shifted(54),
                           C2 => n162, ZN => n285);
   U186 : NAND2_X1 port map( A1 => n288, A2 => n287, ZN => Y(55));
   U187 : NAND2_X1 port map( A1 => n290, A2 => n289, ZN => Y(56));
   U188 : NAND2_X1 port map( A1 => n294, A2 => n293, ZN => Y(58));
   U189 : AOI222_X1 port map( A1 => A_shifted(58), A2 => n182, B1 => 
                           zeroSignal(58), B2 => n173, C1 => A_neg_shifted(58),
                           C2 => n161, ZN => n293);
   U190 : NAND2_X1 port map( A1 => n278, A2 => n277, ZN => Y(50));
   U191 : AOI22_X1 port map( A1 => A_neg(50), A2 => n155, B1 => A_signal(50), 
                           B2 => n147, ZN => n278);
   U192 : AOI222_X1 port map( A1 => A_shifted(50), A2 => n181, B1 => 
                           zeroSignal(50), B2 => n172, C1 => A_neg_shifted(50),
                           C2 => n162, ZN => n277);
   U193 : NAND2_X1 port map( A1 => n300, A2 => n299, ZN => Y(60));
   U194 : AOI222_X1 port map( A1 => A_shifted(60), A2 => n182, B1 => 
                           zeroSignal(60), B2 => n173, C1 => A_neg_shifted(60),
                           C2 => n161, ZN => n299);
   U195 : AOI22_X1 port map( A1 => A_neg(60), A2 => n156, B1 => A_signal(60), 
                           B2 => n148, ZN => n300);
   U196 : NAND2_X1 port map( A1 => n296, A2 => n295, ZN => Y(59));
   U197 : AOI22_X1 port map( A1 => A_neg(59), A2 => n156, B1 => A_signal(59), 
                           B2 => n148, ZN => n296);
   U198 : NAND2_X1 port map( A1 => n292, A2 => n291, ZN => Y(57));
   U199 : AOI22_X1 port map( A1 => A_neg(57), A2 => n156, B1 => A_signal(57), 
                           B2 => n148, ZN => n292);
   U200 : NAND2_X1 port map( A1 => n268, A2 => n267, ZN => Y(46));
   U201 : AOI22_X1 port map( A1 => A_neg(46), A2 => n155, B1 => A_signal(46), 
                           B2 => n147, ZN => n268);
   U202 : AOI222_X1 port map( A1 => A_shifted(46), A2 => n181, B1 => 
                           zeroSignal(46), B2 => n172, C1 => A_neg_shifted(46),
                           C2 => n162, ZN => n267);
   U203 : NAND2_X1 port map( A1 => n188, A2 => n187, ZN => Y(0));
   U204 : AOI22_X1 port map( A1 => A_neg(0), A2 => n152, B1 => A_signal(0), B2 
                           => n144, ZN => n188);
   U205 : AOI222_X1 port map( A1 => A_shifted(0), A2 => n178, B1 => 
                           zeroSignal(0), B2 => n169, C1 => A_neg_shifted(0), 
                           C2 => n166, ZN => n187);
   U206 : NAND2_X1 port map( A1 => n210, A2 => n209, ZN => Y(1));
   U207 : AOI22_X1 port map( A1 => A_neg(1), A2 => n152, B1 => A_signal(1), B2 
                           => n144, ZN => n210);
   U208 : AOI222_X1 port map( A1 => A_shifted(1), A2 => n178, B1 => 
                           zeroSignal(1), B2 => n169, C1 => A_neg_shifted(1), 
                           C2 => n165, ZN => n209);
   U209 : NAND2_X1 port map( A1 => n232, A2 => n231, ZN => Y(2));
   U210 : AOI22_X1 port map( A1 => A_neg(2), A2 => n153, B1 => A_signal(2), B2 
                           => n145, ZN => n232);
   U211 : AOI222_X1 port map( A1 => A_shifted(2), A2 => n179, B1 => 
                           zeroSignal(2), B2 => n170, C1 => A_neg_shifted(2), 
                           C2 => n164, ZN => n231);
   U212 : NAND2_X1 port map( A1 => n254, A2 => n253, ZN => Y(3));
   U213 : AOI22_X1 port map( A1 => A_neg(3), A2 => n154, B1 => A_signal(3), B2 
                           => n146, ZN => n254);
   U214 : AOI222_X1 port map( A1 => A_shifted(3), A2 => n180, B1 => 
                           zeroSignal(3), B2 => n171, C1 => A_neg_shifted(3), 
                           C2 => n163, ZN => n253);
   U215 : NAND2_X1 port map( A1 => n276, A2 => n275, ZN => Y(4));
   U216 : AOI22_X1 port map( A1 => A_neg(4), A2 => n155, B1 => A_signal(4), B2 
                           => n147, ZN => n276);
   U217 : AOI222_X1 port map( A1 => A_shifted(4), A2 => n181, B1 => 
                           zeroSignal(4), B2 => n172, C1 => A_neg_shifted(4), 
                           C2 => n162, ZN => n275);
   U218 : NAND2_X1 port map( A1 => n298, A2 => n297, ZN => Y(5));
   U219 : AOI22_X1 port map( A1 => A_neg(5), A2 => n156, B1 => A_signal(5), B2 
                           => n148, ZN => n298);
   U220 : AOI222_X1 port map( A1 => A_shifted(5), A2 => n182, B1 => 
                           zeroSignal(5), B2 => n173, C1 => A_neg_shifted(5), 
                           C2 => n161, ZN => n297);
   U221 : NAND2_X1 port map( A1 => n308, A2 => n307, ZN => Y(6));
   U222 : AOI22_X1 port map( A1 => A_neg(6), A2 => n157, B1 => A_signal(6), B2 
                           => n149, ZN => n308);
   U223 : AOI222_X1 port map( A1 => A_shifted(6), A2 => n183, B1 => 
                           zeroSignal(6), B2 => n174, C1 => A_neg_shifted(6), 
                           C2 => n161, ZN => n307);
   U224 : NAND2_X1 port map( A1 => n310, A2 => n309, ZN => Y(7));
   U225 : AOI22_X1 port map( A1 => A_neg(7), A2 => n157, B1 => A_signal(7), B2 
                           => n149, ZN => n310);
   U226 : AOI222_X1 port map( A1 => A_shifted(7), A2 => n183, B1 => 
                           zeroSignal(7), B2 => n174, C1 => A_neg_shifted(7), 
                           C2 => n161, ZN => n309);
   U227 : AOI222_X1 port map( A1 => A_shifted(59), A2 => n182, B1 => 
                           zeroSignal(59), B2 => n173, C1 => A_neg_shifted(59),
                           C2 => n161, ZN => n295);
   U228 : AOI22_X1 port map( A1 => A_neg(58), A2 => n156, B1 => A_signal(58), 
                           B2 => n148, ZN => n294);
   U229 : AOI222_X1 port map( A1 => A_shifted(62), A2 => n182, B1 => 
                           zeroSignal(62), B2 => n173, C1 => A_neg_shifted(62),
                           C2 => n161, ZN => n303);
   U230 : AOI22_X1 port map( A1 => A_neg(61), A2 => n156, B1 => A_signal(61), 
                           B2 => n148, ZN => n302);
   U231 : AOI222_X1 port map( A1 => A_shifted(57), A2 => n182, B1 => 
                           zeroSignal(57), B2 => n173, C1 => A_neg_shifted(57),
                           C2 => n161, ZN => n291);
   U232 : AOI22_X1 port map( A1 => A_neg(56), A2 => n156, B1 => A_signal(56), 
                           B2 => n148, ZN => n290);
   U233 : AOI222_X1 port map( A1 => A_shifted(55), A2 => n182, B1 => 
                           zeroSignal(55), B2 => n173, C1 => A_neg_shifted(55),
                           C2 => n162, ZN => n287);
   U234 : AOI22_X1 port map( A1 => A_neg(54), A2 => n156, B1 => A_signal(54), 
                           B2 => n148, ZN => n286);
   U235 : AOI222_X1 port map( A1 => A_shifted(56), A2 => n182, B1 => 
                           zeroSignal(56), B2 => n173, C1 => A_neg_shifted(56),
                           C2 => n162, ZN => n289);
   U236 : AOI22_X1 port map( A1 => A_neg(55), A2 => n156, B1 => A_signal(55), 
                           B2 => n148, ZN => n288);
   U237 : AOI222_X1 port map( A1 => A_shifted(53), A2 => n182, B1 => 
                           zeroSignal(53), B2 => n173, C1 => A_neg_shifted(53),
                           C2 => n162, ZN => n283);
   U238 : AOI22_X1 port map( A1 => A_neg(52), A2 => n155, B1 => A_signal(52), 
                           B2 => n147, ZN => n282);
   U239 : AOI222_X1 port map( A1 => A_shifted(9), A2 => n183, B1 => 
                           zeroSignal(9), B2 => n174, C1 => A_neg_shifted(9), 
                           C2 => n161, ZN => n315);
   U240 : AOI22_X1 port map( A1 => A_neg(8), A2 => n157, B1 => A_signal(8), B2 
                           => n149, ZN => n312);
   U241 : NAND2_X1 port map( A1 => n316, A2 => n315, ZN => Y(9));
   U242 : NAND2_X1 port map( A1 => n312, A2 => n311, ZN => Y(8));

end SYN_BEHAVIORAL_2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity MUX51_MuxNbit64_27 is

   port( zeroSignal, A_signal, A_neg, A_shifted, A_neg_shifted : in 
         std_logic_vector (63 downto 0);  Sel : in std_logic_vector (2 downto 
         0);  Y : out std_logic_vector (63 downto 0));

end MUX51_MuxNbit64_27;

architecture SYN_BEHAVIORAL_2 of MUX51_MuxNbit64_27 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, 
      n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, 
      n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, 
      n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, 
      n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, 
      n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, 
      n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, 
      n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, 
      n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, 
      n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, 
      n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, 
      n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, 
      n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, 
      n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, 
      n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319 : 
      std_logic;

begin
   
   U1 : BUF_X1 port map( A => n141, Z => n185);
   U2 : BUF_X1 port map( A => n142, Z => n167);
   U3 : BUF_X1 port map( A => n160, Z => n159);
   U4 : BUF_X1 port map( A => n151, Z => n150);
   U5 : BUF_X1 port map( A => n142, Z => n168);
   U6 : BUF_X1 port map( A => n141, Z => n184);
   U7 : BUF_X1 port map( A => n160, Z => n158);
   U8 : BUF_X1 port map( A => n151, Z => n149);
   U9 : BUF_X1 port map( A => n177, Z => n176);
   U10 : BUF_X1 port map( A => n177, Z => n175);
   U11 : NOR3_X1 port map( A1 => n318, A2 => Sel(2), A3 => n319, ZN => n141);
   U12 : AND3_X1 port map( A1 => n318, A2 => n319, A3 => Sel(2), ZN => n142);
   U13 : BUF_X1 port map( A => n159, Z => n152);
   U14 : BUF_X1 port map( A => n185, Z => n178);
   U15 : BUF_X1 port map( A => n150, Z => n143);
   U16 : BUF_X1 port map( A => n167, Z => n166);
   U17 : BUF_X1 port map( A => n167, Z => n165);
   U18 : BUF_X1 port map( A => n185, Z => n179);
   U19 : BUF_X1 port map( A => n159, Z => n153);
   U20 : BUF_X1 port map( A => n150, Z => n144);
   U21 : BUF_X1 port map( A => n167, Z => n164);
   U22 : BUF_X1 port map( A => n185, Z => n180);
   U23 : BUF_X1 port map( A => n159, Z => n154);
   U24 : BUF_X1 port map( A => n150, Z => n145);
   U25 : BUF_X1 port map( A => n168, Z => n163);
   U26 : BUF_X1 port map( A => n184, Z => n181);
   U27 : BUF_X1 port map( A => n158, Z => n155);
   U28 : BUF_X1 port map( A => n149, Z => n146);
   U29 : BUF_X1 port map( A => n168, Z => n162);
   U30 : BUF_X1 port map( A => n158, Z => n156);
   U31 : BUF_X1 port map( A => n184, Z => n182);
   U32 : BUF_X1 port map( A => n149, Z => n147);
   U33 : BUF_X1 port map( A => n168, Z => n161);
   U34 : BUF_X1 port map( A => n176, Z => n170);
   U35 : BUF_X1 port map( A => n176, Z => n171);
   U36 : BUF_X1 port map( A => n175, Z => n172);
   U37 : BUF_X1 port map( A => n176, Z => n169);
   U38 : BUF_X1 port map( A => n175, Z => n173);
   U39 : BUF_X1 port map( A => n158, Z => n157);
   U40 : BUF_X1 port map( A => n149, Z => n148);
   U41 : BUF_X1 port map( A => n175, Z => n174);
   U42 : BUF_X1 port map( A => n184, Z => n183);
   U43 : INV_X1 port map( A => Sel(1), ZN => n319);
   U44 : BUF_X1 port map( A => n314, Z => n160);
   U45 : NOR3_X1 port map( A1 => Sel(0), A2 => Sel(2), A3 => n319, ZN => n314);
   U46 : INV_X1 port map( A => Sel(0), ZN => n318);
   U47 : BUF_X1 port map( A => n313, Z => n151);
   U48 : NOR3_X1 port map( A1 => Sel(1), A2 => Sel(2), A3 => n318, ZN => n313);
   U49 : BUF_X1 port map( A => n315, Z => n177);
   U50 : NOR2_X1 port map( A1 => n166, A2 => n186, ZN => n315);
   U51 : AOI21_X1 port map( B1 => n318, B2 => n319, A => Sel(2), ZN => n186);
   U52 : AOI22_X1 port map( A1 => A_neg(11), A2 => n152, B1 => A_signal(11), B2
                           => n143, ZN => n192);
   U53 : AOI222_X1 port map( A1 => A_shifted(10), A2 => n178, B1 => 
                           zeroSignal(10), B2 => n169, C1 => A_neg_shifted(10),
                           C2 => n166, ZN => n189);
   U54 : NAND2_X1 port map( A1 => n194, A2 => n193, ZN => Y(12));
   U55 : AOI22_X1 port map( A1 => A_neg(12), A2 => n152, B1 => A_signal(12), B2
                           => n143, ZN => n194);
   U56 : AOI222_X1 port map( A1 => A_shifted(12), A2 => n178, B1 => 
                           zeroSignal(12), B2 => n169, C1 => A_neg_shifted(12),
                           C2 => n166, ZN => n193);
   U57 : NAND2_X1 port map( A1 => n196, A2 => n195, ZN => Y(13));
   U58 : AOI22_X1 port map( A1 => A_neg(13), A2 => n152, B1 => A_signal(13), B2
                           => n143, ZN => n196);
   U59 : AOI222_X1 port map( A1 => A_shifted(13), A2 => n178, B1 => 
                           zeroSignal(13), B2 => n169, C1 => A_neg_shifted(13),
                           C2 => n165, ZN => n195);
   U60 : NAND2_X1 port map( A1 => n198, A2 => n197, ZN => Y(14));
   U61 : AOI22_X1 port map( A1 => A_neg(14), A2 => n152, B1 => A_signal(14), B2
                           => n143, ZN => n198);
   U62 : AOI222_X1 port map( A1 => A_shifted(14), A2 => n178, B1 => 
                           zeroSignal(14), B2 => n169, C1 => A_neg_shifted(14),
                           C2 => n165, ZN => n197);
   U63 : NAND2_X1 port map( A1 => n200, A2 => n199, ZN => Y(15));
   U64 : AOI22_X1 port map( A1 => A_neg(15), A2 => n152, B1 => A_signal(15), B2
                           => n143, ZN => n200);
   U65 : AOI222_X1 port map( A1 => A_shifted(15), A2 => n178, B1 => 
                           zeroSignal(15), B2 => n169, C1 => A_neg_shifted(15),
                           C2 => n165, ZN => n199);
   U66 : NAND2_X1 port map( A1 => n202, A2 => n201, ZN => Y(16));
   U67 : AOI22_X1 port map( A1 => A_neg(16), A2 => n152, B1 => A_signal(16), B2
                           => n143, ZN => n202);
   U68 : AOI222_X1 port map( A1 => A_shifted(16), A2 => n178, B1 => 
                           zeroSignal(16), B2 => n169, C1 => A_neg_shifted(16),
                           C2 => n165, ZN => n201);
   U69 : NAND2_X1 port map( A1 => n306, A2 => n305, ZN => Y(63));
   U70 : AOI222_X1 port map( A1 => A_shifted(63), A2 => n182, B1 => 
                           zeroSignal(63), B2 => n173, C1 => A_neg_shifted(63),
                           C2 => n161, ZN => n305);
   U71 : NAND2_X1 port map( A1 => n204, A2 => n203, ZN => Y(17));
   U72 : AOI22_X1 port map( A1 => A_neg(17), A2 => n152, B1 => A_signal(17), B2
                           => n143, ZN => n204);
   U73 : AOI222_X1 port map( A1 => A_shifted(17), A2 => n178, B1 => 
                           zeroSignal(17), B2 => n169, C1 => A_neg_shifted(17),
                           C2 => n165, ZN => n203);
   U74 : NAND2_X1 port map( A1 => n212, A2 => n211, ZN => Y(20));
   U75 : AOI222_X1 port map( A1 => A_shifted(20), A2 => n179, B1 => 
                           zeroSignal(20), B2 => n170, C1 => A_neg_shifted(20),
                           C2 => n165, ZN => n211);
   U76 : AOI22_X1 port map( A1 => A_neg(20), A2 => n153, B1 => A_signal(20), B2
                           => n144, ZN => n212);
   U77 : NAND2_X1 port map( A1 => n214, A2 => n213, ZN => Y(21));
   U78 : AOI222_X1 port map( A1 => A_shifted(21), A2 => n179, B1 => 
                           zeroSignal(21), B2 => n170, C1 => A_neg_shifted(21),
                           C2 => n165, ZN => n213);
   U79 : AOI22_X1 port map( A1 => A_neg(21), A2 => n153, B1 => A_signal(21), B2
                           => n144, ZN => n214);
   U80 : NAND2_X1 port map( A1 => n216, A2 => n215, ZN => Y(22));
   U81 : AOI222_X1 port map( A1 => A_shifted(22), A2 => n179, B1 => 
                           zeroSignal(22), B2 => n170, C1 => A_neg_shifted(22),
                           C2 => n165, ZN => n215);
   U82 : AOI22_X1 port map( A1 => A_neg(22), A2 => n153, B1 => A_signal(22), B2
                           => n144, ZN => n216);
   U83 : NAND2_X1 port map( A1 => n218, A2 => n217, ZN => Y(23));
   U84 : AOI222_X1 port map( A1 => A_shifted(23), A2 => n179, B1 => 
                           zeroSignal(23), B2 => n170, C1 => A_neg_shifted(23),
                           C2 => n165, ZN => n217);
   U85 : AOI22_X1 port map( A1 => A_neg(23), A2 => n153, B1 => A_signal(23), B2
                           => n144, ZN => n218);
   U86 : NAND2_X1 port map( A1 => n222, A2 => n221, ZN => Y(25));
   U87 : AOI222_X1 port map( A1 => A_shifted(25), A2 => n179, B1 => 
                           zeroSignal(25), B2 => n170, C1 => A_neg_shifted(25),
                           C2 => n164, ZN => n221);
   U88 : AOI22_X1 port map( A1 => A_neg(25), A2 => n153, B1 => A_signal(25), B2
                           => n144, ZN => n222);
   U89 : NAND2_X1 port map( A1 => n224, A2 => n223, ZN => Y(26));
   U90 : AOI222_X1 port map( A1 => A_shifted(26), A2 => n179, B1 => 
                           zeroSignal(26), B2 => n170, C1 => A_neg_shifted(26),
                           C2 => n164, ZN => n223);
   U91 : AOI22_X1 port map( A1 => A_neg(26), A2 => n153, B1 => A_signal(26), B2
                           => n144, ZN => n224);
   U92 : NAND2_X1 port map( A1 => n226, A2 => n225, ZN => Y(27));
   U93 : AOI222_X1 port map( A1 => A_shifted(27), A2 => n179, B1 => 
                           zeroSignal(27), B2 => n170, C1 => A_neg_shifted(27),
                           C2 => n164, ZN => n225);
   U94 : AOI22_X1 port map( A1 => A_neg(27), A2 => n153, B1 => A_signal(27), B2
                           => n144, ZN => n226);
   U95 : NAND2_X1 port map( A1 => n220, A2 => n219, ZN => Y(24));
   U96 : AOI22_X1 port map( A1 => A_neg(24), A2 => n153, B1 => A_signal(24), B2
                           => n144, ZN => n220);
   U97 : AOI222_X1 port map( A1 => A_shifted(24), A2 => n179, B1 => 
                           zeroSignal(24), B2 => n170, C1 => A_neg_shifted(24),
                           C2 => n164, ZN => n219);
   U98 : NAND2_X1 port map( A1 => n206, A2 => n205, ZN => Y(18));
   U99 : AOI22_X1 port map( A1 => A_neg(18), A2 => n152, B1 => A_signal(18), B2
                           => n143, ZN => n206);
   U100 : AOI222_X1 port map( A1 => A_shifted(18), A2 => n178, B1 => 
                           zeroSignal(18), B2 => n169, C1 => A_neg_shifted(18),
                           C2 => n165, ZN => n205);
   U101 : NAND2_X1 port map( A1 => n270, A2 => n269, ZN => Y(47));
   U102 : AOI22_X1 port map( A1 => A_neg(47), A2 => n155, B1 => A_signal(47), 
                           B2 => n146, ZN => n270);
   U103 : AOI222_X1 port map( A1 => A_shifted(47), A2 => n181, B1 => 
                           zeroSignal(47), B2 => n172, C1 => A_neg_shifted(47),
                           C2 => n162, ZN => n269);
   U104 : NAND2_X1 port map( A1 => n230, A2 => n229, ZN => Y(29));
   U105 : AOI222_X1 port map( A1 => A_shifted(29), A2 => n179, B1 => 
                           zeroSignal(29), B2 => n170, C1 => A_neg_shifted(29),
                           C2 => n164, ZN => n229);
   U106 : AOI22_X1 port map( A1 => A_neg(29), A2 => n153, B1 => A_signal(29), 
                           B2 => n144, ZN => n230);
   U107 : NAND2_X1 port map( A1 => n234, A2 => n233, ZN => Y(30));
   U108 : AOI222_X1 port map( A1 => A_shifted(30), A2 => n179, B1 => 
                           zeroSignal(30), B2 => n170, C1 => A_neg_shifted(30),
                           C2 => n164, ZN => n233);
   U109 : AOI22_X1 port map( A1 => A_neg(30), A2 => n153, B1 => A_signal(30), 
                           B2 => n144, ZN => n234);
   U110 : NAND2_X1 port map( A1 => n236, A2 => n235, ZN => Y(31));
   U111 : AOI222_X1 port map( A1 => A_shifted(31), A2 => n180, B1 => 
                           zeroSignal(31), B2 => n171, C1 => A_neg_shifted(31),
                           C2 => n164, ZN => n235);
   U112 : AOI22_X1 port map( A1 => A_neg(31), A2 => n154, B1 => A_signal(31), 
                           B2 => n145, ZN => n236);
   U113 : NAND2_X1 port map( A1 => n238, A2 => n237, ZN => Y(32));
   U114 : AOI222_X1 port map( A1 => A_shifted(32), A2 => n180, B1 => 
                           zeroSignal(32), B2 => n171, C1 => A_neg_shifted(32),
                           C2 => n164, ZN => n237);
   U115 : AOI22_X1 port map( A1 => A_neg(32), A2 => n154, B1 => A_signal(32), 
                           B2 => n145, ZN => n238);
   U116 : NAND2_X1 port map( A1 => n228, A2 => n227, ZN => Y(28));
   U117 : AOI22_X1 port map( A1 => A_neg(28), A2 => n153, B1 => A_signal(28), 
                           B2 => n144, ZN => n228);
   U118 : AOI222_X1 port map( A1 => A_shifted(28), A2 => n179, B1 => 
                           zeroSignal(28), B2 => n170, C1 => A_neg_shifted(28),
                           C2 => n164, ZN => n227);
   U119 : NAND2_X1 port map( A1 => n244, A2 => n243, ZN => Y(35));
   U120 : AOI222_X1 port map( A1 => A_shifted(35), A2 => n180, B1 => 
                           zeroSignal(35), B2 => n171, C1 => A_neg_shifted(35),
                           C2 => n163, ZN => n243);
   U121 : AOI22_X1 port map( A1 => A_neg(35), A2 => n154, B1 => A_signal(35), 
                           B2 => n145, ZN => n244);
   U122 : NAND2_X1 port map( A1 => n240, A2 => n239, ZN => Y(33));
   U123 : AOI222_X1 port map( A1 => A_shifted(33), A2 => n180, B1 => 
                           zeroSignal(33), B2 => n171, C1 => A_neg_shifted(33),
                           C2 => n164, ZN => n239);
   U124 : AOI22_X1 port map( A1 => A_neg(33), A2 => n154, B1 => A_signal(33), 
                           B2 => n145, ZN => n240);
   U125 : NAND2_X1 port map( A1 => n248, A2 => n247, ZN => Y(37));
   U126 : AOI222_X1 port map( A1 => A_shifted(37), A2 => n180, B1 => 
                           zeroSignal(37), B2 => n171, C1 => A_neg_shifted(37),
                           C2 => n163, ZN => n247);
   U127 : AOI22_X1 port map( A1 => A_neg(37), A2 => n154, B1 => A_signal(37), 
                           B2 => n145, ZN => n248);
   U128 : NAND2_X1 port map( A1 => n246, A2 => n245, ZN => Y(36));
   U129 : AOI222_X1 port map( A1 => A_shifted(36), A2 => n180, B1 => 
                           zeroSignal(36), B2 => n171, C1 => A_neg_shifted(36),
                           C2 => n163, ZN => n245);
   U130 : AOI22_X1 port map( A1 => A_neg(36), A2 => n154, B1 => A_signal(36), 
                           B2 => n145, ZN => n246);
   U131 : NAND2_X1 port map( A1 => n252, A2 => n251, ZN => Y(39));
   U132 : AOI222_X1 port map( A1 => A_shifted(39), A2 => n180, B1 => 
                           zeroSignal(39), B2 => n171, C1 => A_neg_shifted(39),
                           C2 => n163, ZN => n251);
   U133 : AOI22_X1 port map( A1 => A_neg(39), A2 => n154, B1 => A_signal(39), 
                           B2 => n145, ZN => n252);
   U134 : NAND2_X1 port map( A1 => n242, A2 => n241, ZN => Y(34));
   U135 : AOI22_X1 port map( A1 => A_neg(34), A2 => n154, B1 => A_signal(34), 
                           B2 => n145, ZN => n242);
   U136 : AOI222_X1 port map( A1 => A_shifted(34), A2 => n180, B1 => 
                           zeroSignal(34), B2 => n171, C1 => A_neg_shifted(34),
                           C2 => n164, ZN => n241);
   U137 : NAND2_X1 port map( A1 => n208, A2 => n207, ZN => Y(19));
   U138 : AOI22_X1 port map( A1 => A_neg(19), A2 => n152, B1 => A_signal(19), 
                           B2 => n143, ZN => n208);
   U139 : AOI222_X1 port map( A1 => A_shifted(19), A2 => n178, B1 => 
                           zeroSignal(19), B2 => n169, C1 => A_neg_shifted(19),
                           C2 => n165, ZN => n207);
   U140 : NAND2_X1 port map( A1 => n250, A2 => n249, ZN => Y(38));
   U141 : AOI222_X1 port map( A1 => A_shifted(38), A2 => n180, B1 => 
                           zeroSignal(38), B2 => n171, C1 => A_neg_shifted(38),
                           C2 => n163, ZN => n249);
   U142 : AOI22_X1 port map( A1 => A_neg(38), A2 => n154, B1 => A_signal(38), 
                           B2 => n145, ZN => n250);
   U143 : NAND2_X1 port map( A1 => n256, A2 => n255, ZN => Y(40));
   U144 : AOI222_X1 port map( A1 => A_shifted(40), A2 => n180, B1 => 
                           zeroSignal(40), B2 => n171, C1 => A_neg_shifted(40),
                           C2 => n163, ZN => n255);
   U145 : AOI22_X1 port map( A1 => A_neg(40), A2 => n154, B1 => A_signal(40), 
                           B2 => n145, ZN => n256);
   U146 : NAND2_X1 port map( A1 => n262, A2 => n261, ZN => Y(43));
   U147 : AOI222_X1 port map( A1 => A_shifted(43), A2 => n181, B1 => 
                           zeroSignal(43), B2 => n172, C1 => A_neg_shifted(43),
                           C2 => n163, ZN => n261);
   U148 : AOI22_X1 port map( A1 => A_neg(43), A2 => n155, B1 => A_signal(43), 
                           B2 => n146, ZN => n262);
   U149 : NAND2_X1 port map( A1 => n258, A2 => n257, ZN => Y(41));
   U150 : AOI222_X1 port map( A1 => A_shifted(41), A2 => n180, B1 => 
                           zeroSignal(41), B2 => n171, C1 => A_neg_shifted(41),
                           C2 => n163, ZN => n257);
   U151 : AOI22_X1 port map( A1 => A_neg(41), A2 => n154, B1 => A_signal(41), 
                           B2 => n145, ZN => n258);
   U152 : NAND2_X1 port map( A1 => n274, A2 => n273, ZN => Y(49));
   U153 : AOI222_X1 port map( A1 => A_shifted(49), A2 => n181, B1 => 
                           zeroSignal(49), B2 => n172, C1 => A_neg_shifted(49),
                           C2 => n162, ZN => n273);
   U154 : AOI22_X1 port map( A1 => A_neg(49), A2 => n155, B1 => A_signal(49), 
                           B2 => n146, ZN => n274);
   U155 : NAND2_X1 port map( A1 => n260, A2 => n259, ZN => Y(42));
   U156 : AOI222_X1 port map( A1 => A_shifted(42), A2 => n181, B1 => 
                           zeroSignal(42), B2 => n172, C1 => A_neg_shifted(42),
                           C2 => n163, ZN => n259);
   U157 : AOI22_X1 port map( A1 => A_neg(42), A2 => n155, B1 => A_signal(42), 
                           B2 => n146, ZN => n260);
   U158 : NAND2_X1 port map( A1 => n278, A2 => n277, ZN => Y(50));
   U159 : AOI222_X1 port map( A1 => A_shifted(50), A2 => n181, B1 => 
                           zeroSignal(50), B2 => n172, C1 => A_neg_shifted(50),
                           C2 => n162, ZN => n277);
   U160 : AOI22_X1 port map( A1 => A_neg(50), A2 => n155, B1 => A_signal(50), 
                           B2 => n146, ZN => n278);
   U161 : NAND2_X1 port map( A1 => n272, A2 => n271, ZN => Y(48));
   U162 : AOI222_X1 port map( A1 => A_shifted(48), A2 => n181, B1 => 
                           zeroSignal(48), B2 => n172, C1 => A_neg_shifted(48),
                           C2 => n162, ZN => n271);
   U163 : AOI22_X1 port map( A1 => A_neg(48), A2 => n155, B1 => A_signal(48), 
                           B2 => n146, ZN => n272);
   U164 : NAND2_X1 port map( A1 => n264, A2 => n263, ZN => Y(44));
   U165 : AOI222_X1 port map( A1 => A_shifted(44), A2 => n181, B1 => 
                           zeroSignal(44), B2 => n172, C1 => A_neg_shifted(44),
                           C2 => n163, ZN => n263);
   U166 : AOI22_X1 port map( A1 => A_neg(44), A2 => n155, B1 => A_signal(44), 
                           B2 => n146, ZN => n264);
   U167 : NAND2_X1 port map( A1 => n280, A2 => n279, ZN => Y(51));
   U168 : AOI22_X1 port map( A1 => A_neg(51), A2 => n155, B1 => A_signal(51), 
                           B2 => n146, ZN => n280);
   U169 : AOI222_X1 port map( A1 => A_shifted(51), A2 => n181, B1 => 
                           zeroSignal(51), B2 => n172, C1 => A_neg_shifted(51),
                           C2 => n162, ZN => n279);
   U170 : NAND2_X1 port map( A1 => n266, A2 => n265, ZN => Y(45));
   U171 : AOI222_X1 port map( A1 => A_shifted(45), A2 => n181, B1 => 
                           zeroSignal(45), B2 => n172, C1 => A_neg_shifted(45),
                           C2 => n163, ZN => n265);
   U172 : AOI22_X1 port map( A1 => A_neg(45), A2 => n155, B1 => A_signal(45), 
                           B2 => n146, ZN => n266);
   U173 : NAND2_X1 port map( A1 => n268, A2 => n267, ZN => Y(46));
   U174 : AOI222_X1 port map( A1 => A_shifted(46), A2 => n181, B1 => 
                           zeroSignal(46), B2 => n172, C1 => A_neg_shifted(46),
                           C2 => n162, ZN => n267);
   U175 : AOI22_X1 port map( A1 => A_neg(46), A2 => n155, B1 => A_signal(46), 
                           B2 => n146, ZN => n268);
   U176 : NAND2_X1 port map( A1 => n284, A2 => n283, ZN => Y(53));
   U177 : AOI222_X1 port map( A1 => A_shifted(53), A2 => n182, B1 => 
                           zeroSignal(53), B2 => n173, C1 => A_neg_shifted(53),
                           C2 => n162, ZN => n283);
   U178 : AOI22_X1 port map( A1 => A_neg(53), A2 => n156, B1 => A_signal(53), 
                           B2 => n147, ZN => n284);
   U179 : NAND2_X1 port map( A1 => n286, A2 => n285, ZN => Y(54));
   U180 : AOI222_X1 port map( A1 => A_shifted(54), A2 => n182, B1 => 
                           zeroSignal(54), B2 => n173, C1 => A_neg_shifted(54),
                           C2 => n162, ZN => n285);
   U181 : NAND2_X1 port map( A1 => n290, A2 => n289, ZN => Y(56));
   U182 : AOI222_X1 port map( A1 => A_shifted(56), A2 => n182, B1 => 
                           zeroSignal(56), B2 => n173, C1 => A_neg_shifted(56),
                           C2 => n162, ZN => n289);
   U183 : NAND2_X1 port map( A1 => n292, A2 => n291, ZN => Y(57));
   U184 : NAND2_X1 port map( A1 => n294, A2 => n293, ZN => Y(58));
   U185 : NAND2_X1 port map( A1 => n282, A2 => n281, ZN => Y(52));
   U186 : AOI22_X1 port map( A1 => A_neg(52), A2 => n155, B1 => A_signal(52), 
                           B2 => n146, ZN => n282);
   U187 : AOI222_X1 port map( A1 => A_shifted(52), A2 => n181, B1 => 
                           zeroSignal(52), B2 => n172, C1 => A_neg_shifted(52),
                           C2 => n162, ZN => n281);
   U188 : NAND2_X1 port map( A1 => n300, A2 => n299, ZN => Y(60));
   U189 : AOI222_X1 port map( A1 => A_shifted(60), A2 => n182, B1 => 
                           zeroSignal(60), B2 => n173, C1 => A_neg_shifted(60),
                           C2 => n161, ZN => n299);
   U190 : NAND2_X1 port map( A1 => n288, A2 => n287, ZN => Y(55));
   U191 : AOI22_X1 port map( A1 => A_neg(55), A2 => n156, B1 => A_signal(55), 
                           B2 => n147, ZN => n288);
   U192 : NAND2_X1 port map( A1 => n304, A2 => n303, ZN => Y(62));
   U193 : AOI222_X1 port map( A1 => A_shifted(62), A2 => n182, B1 => 
                           zeroSignal(62), B2 => n173, C1 => A_neg_shifted(62),
                           C2 => n161, ZN => n303);
   U194 : AOI22_X1 port map( A1 => A_neg(62), A2 => n156, B1 => A_signal(62), 
                           B2 => n147, ZN => n304);
   U195 : NAND2_X1 port map( A1 => n302, A2 => n301, ZN => Y(61));
   U196 : AOI22_X1 port map( A1 => A_neg(61), A2 => n156, B1 => A_signal(61), 
                           B2 => n147, ZN => n302);
   U197 : NAND2_X1 port map( A1 => n296, A2 => n295, ZN => Y(59));
   U198 : AOI22_X1 port map( A1 => A_neg(59), A2 => n156, B1 => A_signal(59), 
                           B2 => n147, ZN => n296);
   U199 : NAND2_X1 port map( A1 => n188, A2 => n187, ZN => Y(0));
   U200 : AOI22_X1 port map( A1 => A_neg(0), A2 => n152, B1 => A_signal(0), B2 
                           => n143, ZN => n188);
   U201 : AOI222_X1 port map( A1 => A_shifted(0), A2 => n178, B1 => 
                           zeroSignal(0), B2 => n169, C1 => A_neg_shifted(0), 
                           C2 => n166, ZN => n187);
   U202 : NAND2_X1 port map( A1 => n210, A2 => n209, ZN => Y(1));
   U203 : AOI22_X1 port map( A1 => A_neg(1), A2 => n152, B1 => A_signal(1), B2 
                           => n143, ZN => n210);
   U204 : AOI222_X1 port map( A1 => A_shifted(1), A2 => n178, B1 => 
                           zeroSignal(1), B2 => n169, C1 => A_neg_shifted(1), 
                           C2 => n165, ZN => n209);
   U205 : NAND2_X1 port map( A1 => n232, A2 => n231, ZN => Y(2));
   U206 : AOI22_X1 port map( A1 => A_neg(2), A2 => n153, B1 => A_signal(2), B2 
                           => n144, ZN => n232);
   U207 : AOI222_X1 port map( A1 => A_shifted(2), A2 => n179, B1 => 
                           zeroSignal(2), B2 => n170, C1 => A_neg_shifted(2), 
                           C2 => n164, ZN => n231);
   U208 : NAND2_X1 port map( A1 => n254, A2 => n253, ZN => Y(3));
   U209 : AOI22_X1 port map( A1 => A_neg(3), A2 => n154, B1 => A_signal(3), B2 
                           => n145, ZN => n254);
   U210 : AOI222_X1 port map( A1 => A_shifted(3), A2 => n180, B1 => 
                           zeroSignal(3), B2 => n171, C1 => A_neg_shifted(3), 
                           C2 => n163, ZN => n253);
   U211 : NAND2_X1 port map( A1 => n276, A2 => n275, ZN => Y(4));
   U212 : AOI22_X1 port map( A1 => A_neg(4), A2 => n155, B1 => A_signal(4), B2 
                           => n146, ZN => n276);
   U213 : AOI222_X1 port map( A1 => A_shifted(4), A2 => n181, B1 => 
                           zeroSignal(4), B2 => n172, C1 => A_neg_shifted(4), 
                           C2 => n162, ZN => n275);
   U214 : NAND2_X1 port map( A1 => n298, A2 => n297, ZN => Y(5));
   U215 : AOI22_X1 port map( A1 => A_neg(5), A2 => n156, B1 => A_signal(5), B2 
                           => n147, ZN => n298);
   U216 : AOI222_X1 port map( A1 => A_shifted(5), A2 => n182, B1 => 
                           zeroSignal(5), B2 => n173, C1 => A_neg_shifted(5), 
                           C2 => n161, ZN => n297);
   U217 : NAND2_X1 port map( A1 => n308, A2 => n307, ZN => Y(6));
   U218 : AOI22_X1 port map( A1 => A_neg(6), A2 => n157, B1 => A_signal(6), B2 
                           => n148, ZN => n308);
   U219 : AOI222_X1 port map( A1 => A_shifted(6), A2 => n183, B1 => 
                           zeroSignal(6), B2 => n174, C1 => A_neg_shifted(6), 
                           C2 => n161, ZN => n307);
   U220 : NAND2_X1 port map( A1 => n310, A2 => n309, ZN => Y(7));
   U221 : AOI22_X1 port map( A1 => A_neg(7), A2 => n157, B1 => A_signal(7), B2 
                           => n148, ZN => n310);
   U222 : AOI222_X1 port map( A1 => A_shifted(7), A2 => n183, B1 => 
                           zeroSignal(7), B2 => n174, C1 => A_neg_shifted(7), 
                           C2 => n161, ZN => n309);
   U223 : NAND2_X1 port map( A1 => n312, A2 => n311, ZN => Y(8));
   U224 : AOI22_X1 port map( A1 => A_neg(8), A2 => n157, B1 => A_signal(8), B2 
                           => n148, ZN => n312);
   U225 : AOI222_X1 port map( A1 => A_shifted(8), A2 => n183, B1 => 
                           zeroSignal(8), B2 => n174, C1 => A_neg_shifted(8), 
                           C2 => n161, ZN => n311);
   U226 : NAND2_X1 port map( A1 => n317, A2 => n316, ZN => Y(9));
   U227 : AOI22_X1 port map( A1 => A_neg(9), A2 => n157, B1 => A_signal(9), B2 
                           => n148, ZN => n317);
   U228 : AOI222_X1 port map( A1 => A_shifted(9), A2 => n183, B1 => 
                           zeroSignal(9), B2 => n174, C1 => A_neg_shifted(9), 
                           C2 => n161, ZN => n316);
   U229 : AOI222_X1 port map( A1 => A_shifted(61), A2 => n182, B1 => 
                           zeroSignal(61), B2 => n173, C1 => A_neg_shifted(61),
                           C2 => n161, ZN => n301);
   U230 : AOI22_X1 port map( A1 => A_neg(60), A2 => n156, B1 => A_signal(60), 
                           B2 => n147, ZN => n300);
   U231 : AOI22_X1 port map( A1 => A_neg(63), A2 => n156, B1 => A_signal(63), 
                           B2 => n147, ZN => n306);
   U232 : AOI222_X1 port map( A1 => A_shifted(59), A2 => n182, B1 => 
                           zeroSignal(59), B2 => n173, C1 => A_neg_shifted(59),
                           C2 => n161, ZN => n295);
   U233 : AOI22_X1 port map( A1 => A_neg(58), A2 => n156, B1 => A_signal(58), 
                           B2 => n147, ZN => n294);
   U234 : AOI222_X1 port map( A1 => A_shifted(57), A2 => n182, B1 => 
                           zeroSignal(57), B2 => n173, C1 => A_neg_shifted(57),
                           C2 => n161, ZN => n291);
   U235 : AOI22_X1 port map( A1 => A_neg(56), A2 => n156, B1 => A_signal(56), 
                           B2 => n147, ZN => n290);
   U236 : AOI222_X1 port map( A1 => A_shifted(58), A2 => n182, B1 => 
                           zeroSignal(58), B2 => n173, C1 => A_neg_shifted(58),
                           C2 => n161, ZN => n293);
   U237 : AOI22_X1 port map( A1 => A_neg(57), A2 => n156, B1 => A_signal(57), 
                           B2 => n147, ZN => n292);
   U238 : AOI222_X1 port map( A1 => A_shifted(55), A2 => n182, B1 => 
                           zeroSignal(55), B2 => n173, C1 => A_neg_shifted(55),
                           C2 => n162, ZN => n287);
   U239 : AOI22_X1 port map( A1 => A_neg(54), A2 => n156, B1 => A_signal(54), 
                           B2 => n147, ZN => n286);
   U240 : AOI222_X1 port map( A1 => A_shifted(11), A2 => n178, B1 => 
                           zeroSignal(11), B2 => n169, C1 => A_neg_shifted(11),
                           C2 => n166, ZN => n191);
   U241 : AOI22_X1 port map( A1 => A_neg(10), A2 => n152, B1 => A_signal(10), 
                           B2 => n143, ZN => n190);
   U242 : NAND2_X1 port map( A1 => n192, A2 => n191, ZN => Y(11));
   U243 : NAND2_X1 port map( A1 => n190, A2 => n189, ZN => Y(10));

end SYN_BEHAVIORAL_2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity MUX51_MuxNbit64_26 is

   port( zeroSignal, A_signal, A_neg, A_shifted, A_neg_shifted : in 
         std_logic_vector (63 downto 0);  Sel : in std_logic_vector (2 downto 
         0);  Y : out std_logic_vector (63 downto 0));

end MUX51_MuxNbit64_26;

architecture SYN_BEHAVIORAL_2 of MUX51_MuxNbit64_26 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, 
      n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, 
      n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, 
      n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, 
      n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, 
      n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, 
      n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, 
      n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, 
      n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, 
      n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, 
      n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, 
      n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, 
      n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, 
      n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, 
      n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, 
      n320 : std_logic;

begin
   
   U1 : AND3_X1 port map( A1 => n319, A2 => n320, A3 => Sel(2), ZN => n141);
   U2 : BUF_X1 port map( A => n141, Z => n166);
   U3 : BUF_X1 port map( A => n185, Z => n184);
   U4 : BUF_X1 port map( A => n159, Z => n158);
   U5 : BUF_X1 port map( A => n150, Z => n149);
   U6 : BUF_X1 port map( A => n141, Z => n167);
   U7 : BUF_X1 port map( A => n185, Z => n183);
   U8 : BUF_X1 port map( A => n159, Z => n157);
   U9 : BUF_X1 port map( A => n150, Z => n148);
   U10 : BUF_X1 port map( A => n176, Z => n175);
   U11 : BUF_X1 port map( A => n176, Z => n174);
   U12 : BUF_X1 port map( A => n158, Z => n151);
   U13 : BUF_X1 port map( A => n184, Z => n177);
   U14 : BUF_X1 port map( A => n149, Z => n142);
   U15 : BUF_X1 port map( A => n166, Z => n164);
   U16 : BUF_X1 port map( A => n184, Z => n178);
   U17 : BUF_X1 port map( A => n158, Z => n152);
   U18 : BUF_X1 port map( A => n149, Z => n143);
   U19 : BUF_X1 port map( A => n166, Z => n163);
   U20 : BUF_X1 port map( A => n184, Z => n179);
   U21 : BUF_X1 port map( A => n158, Z => n153);
   U22 : BUF_X1 port map( A => n149, Z => n144);
   U23 : BUF_X1 port map( A => n167, Z => n162);
   U24 : BUF_X1 port map( A => n183, Z => n180);
   U25 : BUF_X1 port map( A => n157, Z => n154);
   U26 : BUF_X1 port map( A => n148, Z => n145);
   U27 : BUF_X1 port map( A => n167, Z => n161);
   U28 : BUF_X1 port map( A => n157, Z => n155);
   U29 : BUF_X1 port map( A => n183, Z => n181);
   U30 : BUF_X1 port map( A => n148, Z => n146);
   U31 : BUF_X1 port map( A => n167, Z => n160);
   U32 : BUF_X1 port map( A => n175, Z => n169);
   U33 : BUF_X1 port map( A => n175, Z => n170);
   U34 : BUF_X1 port map( A => n174, Z => n171);
   U35 : BUF_X1 port map( A => n175, Z => n168);
   U36 : BUF_X1 port map( A => n174, Z => n172);
   U37 : BUF_X1 port map( A => n166, Z => n165);
   U38 : BUF_X1 port map( A => n157, Z => n156);
   U39 : BUF_X1 port map( A => n148, Z => n147);
   U40 : BUF_X1 port map( A => n174, Z => n173);
   U41 : BUF_X1 port map( A => n183, Z => n182);
   U42 : INV_X1 port map( A => Sel(1), ZN => n320);
   U43 : BUF_X1 port map( A => n314, Z => n159);
   U44 : NOR3_X1 port map( A1 => Sel(0), A2 => Sel(2), A3 => n320, ZN => n314);
   U45 : BUF_X1 port map( A => n316, Z => n185);
   U46 : NOR3_X1 port map( A1 => n319, A2 => Sel(2), A3 => n320, ZN => n316);
   U47 : INV_X1 port map( A => Sel(0), ZN => n319);
   U48 : BUF_X1 port map( A => n313, Z => n150);
   U49 : NOR3_X1 port map( A1 => Sel(1), A2 => Sel(2), A3 => n319, ZN => n313);
   U50 : BUF_X1 port map( A => n315, Z => n176);
   U51 : NOR2_X1 port map( A1 => n165, A2 => n186, ZN => n315);
   U52 : AOI21_X1 port map( B1 => n319, B2 => n320, A => Sel(2), ZN => n186);
   U53 : AOI22_X1 port map( A1 => A_neg(13), A2 => n151, B1 => A_signal(13), B2
                           => n142, ZN => n196);
   U54 : AOI222_X1 port map( A1 => A_shifted(12), A2 => n177, B1 => 
                           zeroSignal(12), B2 => n168, C1 => A_neg_shifted(12),
                           C2 => n165, ZN => n193);
   U55 : NAND2_X1 port map( A1 => n198, A2 => n197, ZN => Y(14));
   U56 : AOI22_X1 port map( A1 => A_neg(14), A2 => n151, B1 => A_signal(14), B2
                           => n142, ZN => n198);
   U57 : AOI222_X1 port map( A1 => A_shifted(14), A2 => n177, B1 => 
                           zeroSignal(14), B2 => n168, C1 => A_neg_shifted(14),
                           C2 => n164, ZN => n197);
   U58 : NAND2_X1 port map( A1 => n200, A2 => n199, ZN => Y(15));
   U59 : AOI22_X1 port map( A1 => A_neg(15), A2 => n151, B1 => A_signal(15), B2
                           => n142, ZN => n200);
   U60 : AOI222_X1 port map( A1 => A_shifted(15), A2 => n177, B1 => 
                           zeroSignal(15), B2 => n168, C1 => A_neg_shifted(15),
                           C2 => n164, ZN => n199);
   U61 : NAND2_X1 port map( A1 => n202, A2 => n201, ZN => Y(16));
   U62 : AOI22_X1 port map( A1 => A_neg(16), A2 => n151, B1 => A_signal(16), B2
                           => n142, ZN => n202);
   U63 : AOI222_X1 port map( A1 => A_shifted(16), A2 => n177, B1 => 
                           zeroSignal(16), B2 => n168, C1 => A_neg_shifted(16),
                           C2 => n164, ZN => n201);
   U64 : NAND2_X1 port map( A1 => n204, A2 => n203, ZN => Y(17));
   U65 : AOI22_X1 port map( A1 => A_neg(17), A2 => n151, B1 => A_signal(17), B2
                           => n142, ZN => n204);
   U66 : AOI222_X1 port map( A1 => A_shifted(17), A2 => n177, B1 => 
                           zeroSignal(17), B2 => n168, C1 => A_neg_shifted(17),
                           C2 => n164, ZN => n203);
   U67 : NAND2_X1 port map( A1 => n206, A2 => n205, ZN => Y(18));
   U68 : AOI22_X1 port map( A1 => A_neg(18), A2 => n151, B1 => A_signal(18), B2
                           => n142, ZN => n206);
   U69 : AOI222_X1 port map( A1 => A_shifted(18), A2 => n177, B1 => 
                           zeroSignal(18), B2 => n168, C1 => A_neg_shifted(18),
                           C2 => n164, ZN => n205);
   U70 : NAND2_X1 port map( A1 => n208, A2 => n207, ZN => Y(19));
   U71 : AOI22_X1 port map( A1 => A_neg(19), A2 => n151, B1 => A_signal(19), B2
                           => n142, ZN => n208);
   U72 : AOI222_X1 port map( A1 => A_shifted(19), A2 => n177, B1 => 
                           zeroSignal(19), B2 => n168, C1 => A_neg_shifted(19),
                           C2 => n164, ZN => n207);
   U73 : NAND2_X1 port map( A1 => n270, A2 => n269, ZN => Y(47));
   U74 : AOI222_X1 port map( A1 => A_shifted(47), A2 => n180, B1 => 
                           zeroSignal(47), B2 => n171, C1 => A_neg_shifted(47),
                           C2 => n161, ZN => n269);
   U75 : AOI22_X1 port map( A1 => A_neg(47), A2 => n154, B1 => A_signal(47), B2
                           => n145, ZN => n270);
   U76 : NAND2_X1 port map( A1 => n216, A2 => n215, ZN => Y(22));
   U77 : AOI222_X1 port map( A1 => A_shifted(22), A2 => n178, B1 => 
                           zeroSignal(22), B2 => n169, C1 => A_neg_shifted(22),
                           C2 => n164, ZN => n215);
   U78 : AOI22_X1 port map( A1 => A_neg(22), A2 => n152, B1 => A_signal(22), B2
                           => n143, ZN => n216);
   U79 : NAND2_X1 port map( A1 => n218, A2 => n217, ZN => Y(23));
   U80 : AOI222_X1 port map( A1 => A_shifted(23), A2 => n178, B1 => 
                           zeroSignal(23), B2 => n169, C1 => A_neg_shifted(23),
                           C2 => n164, ZN => n217);
   U81 : AOI22_X1 port map( A1 => A_neg(23), A2 => n152, B1 => A_signal(23), B2
                           => n143, ZN => n218);
   U82 : NAND2_X1 port map( A1 => n220, A2 => n219, ZN => Y(24));
   U83 : AOI222_X1 port map( A1 => A_shifted(24), A2 => n178, B1 => 
                           zeroSignal(24), B2 => n169, C1 => A_neg_shifted(24),
                           C2 => n163, ZN => n219);
   U84 : AOI22_X1 port map( A1 => A_neg(24), A2 => n152, B1 => A_signal(24), B2
                           => n143, ZN => n220);
   U85 : NAND2_X1 port map( A1 => n272, A2 => n271, ZN => Y(48));
   U86 : AOI222_X1 port map( A1 => A_shifted(48), A2 => n180, B1 => 
                           zeroSignal(48), B2 => n171, C1 => A_neg_shifted(48),
                           C2 => n161, ZN => n271);
   U87 : AOI22_X1 port map( A1 => A_neg(48), A2 => n154, B1 => A_signal(48), B2
                           => n145, ZN => n272);
   U88 : NAND2_X1 port map( A1 => n222, A2 => n221, ZN => Y(25));
   U89 : AOI222_X1 port map( A1 => A_shifted(25), A2 => n178, B1 => 
                           zeroSignal(25), B2 => n169, C1 => A_neg_shifted(25),
                           C2 => n163, ZN => n221);
   U90 : AOI22_X1 port map( A1 => A_neg(25), A2 => n152, B1 => A_signal(25), B2
                           => n143, ZN => n222);
   U91 : NAND2_X1 port map( A1 => n226, A2 => n225, ZN => Y(27));
   U92 : AOI222_X1 port map( A1 => A_shifted(27), A2 => n178, B1 => 
                           zeroSignal(27), B2 => n169, C1 => A_neg_shifted(27),
                           C2 => n163, ZN => n225);
   U93 : AOI22_X1 port map( A1 => A_neg(27), A2 => n152, B1 => A_signal(27), B2
                           => n143, ZN => n226);
   U94 : NAND2_X1 port map( A1 => n228, A2 => n227, ZN => Y(28));
   U95 : AOI222_X1 port map( A1 => A_shifted(28), A2 => n178, B1 => 
                           zeroSignal(28), B2 => n169, C1 => A_neg_shifted(28),
                           C2 => n163, ZN => n227);
   U96 : AOI22_X1 port map( A1 => A_neg(28), A2 => n152, B1 => A_signal(28), B2
                           => n143, ZN => n228);
   U97 : NAND2_X1 port map( A1 => n274, A2 => n273, ZN => Y(49));
   U98 : AOI22_X1 port map( A1 => A_neg(49), A2 => n154, B1 => A_signal(49), B2
                           => n145, ZN => n274);
   U99 : AOI222_X1 port map( A1 => A_shifted(49), A2 => n180, B1 => 
                           zeroSignal(49), B2 => n171, C1 => A_neg_shifted(49),
                           C2 => n161, ZN => n273);
   U100 : NAND2_X1 port map( A1 => n224, A2 => n223, ZN => Y(26));
   U101 : AOI22_X1 port map( A1 => A_neg(26), A2 => n152, B1 => A_signal(26), 
                           B2 => n143, ZN => n224);
   U102 : AOI222_X1 port map( A1 => A_shifted(26), A2 => n178, B1 => 
                           zeroSignal(26), B2 => n169, C1 => A_neg_shifted(26),
                           C2 => n163, ZN => n223);
   U103 : NAND2_X1 port map( A1 => n230, A2 => n229, ZN => Y(29));
   U104 : AOI222_X1 port map( A1 => A_shifted(29), A2 => n178, B1 => 
                           zeroSignal(29), B2 => n169, C1 => A_neg_shifted(29),
                           C2 => n163, ZN => n229);
   U105 : AOI22_X1 port map( A1 => A_neg(29), A2 => n152, B1 => A_signal(29), 
                           B2 => n143, ZN => n230);
   U106 : NAND2_X1 port map( A1 => n212, A2 => n211, ZN => Y(20));
   U107 : AOI22_X1 port map( A1 => A_neg(20), A2 => n152, B1 => A_signal(20), 
                           B2 => n143, ZN => n212);
   U108 : AOI222_X1 port map( A1 => A_shifted(20), A2 => n178, B1 => 
                           zeroSignal(20), B2 => n169, C1 => A_neg_shifted(20),
                           C2 => n164, ZN => n211);
   U109 : NAND2_X1 port map( A1 => n236, A2 => n235, ZN => Y(31));
   U110 : AOI222_X1 port map( A1 => A_shifted(31), A2 => n179, B1 => 
                           zeroSignal(31), B2 => n170, C1 => A_neg_shifted(31),
                           C2 => n163, ZN => n235);
   U111 : AOI22_X1 port map( A1 => A_neg(31), A2 => n153, B1 => A_signal(31), 
                           B2 => n144, ZN => n236);
   U112 : NAND2_X1 port map( A1 => n238, A2 => n237, ZN => Y(32));
   U113 : AOI222_X1 port map( A1 => A_shifted(32), A2 => n179, B1 => 
                           zeroSignal(32), B2 => n170, C1 => A_neg_shifted(32),
                           C2 => n163, ZN => n237);
   U114 : AOI22_X1 port map( A1 => A_neg(32), A2 => n153, B1 => A_signal(32), 
                           B2 => n144, ZN => n238);
   U115 : NAND2_X1 port map( A1 => n240, A2 => n239, ZN => Y(33));
   U116 : AOI222_X1 port map( A1 => A_shifted(33), A2 => n179, B1 => 
                           zeroSignal(33), B2 => n170, C1 => A_neg_shifted(33),
                           C2 => n163, ZN => n239);
   U117 : AOI22_X1 port map( A1 => A_neg(33), A2 => n153, B1 => A_signal(33), 
                           B2 => n144, ZN => n240);
   U118 : NAND2_X1 port map( A1 => n244, A2 => n243, ZN => Y(35));
   U119 : AOI222_X1 port map( A1 => A_shifted(35), A2 => n179, B1 => 
                           zeroSignal(35), B2 => n170, C1 => A_neg_shifted(35),
                           C2 => n162, ZN => n243);
   U120 : AOI22_X1 port map( A1 => A_neg(35), A2 => n153, B1 => A_signal(35), 
                           B2 => n144, ZN => n244);
   U121 : NAND2_X1 port map( A1 => n242, A2 => n241, ZN => Y(34));
   U122 : AOI222_X1 port map( A1 => A_shifted(34), A2 => n179, B1 => 
                           zeroSignal(34), B2 => n170, C1 => A_neg_shifted(34),
                           C2 => n163, ZN => n241);
   U123 : AOI22_X1 port map( A1 => A_neg(34), A2 => n153, B1 => A_signal(34), 
                           B2 => n144, ZN => n242);
   U124 : NAND2_X1 port map( A1 => n234, A2 => n233, ZN => Y(30));
   U125 : AOI22_X1 port map( A1 => A_neg(30), A2 => n152, B1 => A_signal(30), 
                           B2 => n143, ZN => n234);
   U126 : AOI222_X1 port map( A1 => A_shifted(30), A2 => n178, B1 => 
                           zeroSignal(30), B2 => n169, C1 => A_neg_shifted(30),
                           C2 => n163, ZN => n233);
   U127 : NAND2_X1 port map( A1 => n248, A2 => n247, ZN => Y(37));
   U128 : AOI222_X1 port map( A1 => A_shifted(37), A2 => n179, B1 => 
                           zeroSignal(37), B2 => n170, C1 => A_neg_shifted(37),
                           C2 => n162, ZN => n247);
   U129 : AOI22_X1 port map( A1 => A_neg(37), A2 => n153, B1 => A_signal(37), 
                           B2 => n144, ZN => n248);
   U130 : NAND2_X1 port map( A1 => n252, A2 => n251, ZN => Y(39));
   U131 : AOI222_X1 port map( A1 => A_shifted(39), A2 => n179, B1 => 
                           zeroSignal(39), B2 => n170, C1 => A_neg_shifted(39),
                           C2 => n162, ZN => n251);
   U132 : AOI22_X1 port map( A1 => A_neg(39), A2 => n153, B1 => A_signal(39), 
                           B2 => n144, ZN => n252);
   U133 : NAND2_X1 port map( A1 => n250, A2 => n249, ZN => Y(38));
   U134 : AOI222_X1 port map( A1 => A_shifted(38), A2 => n179, B1 => 
                           zeroSignal(38), B2 => n170, C1 => A_neg_shifted(38),
                           C2 => n162, ZN => n249);
   U135 : AOI22_X1 port map( A1 => A_neg(38), A2 => n153, B1 => A_signal(38), 
                           B2 => n144, ZN => n250);
   U136 : NAND2_X1 port map( A1 => n246, A2 => n245, ZN => Y(36));
   U137 : AOI22_X1 port map( A1 => A_neg(36), A2 => n153, B1 => A_signal(36), 
                           B2 => n144, ZN => n246);
   U138 : AOI222_X1 port map( A1 => A_shifted(36), A2 => n179, B1 => 
                           zeroSignal(36), B2 => n170, C1 => A_neg_shifted(36),
                           C2 => n162, ZN => n245);
   U139 : NAND2_X1 port map( A1 => n256, A2 => n255, ZN => Y(40));
   U140 : AOI222_X1 port map( A1 => A_shifted(40), A2 => n179, B1 => 
                           zeroSignal(40), B2 => n170, C1 => A_neg_shifted(40),
                           C2 => n162, ZN => n255);
   U141 : AOI22_X1 port map( A1 => A_neg(40), A2 => n153, B1 => A_signal(40), 
                           B2 => n144, ZN => n256);
   U142 : NAND2_X1 port map( A1 => n266, A2 => n265, ZN => Y(45));
   U143 : AOI222_X1 port map( A1 => A_shifted(45), A2 => n180, B1 => 
                           zeroSignal(45), B2 => n171, C1 => A_neg_shifted(45),
                           C2 => n162, ZN => n265);
   U144 : AOI22_X1 port map( A1 => A_neg(45), A2 => n154, B1 => A_signal(45), 
                           B2 => n145, ZN => n266);
   U145 : NAND2_X1 port map( A1 => n214, A2 => n213, ZN => Y(21));
   U146 : AOI222_X1 port map( A1 => A_shifted(21), A2 => n178, B1 => 
                           zeroSignal(21), B2 => n169, C1 => A_neg_shifted(21),
                           C2 => n164, ZN => n213);
   U147 : AOI22_X1 port map( A1 => A_neg(21), A2 => n152, B1 => A_signal(21), 
                           B2 => n143, ZN => n214);
   U148 : NAND2_X1 port map( A1 => n258, A2 => n257, ZN => Y(41));
   U149 : AOI222_X1 port map( A1 => A_shifted(41), A2 => n179, B1 => 
                           zeroSignal(41), B2 => n170, C1 => A_neg_shifted(41),
                           C2 => n162, ZN => n257);
   U150 : AOI22_X1 port map( A1 => A_neg(41), A2 => n153, B1 => A_signal(41), 
                           B2 => n144, ZN => n258);
   U151 : NAND2_X1 port map( A1 => n260, A2 => n259, ZN => Y(42));
   U152 : AOI222_X1 port map( A1 => A_shifted(42), A2 => n180, B1 => 
                           zeroSignal(42), B2 => n171, C1 => A_neg_shifted(42),
                           C2 => n162, ZN => n259);
   U153 : AOI22_X1 port map( A1 => A_neg(42), A2 => n154, B1 => A_signal(42), 
                           B2 => n145, ZN => n260);
   U154 : NAND2_X1 port map( A1 => n264, A2 => n263, ZN => Y(44));
   U155 : AOI222_X1 port map( A1 => A_shifted(44), A2 => n180, B1 => 
                           zeroSignal(44), B2 => n171, C1 => A_neg_shifted(44),
                           C2 => n162, ZN => n263);
   U156 : AOI22_X1 port map( A1 => A_neg(44), A2 => n154, B1 => A_signal(44), 
                           B2 => n145, ZN => n264);
   U157 : NAND2_X1 port map( A1 => n262, A2 => n261, ZN => Y(43));
   U158 : AOI222_X1 port map( A1 => A_shifted(43), A2 => n180, B1 => 
                           zeroSignal(43), B2 => n171, C1 => A_neg_shifted(43),
                           C2 => n162, ZN => n261);
   U159 : AOI22_X1 port map( A1 => A_neg(43), A2 => n154, B1 => A_signal(43), 
                           B2 => n145, ZN => n262);
   U160 : NAND2_X1 port map( A1 => n282, A2 => n281, ZN => Y(52));
   U161 : AOI222_X1 port map( A1 => A_shifted(52), A2 => n180, B1 => 
                           zeroSignal(52), B2 => n171, C1 => A_neg_shifted(52),
                           C2 => n161, ZN => n281);
   U162 : AOI22_X1 port map( A1 => A_neg(52), A2 => n154, B1 => A_signal(52), 
                           B2 => n145, ZN => n282);
   U163 : NAND2_X1 port map( A1 => n280, A2 => n279, ZN => Y(51));
   U164 : AOI222_X1 port map( A1 => A_shifted(51), A2 => n180, B1 => 
                           zeroSignal(51), B2 => n171, C1 => A_neg_shifted(51),
                           C2 => n161, ZN => n279);
   U165 : AOI22_X1 port map( A1 => A_neg(51), A2 => n154, B1 => A_signal(51), 
                           B2 => n145, ZN => n280);
   U166 : NAND2_X1 port map( A1 => n278, A2 => n277, ZN => Y(50));
   U167 : AOI222_X1 port map( A1 => A_shifted(50), A2 => n180, B1 => 
                           zeroSignal(50), B2 => n171, C1 => A_neg_shifted(50),
                           C2 => n161, ZN => n277);
   U168 : AOI22_X1 port map( A1 => A_neg(50), A2 => n154, B1 => A_signal(50), 
                           B2 => n145, ZN => n278);
   U169 : NAND2_X1 port map( A1 => n268, A2 => n267, ZN => Y(46));
   U170 : AOI22_X1 port map( A1 => A_neg(46), A2 => n154, B1 => A_signal(46), 
                           B2 => n145, ZN => n268);
   U171 : AOI222_X1 port map( A1 => A_shifted(46), A2 => n180, B1 => 
                           zeroSignal(46), B2 => n171, C1 => A_neg_shifted(46),
                           C2 => n161, ZN => n267);
   U172 : NAND2_X1 port map( A1 => n284, A2 => n283, ZN => Y(53));
   U173 : AOI22_X1 port map( A1 => A_neg(53), A2 => n155, B1 => A_signal(53), 
                           B2 => n146, ZN => n284);
   U174 : AOI222_X1 port map( A1 => A_shifted(53), A2 => n181, B1 => 
                           zeroSignal(53), B2 => n172, C1 => A_neg_shifted(53),
                           C2 => n161, ZN => n283);
   U175 : NAND2_X1 port map( A1 => n304, A2 => n303, ZN => Y(62));
   U176 : AOI222_X1 port map( A1 => A_shifted(62), A2 => n181, B1 => 
                           zeroSignal(62), B2 => n172, C1 => A_neg_shifted(62),
                           C2 => n160, ZN => n303);
   U177 : NAND2_X1 port map( A1 => n296, A2 => n295, ZN => Y(59));
   U178 : NAND2_X1 port map( A1 => n290, A2 => n289, ZN => Y(56));
   U179 : AOI222_X1 port map( A1 => A_shifted(56), A2 => n181, B1 => 
                           zeroSignal(56), B2 => n172, C1 => A_neg_shifted(56),
                           C2 => n161, ZN => n289);
   U180 : NAND2_X1 port map( A1 => n288, A2 => n287, ZN => Y(55));
   U181 : AOI222_X1 port map( A1 => A_shifted(55), A2 => n181, B1 => 
                           zeroSignal(55), B2 => n172, C1 => A_neg_shifted(55),
                           C2 => n161, ZN => n287);
   U182 : AOI22_X1 port map( A1 => A_neg(55), A2 => n155, B1 => A_signal(55), 
                           B2 => n146, ZN => n288);
   U183 : NAND2_X1 port map( A1 => n294, A2 => n293, ZN => Y(58));
   U184 : AOI222_X1 port map( A1 => A_shifted(58), A2 => n181, B1 => 
                           zeroSignal(58), B2 => n172, C1 => A_neg_shifted(58),
                           C2 => n160, ZN => n293);
   U185 : NAND2_X1 port map( A1 => n300, A2 => n299, ZN => Y(60));
   U186 : NAND2_X1 port map( A1 => n292, A2 => n291, ZN => Y(57));
   U187 : AOI22_X1 port map( A1 => A_neg(57), A2 => n155, B1 => A_signal(57), 
                           B2 => n146, ZN => n292);
   U188 : NAND2_X1 port map( A1 => n286, A2 => n285, ZN => Y(54));
   U189 : AOI22_X1 port map( A1 => A_neg(54), A2 => n155, B1 => A_signal(54), 
                           B2 => n146, ZN => n286);
   U190 : AOI222_X1 port map( A1 => A_shifted(54), A2 => n181, B1 => 
                           zeroSignal(54), B2 => n172, C1 => A_neg_shifted(54),
                           C2 => n161, ZN => n285);
   U191 : NAND2_X1 port map( A1 => n306, A2 => n305, ZN => Y(63));
   U192 : AOI22_X1 port map( A1 => A_neg(63), A2 => n155, B1 => A_signal(63), 
                           B2 => n146, ZN => n306);
   U193 : NAND2_X1 port map( A1 => n302, A2 => n301, ZN => Y(61));
   U194 : AOI22_X1 port map( A1 => A_neg(61), A2 => n155, B1 => A_signal(61), 
                           B2 => n146, ZN => n302);
   U195 : NAND2_X1 port map( A1 => n188, A2 => n187, ZN => Y(0));
   U196 : AOI22_X1 port map( A1 => A_neg(0), A2 => n151, B1 => A_signal(0), B2 
                           => n142, ZN => n188);
   U197 : AOI222_X1 port map( A1 => A_shifted(0), A2 => n177, B1 => 
                           zeroSignal(0), B2 => n168, C1 => A_neg_shifted(0), 
                           C2 => n165, ZN => n187);
   U198 : NAND2_X1 port map( A1 => n210, A2 => n209, ZN => Y(1));
   U199 : AOI22_X1 port map( A1 => A_neg(1), A2 => n151, B1 => A_signal(1), B2 
                           => n142, ZN => n210);
   U200 : AOI222_X1 port map( A1 => A_shifted(1), A2 => n177, B1 => 
                           zeroSignal(1), B2 => n168, C1 => A_neg_shifted(1), 
                           C2 => n164, ZN => n209);
   U201 : NAND2_X1 port map( A1 => n232, A2 => n231, ZN => Y(2));
   U202 : AOI22_X1 port map( A1 => A_neg(2), A2 => n152, B1 => A_signal(2), B2 
                           => n143, ZN => n232);
   U203 : AOI222_X1 port map( A1 => A_shifted(2), A2 => n178, B1 => 
                           zeroSignal(2), B2 => n169, C1 => A_neg_shifted(2), 
                           C2 => n163, ZN => n231);
   U204 : NAND2_X1 port map( A1 => n254, A2 => n253, ZN => Y(3));
   U205 : AOI22_X1 port map( A1 => A_neg(3), A2 => n153, B1 => A_signal(3), B2 
                           => n144, ZN => n254);
   U206 : AOI222_X1 port map( A1 => A_shifted(3), A2 => n179, B1 => 
                           zeroSignal(3), B2 => n170, C1 => A_neg_shifted(3), 
                           C2 => n162, ZN => n253);
   U207 : NAND2_X1 port map( A1 => n276, A2 => n275, ZN => Y(4));
   U208 : AOI22_X1 port map( A1 => A_neg(4), A2 => n154, B1 => A_signal(4), B2 
                           => n145, ZN => n276);
   U209 : AOI222_X1 port map( A1 => A_shifted(4), A2 => n180, B1 => 
                           zeroSignal(4), B2 => n171, C1 => A_neg_shifted(4), 
                           C2 => n161, ZN => n275);
   U210 : NAND2_X1 port map( A1 => n298, A2 => n297, ZN => Y(5));
   U211 : AOI22_X1 port map( A1 => A_neg(5), A2 => n155, B1 => A_signal(5), B2 
                           => n146, ZN => n298);
   U212 : AOI222_X1 port map( A1 => A_shifted(5), A2 => n181, B1 => 
                           zeroSignal(5), B2 => n172, C1 => A_neg_shifted(5), 
                           C2 => n160, ZN => n297);
   U213 : NAND2_X1 port map( A1 => n308, A2 => n307, ZN => Y(6));
   U214 : AOI22_X1 port map( A1 => A_neg(6), A2 => n156, B1 => A_signal(6), B2 
                           => n147, ZN => n308);
   U215 : AOI222_X1 port map( A1 => A_shifted(6), A2 => n182, B1 => 
                           zeroSignal(6), B2 => n173, C1 => A_neg_shifted(6), 
                           C2 => n160, ZN => n307);
   U216 : NAND2_X1 port map( A1 => n310, A2 => n309, ZN => Y(7));
   U217 : AOI22_X1 port map( A1 => A_neg(7), A2 => n156, B1 => A_signal(7), B2 
                           => n147, ZN => n310);
   U218 : AOI222_X1 port map( A1 => A_shifted(7), A2 => n182, B1 => 
                           zeroSignal(7), B2 => n173, C1 => A_neg_shifted(7), 
                           C2 => n160, ZN => n309);
   U219 : NAND2_X1 port map( A1 => n312, A2 => n311, ZN => Y(8));
   U220 : AOI22_X1 port map( A1 => A_neg(8), A2 => n156, B1 => A_signal(8), B2 
                           => n147, ZN => n312);
   U221 : AOI222_X1 port map( A1 => A_shifted(8), A2 => n182, B1 => 
                           zeroSignal(8), B2 => n173, C1 => A_neg_shifted(8), 
                           C2 => n160, ZN => n311);
   U222 : NAND2_X1 port map( A1 => n318, A2 => n317, ZN => Y(9));
   U223 : AOI22_X1 port map( A1 => A_neg(9), A2 => n156, B1 => A_signal(9), B2 
                           => n147, ZN => n318);
   U224 : AOI222_X1 port map( A1 => A_shifted(9), A2 => n182, B1 => 
                           zeroSignal(9), B2 => n173, C1 => A_neg_shifted(9), 
                           C2 => n160, ZN => n317);
   U225 : NAND2_X1 port map( A1 => n190, A2 => n189, ZN => Y(10));
   U226 : AOI22_X1 port map( A1 => A_neg(10), A2 => n151, B1 => A_signal(10), 
                           B2 => n142, ZN => n190);
   U227 : AOI222_X1 port map( A1 => A_shifted(10), A2 => n177, B1 => 
                           zeroSignal(10), B2 => n168, C1 => A_neg_shifted(10),
                           C2 => n165, ZN => n189);
   U228 : NAND2_X1 port map( A1 => n192, A2 => n191, ZN => Y(11));
   U229 : AOI22_X1 port map( A1 => A_neg(11), A2 => n151, B1 => A_signal(11), 
                           B2 => n142, ZN => n192);
   U230 : AOI222_X1 port map( A1 => A_shifted(11), A2 => n177, B1 => 
                           zeroSignal(11), B2 => n168, C1 => A_neg_shifted(11),
                           C2 => n165, ZN => n191);
   U231 : AOI222_X1 port map( A1 => A_shifted(63), A2 => n181, B1 => 
                           zeroSignal(63), B2 => n172, C1 => A_neg_shifted(63),
                           C2 => n160, ZN => n305);
   U232 : AOI22_X1 port map( A1 => A_neg(62), A2 => n155, B1 => A_signal(62), 
                           B2 => n146, ZN => n304);
   U233 : AOI222_X1 port map( A1 => A_shifted(61), A2 => n181, B1 => 
                           zeroSignal(61), B2 => n172, C1 => A_neg_shifted(61),
                           C2 => n160, ZN => n301);
   U234 : AOI22_X1 port map( A1 => A_neg(60), A2 => n155, B1 => A_signal(60), 
                           B2 => n146, ZN => n300);
   U235 : AOI222_X1 port map( A1 => A_shifted(59), A2 => n181, B1 => 
                           zeroSignal(59), B2 => n172, C1 => A_neg_shifted(59),
                           C2 => n160, ZN => n295);
   U236 : AOI22_X1 port map( A1 => A_neg(58), A2 => n155, B1 => A_signal(58), 
                           B2 => n146, ZN => n294);
   U237 : AOI222_X1 port map( A1 => A_shifted(60), A2 => n181, B1 => 
                           zeroSignal(60), B2 => n172, C1 => A_neg_shifted(60),
                           C2 => n160, ZN => n299);
   U238 : AOI22_X1 port map( A1 => A_neg(59), A2 => n155, B1 => A_signal(59), 
                           B2 => n146, ZN => n296);
   U239 : AOI222_X1 port map( A1 => A_shifted(57), A2 => n181, B1 => 
                           zeroSignal(57), B2 => n172, C1 => A_neg_shifted(57),
                           C2 => n160, ZN => n291);
   U240 : AOI22_X1 port map( A1 => A_neg(56), A2 => n155, B1 => A_signal(56), 
                           B2 => n146, ZN => n290);
   U241 : AOI222_X1 port map( A1 => A_shifted(13), A2 => n177, B1 => 
                           zeroSignal(13), B2 => n168, C1 => A_neg_shifted(13),
                           C2 => n164, ZN => n195);
   U242 : AOI22_X1 port map( A1 => A_neg(12), A2 => n151, B1 => A_signal(12), 
                           B2 => n142, ZN => n194);
   U243 : NAND2_X1 port map( A1 => n196, A2 => n195, ZN => Y(13));
   U244 : NAND2_X1 port map( A1 => n194, A2 => n193, ZN => Y(12));

end SYN_BEHAVIORAL_2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity MUX51_MuxNbit64_25 is

   port( zeroSignal, A_signal, A_neg, A_shifted, A_neg_shifted : in 
         std_logic_vector (63 downto 0);  Sel : in std_logic_vector (2 downto 
         0);  Y : out std_logic_vector (63 downto 0));

end MUX51_MuxNbit64_25;

architecture SYN_BEHAVIORAL_2 of MUX51_MuxNbit64_25 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, 
      n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, 
      n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, 
      n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, 
      n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, 
      n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, 
      n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, 
      n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, 
      n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, 
      n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, 
      n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, 
      n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, 
      n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, 
      n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, 
      n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, 
      n320 : std_logic;

begin
   
   U1 : AND3_X1 port map( A1 => n319, A2 => n320, A3 => Sel(2), ZN => n141);
   U2 : BUF_X1 port map( A => n141, Z => n166);
   U3 : BUF_X1 port map( A => n185, Z => n184);
   U4 : BUF_X1 port map( A => n159, Z => n158);
   U5 : BUF_X1 port map( A => n150, Z => n149);
   U6 : BUF_X1 port map( A => n141, Z => n167);
   U7 : BUF_X1 port map( A => n185, Z => n183);
   U8 : BUF_X1 port map( A => n159, Z => n157);
   U9 : BUF_X1 port map( A => n150, Z => n148);
   U10 : BUF_X1 port map( A => n176, Z => n175);
   U11 : BUF_X1 port map( A => n176, Z => n174);
   U12 : BUF_X1 port map( A => n158, Z => n151);
   U13 : BUF_X1 port map( A => n184, Z => n177);
   U14 : BUF_X1 port map( A => n149, Z => n142);
   U15 : BUF_X1 port map( A => n166, Z => n164);
   U16 : BUF_X1 port map( A => n184, Z => n178);
   U17 : BUF_X1 port map( A => n158, Z => n152);
   U18 : BUF_X1 port map( A => n149, Z => n143);
   U19 : BUF_X1 port map( A => n166, Z => n163);
   U20 : BUF_X1 port map( A => n184, Z => n179);
   U21 : BUF_X1 port map( A => n158, Z => n153);
   U22 : BUF_X1 port map( A => n149, Z => n144);
   U23 : BUF_X1 port map( A => n167, Z => n162);
   U24 : BUF_X1 port map( A => n183, Z => n180);
   U25 : BUF_X1 port map( A => n157, Z => n154);
   U26 : BUF_X1 port map( A => n148, Z => n145);
   U27 : BUF_X1 port map( A => n167, Z => n161);
   U28 : BUF_X1 port map( A => n183, Z => n181);
   U29 : BUF_X1 port map( A => n157, Z => n155);
   U30 : BUF_X1 port map( A => n148, Z => n146);
   U31 : BUF_X1 port map( A => n167, Z => n160);
   U32 : BUF_X1 port map( A => n175, Z => n169);
   U33 : BUF_X1 port map( A => n175, Z => n170);
   U34 : BUF_X1 port map( A => n174, Z => n171);
   U35 : BUF_X1 port map( A => n175, Z => n168);
   U36 : BUF_X1 port map( A => n174, Z => n172);
   U37 : BUF_X1 port map( A => n166, Z => n165);
   U38 : BUF_X1 port map( A => n157, Z => n156);
   U39 : BUF_X1 port map( A => n148, Z => n147);
   U40 : BUF_X1 port map( A => n174, Z => n173);
   U41 : BUF_X1 port map( A => n183, Z => n182);
   U42 : BUF_X1 port map( A => n314, Z => n159);
   U43 : NOR3_X1 port map( A1 => Sel(0), A2 => Sel(2), A3 => n320, ZN => n314);
   U44 : INV_X1 port map( A => Sel(1), ZN => n320);
   U45 : BUF_X1 port map( A => n316, Z => n185);
   U46 : NOR3_X1 port map( A1 => n319, A2 => Sel(2), A3 => n320, ZN => n316);
   U47 : BUF_X1 port map( A => n313, Z => n150);
   U48 : NOR3_X1 port map( A1 => Sel(1), A2 => Sel(2), A3 => n319, ZN => n313);
   U49 : INV_X1 port map( A => Sel(0), ZN => n319);
   U50 : BUF_X1 port map( A => n315, Z => n176);
   U51 : NOR2_X1 port map( A1 => n165, A2 => n186, ZN => n315);
   U52 : AOI21_X1 port map( B1 => n319, B2 => n320, A => Sel(2), ZN => n186);
   U53 : NAND2_X1 port map( A1 => n200, A2 => n199, ZN => Y(15));
   U54 : AOI22_X1 port map( A1 => A_neg(15), A2 => n151, B1 => A_signal(15), B2
                           => n142, ZN => n200);
   U55 : AOI222_X1 port map( A1 => A_shifted(14), A2 => n177, B1 => 
                           zeroSignal(14), B2 => n168, C1 => A_neg_shifted(14),
                           C2 => n164, ZN => n197);
   U56 : NAND2_X1 port map( A1 => n202, A2 => n201, ZN => Y(16));
   U57 : AOI22_X1 port map( A1 => A_neg(16), A2 => n151, B1 => A_signal(16), B2
                           => n142, ZN => n202);
   U58 : AOI222_X1 port map( A1 => A_shifted(16), A2 => n177, B1 => 
                           zeroSignal(16), B2 => n168, C1 => A_neg_shifted(16),
                           C2 => n164, ZN => n201);
   U59 : NAND2_X1 port map( A1 => n204, A2 => n203, ZN => Y(17));
   U60 : AOI22_X1 port map( A1 => A_neg(17), A2 => n151, B1 => A_signal(17), B2
                           => n142, ZN => n204);
   U61 : AOI222_X1 port map( A1 => A_shifted(17), A2 => n177, B1 => 
                           zeroSignal(17), B2 => n168, C1 => A_neg_shifted(17),
                           C2 => n164, ZN => n203);
   U62 : NAND2_X1 port map( A1 => n206, A2 => n205, ZN => Y(18));
   U63 : AOI22_X1 port map( A1 => A_neg(18), A2 => n151, B1 => A_signal(18), B2
                           => n142, ZN => n206);
   U64 : AOI222_X1 port map( A1 => A_shifted(18), A2 => n177, B1 => 
                           zeroSignal(18), B2 => n168, C1 => A_neg_shifted(18),
                           C2 => n164, ZN => n205);
   U65 : NAND2_X1 port map( A1 => n222, A2 => n221, ZN => Y(25));
   U66 : AOI22_X1 port map( A1 => A_neg(25), A2 => n152, B1 => A_signal(25), B2
                           => n143, ZN => n222);
   U67 : AOI222_X1 port map( A1 => A_shifted(25), A2 => n178, B1 => 
                           zeroSignal(25), B2 => n169, C1 => A_neg_shifted(25),
                           C2 => n163, ZN => n221);
   U68 : NAND2_X1 port map( A1 => n224, A2 => n223, ZN => Y(26));
   U69 : AOI22_X1 port map( A1 => A_neg(26), A2 => n152, B1 => A_signal(26), B2
                           => n143, ZN => n224);
   U70 : AOI222_X1 port map( A1 => A_shifted(26), A2 => n178, B1 => 
                           zeroSignal(26), B2 => n169, C1 => A_neg_shifted(26),
                           C2 => n163, ZN => n223);
   U71 : NAND2_X1 port map( A1 => n208, A2 => n207, ZN => Y(19));
   U72 : AOI22_X1 port map( A1 => A_neg(19), A2 => n151, B1 => A_signal(19), B2
                           => n142, ZN => n208);
   U73 : AOI222_X1 port map( A1 => A_shifted(19), A2 => n177, B1 => 
                           zeroSignal(19), B2 => n168, C1 => A_neg_shifted(19),
                           C2 => n164, ZN => n207);
   U74 : NAND2_X1 port map( A1 => n226, A2 => n225, ZN => Y(27));
   U75 : AOI22_X1 port map( A1 => A_neg(27), A2 => n152, B1 => A_signal(27), B2
                           => n143, ZN => n226);
   U76 : AOI222_X1 port map( A1 => A_shifted(27), A2 => n178, B1 => 
                           zeroSignal(27), B2 => n169, C1 => A_neg_shifted(27),
                           C2 => n163, ZN => n225);
   U77 : NAND2_X1 port map( A1 => n228, A2 => n227, ZN => Y(28));
   U78 : AOI22_X1 port map( A1 => A_neg(28), A2 => n152, B1 => A_signal(28), B2
                           => n143, ZN => n228);
   U79 : AOI222_X1 port map( A1 => A_shifted(28), A2 => n178, B1 => 
                           zeroSignal(28), B2 => n169, C1 => A_neg_shifted(28),
                           C2 => n163, ZN => n227);
   U80 : NAND2_X1 port map( A1 => n234, A2 => n233, ZN => Y(30));
   U81 : AOI22_X1 port map( A1 => A_neg(30), A2 => n152, B1 => A_signal(30), B2
                           => n143, ZN => n234);
   U82 : AOI222_X1 port map( A1 => A_shifted(30), A2 => n178, B1 => 
                           zeroSignal(30), B2 => n169, C1 => A_neg_shifted(30),
                           C2 => n163, ZN => n233);
   U83 : NAND2_X1 port map( A1 => n236, A2 => n235, ZN => Y(31));
   U84 : AOI22_X1 port map( A1 => A_neg(31), A2 => n153, B1 => A_signal(31), B2
                           => n144, ZN => n236);
   U85 : AOI222_X1 port map( A1 => A_shifted(31), A2 => n179, B1 => 
                           zeroSignal(31), B2 => n170, C1 => A_neg_shifted(31),
                           C2 => n163, ZN => n235);
   U86 : NAND2_X1 port map( A1 => n238, A2 => n237, ZN => Y(32));
   U87 : AOI22_X1 port map( A1 => A_neg(32), A2 => n153, B1 => A_signal(32), B2
                           => n144, ZN => n238);
   U88 : AOI222_X1 port map( A1 => A_shifted(32), A2 => n179, B1 => 
                           zeroSignal(32), B2 => n170, C1 => A_neg_shifted(32),
                           C2 => n163, ZN => n237);
   U89 : NAND2_X1 port map( A1 => n244, A2 => n243, ZN => Y(35));
   U90 : AOI22_X1 port map( A1 => A_neg(35), A2 => n153, B1 => A_signal(35), B2
                           => n144, ZN => n244);
   U91 : AOI222_X1 port map( A1 => A_shifted(35), A2 => n179, B1 => 
                           zeroSignal(35), B2 => n170, C1 => A_neg_shifted(35),
                           C2 => n162, ZN => n243);
   U92 : NAND2_X1 port map( A1 => n242, A2 => n241, ZN => Y(34));
   U93 : AOI22_X1 port map( A1 => A_neg(34), A2 => n153, B1 => A_signal(34), B2
                           => n144, ZN => n242);
   U94 : AOI222_X1 port map( A1 => A_shifted(34), A2 => n179, B1 => 
                           zeroSignal(34), B2 => n170, C1 => A_neg_shifted(34),
                           C2 => n163, ZN => n241);
   U95 : NAND2_X1 port map( A1 => n246, A2 => n245, ZN => Y(36));
   U96 : AOI22_X1 port map( A1 => A_neg(36), A2 => n153, B1 => A_signal(36), B2
                           => n144, ZN => n246);
   U97 : AOI222_X1 port map( A1 => A_shifted(36), A2 => n179, B1 => 
                           zeroSignal(36), B2 => n170, C1 => A_neg_shifted(36),
                           C2 => n162, ZN => n245);
   U98 : NAND2_X1 port map( A1 => n270, A2 => n269, ZN => Y(47));
   U99 : AOI222_X1 port map( A1 => A_shifted(47), A2 => n180, B1 => 
                           zeroSignal(47), B2 => n171, C1 => A_neg_shifted(47),
                           C2 => n161, ZN => n269);
   U100 : AOI22_X1 port map( A1 => A_neg(47), A2 => n154, B1 => A_signal(47), 
                           B2 => n145, ZN => n270);
   U101 : NAND2_X1 port map( A1 => n212, A2 => n211, ZN => Y(20));
   U102 : AOI22_X1 port map( A1 => A_neg(20), A2 => n152, B1 => A_signal(20), 
                           B2 => n143, ZN => n212);
   U103 : AOI222_X1 port map( A1 => A_shifted(20), A2 => n178, B1 => 
                           zeroSignal(20), B2 => n169, C1 => A_neg_shifted(20),
                           C2 => n164, ZN => n211);
   U104 : NAND2_X1 port map( A1 => n248, A2 => n247, ZN => Y(37));
   U105 : AOI22_X1 port map( A1 => A_neg(37), A2 => n153, B1 => A_signal(37), 
                           B2 => n144, ZN => n248);
   U106 : AOI222_X1 port map( A1 => A_shifted(37), A2 => n179, B1 => 
                           zeroSignal(37), B2 => n170, C1 => A_neg_shifted(37),
                           C2 => n162, ZN => n247);
   U107 : NAND2_X1 port map( A1 => n250, A2 => n249, ZN => Y(38));
   U108 : AOI22_X1 port map( A1 => A_neg(38), A2 => n153, B1 => A_signal(38), 
                           B2 => n144, ZN => n250);
   U109 : AOI222_X1 port map( A1 => A_shifted(38), A2 => n179, B1 => 
                           zeroSignal(38), B2 => n170, C1 => A_neg_shifted(38),
                           C2 => n162, ZN => n249);
   U110 : NAND2_X1 port map( A1 => n214, A2 => n213, ZN => Y(21));
   U111 : AOI22_X1 port map( A1 => A_neg(21), A2 => n152, B1 => A_signal(21), 
                           B2 => n143, ZN => n214);
   U112 : AOI222_X1 port map( A1 => A_shifted(21), A2 => n178, B1 => 
                           zeroSignal(21), B2 => n169, C1 => A_neg_shifted(21),
                           C2 => n164, ZN => n213);
   U113 : NAND2_X1 port map( A1 => n256, A2 => n255, ZN => Y(40));
   U114 : AOI22_X1 port map( A1 => A_neg(40), A2 => n153, B1 => A_signal(40), 
                           B2 => n144, ZN => n256);
   U115 : AOI222_X1 port map( A1 => A_shifted(40), A2 => n179, B1 => 
                           zeroSignal(40), B2 => n170, C1 => A_neg_shifted(40),
                           C2 => n162, ZN => n255);
   U116 : NAND2_X1 port map( A1 => n216, A2 => n215, ZN => Y(22));
   U117 : AOI22_X1 port map( A1 => A_neg(22), A2 => n152, B1 => A_signal(22), 
                           B2 => n143, ZN => n216);
   U118 : AOI222_X1 port map( A1 => A_shifted(22), A2 => n178, B1 => 
                           zeroSignal(22), B2 => n169, C1 => A_neg_shifted(22),
                           C2 => n164, ZN => n215);
   U119 : NAND2_X1 port map( A1 => n258, A2 => n257, ZN => Y(41));
   U120 : AOI22_X1 port map( A1 => A_neg(41), A2 => n153, B1 => A_signal(41), 
                           B2 => n144, ZN => n258);
   U121 : AOI222_X1 port map( A1 => A_shifted(41), A2 => n179, B1 => 
                           zeroSignal(41), B2 => n170, C1 => A_neg_shifted(41),
                           C2 => n162, ZN => n257);
   U122 : NAND2_X1 port map( A1 => n260, A2 => n259, ZN => Y(42));
   U123 : AOI22_X1 port map( A1 => A_neg(42), A2 => n154, B1 => A_signal(42), 
                           B2 => n145, ZN => n260);
   U124 : AOI222_X1 port map( A1 => A_shifted(42), A2 => n180, B1 => 
                           zeroSignal(42), B2 => n171, C1 => A_neg_shifted(42),
                           C2 => n162, ZN => n259);
   U125 : NAND2_X1 port map( A1 => n218, A2 => n217, ZN => Y(23));
   U126 : AOI22_X1 port map( A1 => A_neg(23), A2 => n152, B1 => A_signal(23), 
                           B2 => n143, ZN => n218);
   U127 : AOI222_X1 port map( A1 => A_shifted(23), A2 => n178, B1 => 
                           zeroSignal(23), B2 => n169, C1 => A_neg_shifted(23),
                           C2 => n164, ZN => n217);
   U128 : NAND2_X1 port map( A1 => n220, A2 => n219, ZN => Y(24));
   U129 : AOI22_X1 port map( A1 => A_neg(24), A2 => n152, B1 => A_signal(24), 
                           B2 => n143, ZN => n220);
   U130 : AOI222_X1 port map( A1 => A_shifted(24), A2 => n178, B1 => 
                           zeroSignal(24), B2 => n169, C1 => A_neg_shifted(24),
                           C2 => n163, ZN => n219);
   U131 : NAND2_X1 port map( A1 => n262, A2 => n261, ZN => Y(43));
   U132 : AOI22_X1 port map( A1 => A_neg(43), A2 => n154, B1 => A_signal(43), 
                           B2 => n145, ZN => n262);
   U133 : AOI222_X1 port map( A1 => A_shifted(43), A2 => n180, B1 => 
                           zeroSignal(43), B2 => n171, C1 => A_neg_shifted(43),
                           C2 => n162, ZN => n261);
   U134 : NAND2_X1 port map( A1 => n264, A2 => n263, ZN => Y(44));
   U135 : AOI22_X1 port map( A1 => A_neg(44), A2 => n154, B1 => A_signal(44), 
                           B2 => n145, ZN => n264);
   U136 : AOI222_X1 port map( A1 => A_shifted(44), A2 => n180, B1 => 
                           zeroSignal(44), B2 => n171, C1 => A_neg_shifted(44),
                           C2 => n162, ZN => n263);
   U137 : NAND2_X1 port map( A1 => n266, A2 => n265, ZN => Y(45));
   U138 : AOI22_X1 port map( A1 => A_neg(45), A2 => n154, B1 => A_signal(45), 
                           B2 => n145, ZN => n266);
   U139 : AOI222_X1 port map( A1 => A_shifted(45), A2 => n180, B1 => 
                           zeroSignal(45), B2 => n171, C1 => A_neg_shifted(45),
                           C2 => n162, ZN => n265);
   U140 : NAND2_X1 port map( A1 => n268, A2 => n267, ZN => Y(46));
   U141 : AOI22_X1 port map( A1 => A_neg(46), A2 => n154, B1 => A_signal(46), 
                           B2 => n145, ZN => n268);
   U142 : AOI222_X1 port map( A1 => A_shifted(46), A2 => n180, B1 => 
                           zeroSignal(46), B2 => n171, C1 => A_neg_shifted(46),
                           C2 => n161, ZN => n267);
   U143 : NAND2_X1 port map( A1 => n272, A2 => n271, ZN => Y(48));
   U144 : AOI22_X1 port map( A1 => A_neg(48), A2 => n154, B1 => A_signal(48), 
                           B2 => n145, ZN => n272);
   U145 : AOI222_X1 port map( A1 => A_shifted(48), A2 => n180, B1 => 
                           zeroSignal(48), B2 => n171, C1 => A_neg_shifted(48),
                           C2 => n161, ZN => n271);
   U146 : NAND2_X1 port map( A1 => n274, A2 => n273, ZN => Y(49));
   U147 : AOI222_X1 port map( A1 => A_shifted(49), A2 => n180, B1 => 
                           zeroSignal(49), B2 => n171, C1 => A_neg_shifted(49),
                           C2 => n161, ZN => n273);
   U148 : AOI22_X1 port map( A1 => A_neg(49), A2 => n154, B1 => A_signal(49), 
                           B2 => n145, ZN => n274);
   U149 : NAND2_X1 port map( A1 => n230, A2 => n229, ZN => Y(29));
   U150 : AOI22_X1 port map( A1 => A_neg(29), A2 => n152, B1 => A_signal(29), 
                           B2 => n143, ZN => n230);
   U151 : AOI222_X1 port map( A1 => A_shifted(29), A2 => n178, B1 => 
                           zeroSignal(29), B2 => n169, C1 => A_neg_shifted(29),
                           C2 => n163, ZN => n229);
   U152 : NAND2_X1 port map( A1 => n278, A2 => n277, ZN => Y(50));
   U153 : AOI222_X1 port map( A1 => A_shifted(50), A2 => n180, B1 => 
                           zeroSignal(50), B2 => n171, C1 => A_neg_shifted(50),
                           C2 => n161, ZN => n277);
   U154 : AOI22_X1 port map( A1 => A_neg(50), A2 => n154, B1 => A_signal(50), 
                           B2 => n145, ZN => n278);
   U155 : NAND2_X1 port map( A1 => n240, A2 => n239, ZN => Y(33));
   U156 : AOI22_X1 port map( A1 => A_neg(33), A2 => n153, B1 => A_signal(33), 
                           B2 => n144, ZN => n240);
   U157 : AOI222_X1 port map( A1 => A_shifted(33), A2 => n179, B1 => 
                           zeroSignal(33), B2 => n170, C1 => A_neg_shifted(33),
                           C2 => n163, ZN => n239);
   U158 : NAND2_X1 port map( A1 => n280, A2 => n279, ZN => Y(51));
   U159 : AOI22_X1 port map( A1 => A_neg(51), A2 => n154, B1 => A_signal(51), 
                           B2 => n145, ZN => n280);
   U160 : AOI222_X1 port map( A1 => A_shifted(51), A2 => n180, B1 => 
                           zeroSignal(51), B2 => n171, C1 => A_neg_shifted(51),
                           C2 => n161, ZN => n279);
   U161 : NAND2_X1 port map( A1 => n252, A2 => n251, ZN => Y(39));
   U162 : AOI22_X1 port map( A1 => A_neg(39), A2 => n153, B1 => A_signal(39), 
                           B2 => n144, ZN => n252);
   U163 : AOI222_X1 port map( A1 => A_shifted(39), A2 => n179, B1 => 
                           zeroSignal(39), B2 => n170, C1 => A_neg_shifted(39),
                           C2 => n162, ZN => n251);
   U164 : NAND2_X1 port map( A1 => n284, A2 => n283, ZN => Y(53));
   U165 : AOI222_X1 port map( A1 => A_shifted(53), A2 => n181, B1 => 
                           zeroSignal(53), B2 => n172, C1 => A_neg_shifted(53),
                           C2 => n161, ZN => n283);
   U166 : AOI22_X1 port map( A1 => A_neg(53), A2 => n155, B1 => A_signal(53), 
                           B2 => n146, ZN => n284);
   U167 : NAND2_X1 port map( A1 => n282, A2 => n281, ZN => Y(52));
   U168 : AOI222_X1 port map( A1 => A_shifted(52), A2 => n180, B1 => 
                           zeroSignal(52), B2 => n171, C1 => A_neg_shifted(52),
                           C2 => n161, ZN => n281);
   U169 : AOI22_X1 port map( A1 => A_neg(52), A2 => n154, B1 => A_signal(52), 
                           B2 => n145, ZN => n282);
   U170 : NAND2_X1 port map( A1 => n286, A2 => n285, ZN => Y(54));
   U171 : AOI222_X1 port map( A1 => A_shifted(54), A2 => n181, B1 => 
                           zeroSignal(54), B2 => n172, C1 => A_neg_shifted(54),
                           C2 => n161, ZN => n285);
   U172 : AOI22_X1 port map( A1 => A_neg(54), A2 => n155, B1 => A_signal(54), 
                           B2 => n146, ZN => n286);
   U173 : NAND2_X1 port map( A1 => n288, A2 => n287, ZN => Y(55));
   U174 : AOI22_X1 port map( A1 => A_neg(55), A2 => n155, B1 => A_signal(55), 
                           B2 => n146, ZN => n288);
   U175 : AOI222_X1 port map( A1 => A_shifted(55), A2 => n181, B1 => 
                           zeroSignal(55), B2 => n172, C1 => A_neg_shifted(55),
                           C2 => n161, ZN => n287);
   U176 : NAND2_X1 port map( A1 => n304, A2 => n303, ZN => Y(62));
   U177 : NAND2_X1 port map( A1 => n294, A2 => n293, ZN => Y(58));
   U178 : AOI222_X1 port map( A1 => A_shifted(58), A2 => n181, B1 => 
                           zeroSignal(58), B2 => n172, C1 => A_neg_shifted(58),
                           C2 => n160, ZN => n293);
   U179 : NAND2_X1 port map( A1 => n302, A2 => n301, ZN => Y(61));
   U180 : NAND2_X1 port map( A1 => n292, A2 => n291, ZN => Y(57));
   U181 : AOI222_X1 port map( A1 => A_shifted(57), A2 => n181, B1 => 
                           zeroSignal(57), B2 => n172, C1 => A_neg_shifted(57),
                           C2 => n160, ZN => n291);
   U182 : AOI22_X1 port map( A1 => A_neg(57), A2 => n155, B1 => A_signal(57), 
                           B2 => n146, ZN => n292);
   U183 : NAND2_X1 port map( A1 => n300, A2 => n299, ZN => Y(60));
   U184 : AOI222_X1 port map( A1 => A_shifted(60), A2 => n181, B1 => 
                           zeroSignal(60), B2 => n172, C1 => A_neg_shifted(60),
                           C2 => n160, ZN => n299);
   U185 : NAND2_X1 port map( A1 => n296, A2 => n295, ZN => Y(59));
   U186 : AOI22_X1 port map( A1 => A_neg(59), A2 => n155, B1 => A_signal(59), 
                           B2 => n146, ZN => n296);
   U187 : NAND2_X1 port map( A1 => n306, A2 => n305, ZN => Y(63));
   U188 : AOI22_X1 port map( A1 => A_neg(63), A2 => n155, B1 => A_signal(63), 
                           B2 => n146, ZN => n306);
   U189 : NAND2_X1 port map( A1 => n290, A2 => n289, ZN => Y(56));
   U190 : AOI22_X1 port map( A1 => A_neg(56), A2 => n155, B1 => A_signal(56), 
                           B2 => n146, ZN => n290);
   U191 : AOI222_X1 port map( A1 => A_shifted(56), A2 => n181, B1 => 
                           zeroSignal(56), B2 => n172, C1 => A_neg_shifted(56),
                           C2 => n161, ZN => n289);
   U192 : NAND2_X1 port map( A1 => n188, A2 => n187, ZN => Y(0));
   U193 : AOI22_X1 port map( A1 => A_neg(0), A2 => n151, B1 => A_signal(0), B2 
                           => n142, ZN => n188);
   U194 : AOI222_X1 port map( A1 => A_shifted(0), A2 => n177, B1 => 
                           zeroSignal(0), B2 => n168, C1 => A_neg_shifted(0), 
                           C2 => n165, ZN => n187);
   U195 : NAND2_X1 port map( A1 => n210, A2 => n209, ZN => Y(1));
   U196 : AOI22_X1 port map( A1 => A_neg(1), A2 => n151, B1 => A_signal(1), B2 
                           => n142, ZN => n210);
   U197 : AOI222_X1 port map( A1 => A_shifted(1), A2 => n177, B1 => 
                           zeroSignal(1), B2 => n168, C1 => A_neg_shifted(1), 
                           C2 => n164, ZN => n209);
   U198 : NAND2_X1 port map( A1 => n232, A2 => n231, ZN => Y(2));
   U199 : AOI22_X1 port map( A1 => A_neg(2), A2 => n152, B1 => A_signal(2), B2 
                           => n143, ZN => n232);
   U200 : AOI222_X1 port map( A1 => A_shifted(2), A2 => n178, B1 => 
                           zeroSignal(2), B2 => n169, C1 => A_neg_shifted(2), 
                           C2 => n163, ZN => n231);
   U201 : NAND2_X1 port map( A1 => n254, A2 => n253, ZN => Y(3));
   U202 : AOI22_X1 port map( A1 => A_neg(3), A2 => n153, B1 => A_signal(3), B2 
                           => n144, ZN => n254);
   U203 : AOI222_X1 port map( A1 => A_shifted(3), A2 => n179, B1 => 
                           zeroSignal(3), B2 => n170, C1 => A_neg_shifted(3), 
                           C2 => n162, ZN => n253);
   U204 : NAND2_X1 port map( A1 => n276, A2 => n275, ZN => Y(4));
   U205 : AOI22_X1 port map( A1 => A_neg(4), A2 => n154, B1 => A_signal(4), B2 
                           => n145, ZN => n276);
   U206 : AOI222_X1 port map( A1 => A_shifted(4), A2 => n180, B1 => 
                           zeroSignal(4), B2 => n171, C1 => A_neg_shifted(4), 
                           C2 => n161, ZN => n275);
   U207 : NAND2_X1 port map( A1 => n298, A2 => n297, ZN => Y(5));
   U208 : AOI22_X1 port map( A1 => A_neg(5), A2 => n155, B1 => A_signal(5), B2 
                           => n146, ZN => n298);
   U209 : AOI222_X1 port map( A1 => A_shifted(5), A2 => n181, B1 => 
                           zeroSignal(5), B2 => n172, C1 => A_neg_shifted(5), 
                           C2 => n160, ZN => n297);
   U210 : NAND2_X1 port map( A1 => n308, A2 => n307, ZN => Y(6));
   U211 : AOI22_X1 port map( A1 => A_neg(6), A2 => n156, B1 => A_signal(6), B2 
                           => n147, ZN => n308);
   U212 : AOI222_X1 port map( A1 => A_shifted(6), A2 => n182, B1 => 
                           zeroSignal(6), B2 => n173, C1 => A_neg_shifted(6), 
                           C2 => n160, ZN => n307);
   U213 : NAND2_X1 port map( A1 => n310, A2 => n309, ZN => Y(7));
   U214 : AOI22_X1 port map( A1 => A_neg(7), A2 => n156, B1 => A_signal(7), B2 
                           => n147, ZN => n310);
   U215 : AOI222_X1 port map( A1 => A_shifted(7), A2 => n182, B1 => 
                           zeroSignal(7), B2 => n173, C1 => A_neg_shifted(7), 
                           C2 => n160, ZN => n309);
   U216 : NAND2_X1 port map( A1 => n312, A2 => n311, ZN => Y(8));
   U217 : AOI22_X1 port map( A1 => A_neg(8), A2 => n156, B1 => A_signal(8), B2 
                           => n147, ZN => n312);
   U218 : AOI222_X1 port map( A1 => A_shifted(8), A2 => n182, B1 => 
                           zeroSignal(8), B2 => n173, C1 => A_neg_shifted(8), 
                           C2 => n160, ZN => n311);
   U219 : NAND2_X1 port map( A1 => n318, A2 => n317, ZN => Y(9));
   U220 : AOI22_X1 port map( A1 => A_neg(9), A2 => n156, B1 => A_signal(9), B2 
                           => n147, ZN => n318);
   U221 : AOI222_X1 port map( A1 => A_shifted(9), A2 => n182, B1 => 
                           zeroSignal(9), B2 => n173, C1 => A_neg_shifted(9), 
                           C2 => n160, ZN => n317);
   U222 : NAND2_X1 port map( A1 => n190, A2 => n189, ZN => Y(10));
   U223 : AOI22_X1 port map( A1 => A_neg(10), A2 => n151, B1 => A_signal(10), 
                           B2 => n142, ZN => n190);
   U224 : AOI222_X1 port map( A1 => A_shifted(10), A2 => n177, B1 => 
                           zeroSignal(10), B2 => n168, C1 => A_neg_shifted(10),
                           C2 => n165, ZN => n189);
   U225 : NAND2_X1 port map( A1 => n192, A2 => n191, ZN => Y(11));
   U226 : AOI22_X1 port map( A1 => A_neg(11), A2 => n151, B1 => A_signal(11), 
                           B2 => n142, ZN => n192);
   U227 : AOI222_X1 port map( A1 => A_shifted(11), A2 => n177, B1 => 
                           zeroSignal(11), B2 => n168, C1 => A_neg_shifted(11),
                           C2 => n165, ZN => n191);
   U228 : NAND2_X1 port map( A1 => n194, A2 => n193, ZN => Y(12));
   U229 : AOI22_X1 port map( A1 => A_neg(12), A2 => n151, B1 => A_signal(12), 
                           B2 => n142, ZN => n194);
   U230 : AOI222_X1 port map( A1 => A_shifted(12), A2 => n177, B1 => 
                           zeroSignal(12), B2 => n168, C1 => A_neg_shifted(12),
                           C2 => n165, ZN => n193);
   U231 : NAND2_X1 port map( A1 => n196, A2 => n195, ZN => Y(13));
   U232 : AOI22_X1 port map( A1 => A_neg(13), A2 => n151, B1 => A_signal(13), 
                           B2 => n142, ZN => n196);
   U233 : AOI222_X1 port map( A1 => A_shifted(13), A2 => n177, B1 => 
                           zeroSignal(13), B2 => n168, C1 => A_neg_shifted(13),
                           C2 => n164, ZN => n195);
   U234 : AOI222_X1 port map( A1 => A_shifted(63), A2 => n181, B1 => 
                           zeroSignal(63), B2 => n172, C1 => A_neg_shifted(63),
                           C2 => n160, ZN => n305);
   U235 : AOI22_X1 port map( A1 => A_neg(62), A2 => n155, B1 => A_signal(62), 
                           B2 => n146, ZN => n304);
   U236 : AOI222_X1 port map( A1 => A_shifted(61), A2 => n181, B1 => 
                           zeroSignal(61), B2 => n172, C1 => A_neg_shifted(61),
                           C2 => n160, ZN => n301);
   U237 : AOI22_X1 port map( A1 => A_neg(60), A2 => n155, B1 => A_signal(60), 
                           B2 => n146, ZN => n300);
   U238 : AOI222_X1 port map( A1 => A_shifted(62), A2 => n181, B1 => 
                           zeroSignal(62), B2 => n172, C1 => A_neg_shifted(62),
                           C2 => n160, ZN => n303);
   U239 : AOI22_X1 port map( A1 => A_neg(61), A2 => n155, B1 => A_signal(61), 
                           B2 => n146, ZN => n302);
   U240 : AOI222_X1 port map( A1 => A_shifted(59), A2 => n181, B1 => 
                           zeroSignal(59), B2 => n172, C1 => A_neg_shifted(59),
                           C2 => n160, ZN => n295);
   U241 : AOI22_X1 port map( A1 => A_neg(58), A2 => n155, B1 => A_signal(58), 
                           B2 => n146, ZN => n294);
   U242 : AOI22_X1 port map( A1 => A_neg(14), A2 => n151, B1 => A_signal(14), 
                           B2 => n142, ZN => n198);
   U243 : AOI222_X1 port map( A1 => A_shifted(15), A2 => n177, B1 => 
                           zeroSignal(15), B2 => n168, C1 => A_neg_shifted(15),
                           C2 => n164, ZN => n199);
   U244 : NAND2_X1 port map( A1 => n198, A2 => n197, ZN => Y(14));

end SYN_BEHAVIORAL_2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity MUX51_MuxNbit64_24 is

   port( zeroSignal, A_signal, A_neg, A_shifted, A_neg_shifted : in 
         std_logic_vector (63 downto 0);  Sel : in std_logic_vector (2 downto 
         0);  Y : out std_logic_vector (63 downto 0));

end MUX51_MuxNbit64_24;

architecture SYN_BEHAVIORAL_2 of MUX51_MuxNbit64_24 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, 
      n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, 
      n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, 
      n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, 
      n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, 
      n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, 
      n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, 
      n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, 
      n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, 
      n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, 
      n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, 
      n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, 
      n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, 
      n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, 
      n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, 
      n320 : std_logic;

begin
   
   U1 : AND3_X1 port map( A1 => n319, A2 => n320, A3 => Sel(2), ZN => n141);
   U2 : BUF_X1 port map( A => n141, Z => n166);
   U3 : BUF_X1 port map( A => n185, Z => n184);
   U4 : BUF_X1 port map( A => n159, Z => n158);
   U5 : BUF_X1 port map( A => n150, Z => n149);
   U6 : BUF_X1 port map( A => n141, Z => n167);
   U7 : BUF_X1 port map( A => n185, Z => n183);
   U8 : BUF_X1 port map( A => n159, Z => n157);
   U9 : BUF_X1 port map( A => n150, Z => n148);
   U10 : BUF_X1 port map( A => n176, Z => n175);
   U11 : BUF_X1 port map( A => n176, Z => n174);
   U12 : BUF_X1 port map( A => n158, Z => n151);
   U13 : BUF_X1 port map( A => n184, Z => n177);
   U14 : BUF_X1 port map( A => n149, Z => n142);
   U15 : BUF_X1 port map( A => n166, Z => n164);
   U16 : BUF_X1 port map( A => n184, Z => n178);
   U17 : BUF_X1 port map( A => n158, Z => n152);
   U18 : BUF_X1 port map( A => n149, Z => n143);
   U19 : BUF_X1 port map( A => n166, Z => n163);
   U20 : BUF_X1 port map( A => n184, Z => n179);
   U21 : BUF_X1 port map( A => n158, Z => n153);
   U22 : BUF_X1 port map( A => n149, Z => n144);
   U23 : BUF_X1 port map( A => n167, Z => n162);
   U24 : BUF_X1 port map( A => n183, Z => n180);
   U25 : BUF_X1 port map( A => n157, Z => n154);
   U26 : BUF_X1 port map( A => n148, Z => n145);
   U27 : BUF_X1 port map( A => n167, Z => n161);
   U28 : BUF_X1 port map( A => n183, Z => n181);
   U29 : BUF_X1 port map( A => n157, Z => n155);
   U30 : BUF_X1 port map( A => n148, Z => n146);
   U31 : BUF_X1 port map( A => n167, Z => n160);
   U32 : BUF_X1 port map( A => n175, Z => n169);
   U33 : BUF_X1 port map( A => n175, Z => n170);
   U34 : BUF_X1 port map( A => n174, Z => n171);
   U35 : BUF_X1 port map( A => n175, Z => n168);
   U36 : BUF_X1 port map( A => n174, Z => n172);
   U37 : BUF_X1 port map( A => n166, Z => n165);
   U38 : BUF_X1 port map( A => n157, Z => n156);
   U39 : BUF_X1 port map( A => n148, Z => n147);
   U40 : BUF_X1 port map( A => n174, Z => n173);
   U41 : BUF_X1 port map( A => n183, Z => n182);
   U42 : BUF_X1 port map( A => n314, Z => n159);
   U43 : NOR3_X1 port map( A1 => Sel(0), A2 => Sel(2), A3 => n320, ZN => n314);
   U44 : INV_X1 port map( A => Sel(1), ZN => n320);
   U45 : BUF_X1 port map( A => n316, Z => n185);
   U46 : NOR3_X1 port map( A1 => n319, A2 => Sel(2), A3 => n320, ZN => n316);
   U47 : BUF_X1 port map( A => n313, Z => n150);
   U48 : NOR3_X1 port map( A1 => Sel(1), A2 => Sel(2), A3 => n319, ZN => n313);
   U49 : INV_X1 port map( A => Sel(0), ZN => n319);
   U50 : BUF_X1 port map( A => n315, Z => n176);
   U51 : NOR2_X1 port map( A1 => n165, A2 => n186, ZN => n315);
   U52 : AOI21_X1 port map( B1 => n319, B2 => n320, A => Sel(2), ZN => n186);
   U53 : NAND2_X1 port map( A1 => n204, A2 => n203, ZN => Y(17));
   U54 : AOI22_X1 port map( A1 => A_neg(17), A2 => n151, B1 => A_signal(17), B2
                           => n142, ZN => n204);
   U55 : NAND2_X1 port map( A1 => n202, A2 => n201, ZN => Y(16));
   U56 : AOI222_X1 port map( A1 => A_shifted(16), A2 => n177, B1 => 
                           zeroSignal(16), B2 => n168, C1 => A_neg_shifted(16),
                           C2 => n164, ZN => n201);
   U57 : NAND2_X1 port map( A1 => n206, A2 => n205, ZN => Y(18));
   U58 : AOI22_X1 port map( A1 => A_neg(18), A2 => n151, B1 => A_signal(18), B2
                           => n142, ZN => n206);
   U59 : AOI222_X1 port map( A1 => A_shifted(18), A2 => n177, B1 => 
                           zeroSignal(18), B2 => n168, C1 => A_neg_shifted(18),
                           C2 => n164, ZN => n205);
   U60 : NAND2_X1 port map( A1 => n208, A2 => n207, ZN => Y(19));
   U61 : AOI22_X1 port map( A1 => A_neg(19), A2 => n151, B1 => A_signal(19), B2
                           => n142, ZN => n208);
   U62 : AOI222_X1 port map( A1 => A_shifted(19), A2 => n177, B1 => 
                           zeroSignal(19), B2 => n168, C1 => A_neg_shifted(19),
                           C2 => n164, ZN => n207);
   U63 : NAND2_X1 port map( A1 => n212, A2 => n211, ZN => Y(20));
   U64 : AOI22_X1 port map( A1 => A_neg(20), A2 => n152, B1 => A_signal(20), B2
                           => n143, ZN => n212);
   U65 : AOI222_X1 port map( A1 => A_shifted(20), A2 => n178, B1 => 
                           zeroSignal(20), B2 => n169, C1 => A_neg_shifted(20),
                           C2 => n164, ZN => n211);
   U66 : NAND2_X1 port map( A1 => n228, A2 => n227, ZN => Y(28));
   U67 : AOI222_X1 port map( A1 => A_shifted(28), A2 => n178, B1 => 
                           zeroSignal(28), B2 => n169, C1 => A_neg_shifted(28),
                           C2 => n163, ZN => n227);
   U68 : AOI22_X1 port map( A1 => A_neg(28), A2 => n152, B1 => A_signal(28), B2
                           => n143, ZN => n228);
   U69 : NAND2_X1 port map( A1 => n224, A2 => n223, ZN => Y(26));
   U70 : AOI222_X1 port map( A1 => A_shifted(26), A2 => n178, B1 => 
                           zeroSignal(26), B2 => n169, C1 => A_neg_shifted(26),
                           C2 => n163, ZN => n223);
   U71 : AOI22_X1 port map( A1 => A_neg(26), A2 => n152, B1 => A_signal(26), B2
                           => n143, ZN => n224);
   U72 : NAND2_X1 port map( A1 => n226, A2 => n225, ZN => Y(27));
   U73 : AOI222_X1 port map( A1 => A_shifted(27), A2 => n178, B1 => 
                           zeroSignal(27), B2 => n169, C1 => A_neg_shifted(27),
                           C2 => n163, ZN => n225);
   U74 : AOI22_X1 port map( A1 => A_neg(27), A2 => n152, B1 => A_signal(27), B2
                           => n143, ZN => n226);
   U75 : NAND2_X1 port map( A1 => n236, A2 => n235, ZN => Y(31));
   U76 : AOI222_X1 port map( A1 => A_shifted(31), A2 => n179, B1 => 
                           zeroSignal(31), B2 => n170, C1 => A_neg_shifted(31),
                           C2 => n163, ZN => n235);
   U77 : AOI22_X1 port map( A1 => A_neg(31), A2 => n153, B1 => A_signal(31), B2
                           => n144, ZN => n236);
   U78 : NAND2_X1 port map( A1 => n230, A2 => n229, ZN => Y(29));
   U79 : AOI222_X1 port map( A1 => A_shifted(29), A2 => n178, B1 => 
                           zeroSignal(29), B2 => n169, C1 => A_neg_shifted(29),
                           C2 => n163, ZN => n229);
   U80 : AOI22_X1 port map( A1 => A_neg(29), A2 => n152, B1 => A_signal(29), B2
                           => n143, ZN => n230);
   U81 : NAND2_X1 port map( A1 => n238, A2 => n237, ZN => Y(32));
   U82 : AOI222_X1 port map( A1 => A_shifted(32), A2 => n179, B1 => 
                           zeroSignal(32), B2 => n170, C1 => A_neg_shifted(32),
                           C2 => n163, ZN => n237);
   U83 : AOI22_X1 port map( A1 => A_neg(32), A2 => n153, B1 => A_signal(32), B2
                           => n144, ZN => n238);
   U84 : NAND2_X1 port map( A1 => n244, A2 => n243, ZN => Y(35));
   U85 : AOI222_X1 port map( A1 => A_shifted(35), A2 => n179, B1 => 
                           zeroSignal(35), B2 => n170, C1 => A_neg_shifted(35),
                           C2 => n162, ZN => n243);
   U86 : AOI22_X1 port map( A1 => A_neg(35), A2 => n153, B1 => A_signal(35), B2
                           => n144, ZN => n244);
   U87 : NAND2_X1 port map( A1 => n240, A2 => n239, ZN => Y(33));
   U88 : AOI222_X1 port map( A1 => A_shifted(33), A2 => n179, B1 => 
                           zeroSignal(33), B2 => n170, C1 => A_neg_shifted(33),
                           C2 => n163, ZN => n239);
   U89 : AOI22_X1 port map( A1 => A_neg(33), A2 => n153, B1 => A_signal(33), B2
                           => n144, ZN => n240);
   U90 : NAND2_X1 port map( A1 => n248, A2 => n247, ZN => Y(37));
   U91 : AOI222_X1 port map( A1 => A_shifted(37), A2 => n179, B1 => 
                           zeroSignal(37), B2 => n170, C1 => A_neg_shifted(37),
                           C2 => n162, ZN => n247);
   U92 : AOI22_X1 port map( A1 => A_neg(37), A2 => n153, B1 => A_signal(37), B2
                           => n144, ZN => n248);
   U93 : NAND2_X1 port map( A1 => n214, A2 => n213, ZN => Y(21));
   U94 : AOI22_X1 port map( A1 => A_neg(21), A2 => n152, B1 => A_signal(21), B2
                           => n143, ZN => n214);
   U95 : AOI222_X1 port map( A1 => A_shifted(21), A2 => n178, B1 => 
                           zeroSignal(21), B2 => n169, C1 => A_neg_shifted(21),
                           C2 => n164, ZN => n213);
   U96 : NAND2_X1 port map( A1 => n252, A2 => n251, ZN => Y(39));
   U97 : AOI222_X1 port map( A1 => A_shifted(39), A2 => n179, B1 => 
                           zeroSignal(39), B2 => n170, C1 => A_neg_shifted(39),
                           C2 => n162, ZN => n251);
   U98 : AOI22_X1 port map( A1 => A_neg(39), A2 => n153, B1 => A_signal(39), B2
                           => n144, ZN => n252);
   U99 : NAND2_X1 port map( A1 => n234, A2 => n233, ZN => Y(30));
   U100 : AOI22_X1 port map( A1 => A_neg(30), A2 => n152, B1 => A_signal(30), 
                           B2 => n143, ZN => n234);
   U101 : AOI222_X1 port map( A1 => A_shifted(30), A2 => n178, B1 => 
                           zeroSignal(30), B2 => n169, C1 => A_neg_shifted(30),
                           C2 => n163, ZN => n233);
   U102 : NAND2_X1 port map( A1 => n246, A2 => n245, ZN => Y(36));
   U103 : AOI222_X1 port map( A1 => A_shifted(36), A2 => n179, B1 => 
                           zeroSignal(36), B2 => n170, C1 => A_neg_shifted(36),
                           C2 => n162, ZN => n245);
   U104 : AOI22_X1 port map( A1 => A_neg(36), A2 => n153, B1 => A_signal(36), 
                           B2 => n144, ZN => n246);
   U105 : NAND2_X1 port map( A1 => n250, A2 => n249, ZN => Y(38));
   U106 : AOI222_X1 port map( A1 => A_shifted(38), A2 => n179, B1 => 
                           zeroSignal(38), B2 => n170, C1 => A_neg_shifted(38),
                           C2 => n162, ZN => n249);
   U107 : AOI22_X1 port map( A1 => A_neg(38), A2 => n153, B1 => A_signal(38), 
                           B2 => n144, ZN => n250);
   U108 : NAND2_X1 port map( A1 => n258, A2 => n257, ZN => Y(41));
   U109 : AOI222_X1 port map( A1 => A_shifted(41), A2 => n179, B1 => 
                           zeroSignal(41), B2 => n170, C1 => A_neg_shifted(41),
                           C2 => n162, ZN => n257);
   U110 : AOI22_X1 port map( A1 => A_neg(41), A2 => n153, B1 => A_signal(41), 
                           B2 => n144, ZN => n258);
   U111 : NAND2_X1 port map( A1 => n242, A2 => n241, ZN => Y(34));
   U112 : AOI22_X1 port map( A1 => A_neg(34), A2 => n153, B1 => A_signal(34), 
                           B2 => n144, ZN => n242);
   U113 : AOI222_X1 port map( A1 => A_shifted(34), A2 => n179, B1 => 
                           zeroSignal(34), B2 => n170, C1 => A_neg_shifted(34),
                           C2 => n163, ZN => n241);
   U114 : NAND2_X1 port map( A1 => n260, A2 => n259, ZN => Y(42));
   U115 : AOI222_X1 port map( A1 => A_shifted(42), A2 => n180, B1 => 
                           zeroSignal(42), B2 => n171, C1 => A_neg_shifted(42),
                           C2 => n162, ZN => n259);
   U116 : AOI22_X1 port map( A1 => A_neg(42), A2 => n154, B1 => A_signal(42), 
                           B2 => n145, ZN => n260);
   U117 : NAND2_X1 port map( A1 => n262, A2 => n261, ZN => Y(43));
   U118 : AOI222_X1 port map( A1 => A_shifted(43), A2 => n180, B1 => 
                           zeroSignal(43), B2 => n171, C1 => A_neg_shifted(43),
                           C2 => n162, ZN => n261);
   U119 : AOI22_X1 port map( A1 => A_neg(43), A2 => n154, B1 => A_signal(43), 
                           B2 => n145, ZN => n262);
   U120 : NAND2_X1 port map( A1 => n264, A2 => n263, ZN => Y(44));
   U121 : AOI222_X1 port map( A1 => A_shifted(44), A2 => n180, B1 => 
                           zeroSignal(44), B2 => n171, C1 => A_neg_shifted(44),
                           C2 => n162, ZN => n263);
   U122 : AOI22_X1 port map( A1 => A_neg(44), A2 => n154, B1 => A_signal(44), 
                           B2 => n145, ZN => n264);
   U123 : NAND2_X1 port map( A1 => n266, A2 => n265, ZN => Y(45));
   U124 : AOI222_X1 port map( A1 => A_shifted(45), A2 => n180, B1 => 
                           zeroSignal(45), B2 => n171, C1 => A_neg_shifted(45),
                           C2 => n162, ZN => n265);
   U125 : AOI22_X1 port map( A1 => A_neg(45), A2 => n154, B1 => A_signal(45), 
                           B2 => n145, ZN => n266);
   U126 : NAND2_X1 port map( A1 => n274, A2 => n273, ZN => Y(49));
   U127 : AOI222_X1 port map( A1 => A_shifted(49), A2 => n180, B1 => 
                           zeroSignal(49), B2 => n171, C1 => A_neg_shifted(49),
                           C2 => n161, ZN => n273);
   U128 : AOI22_X1 port map( A1 => A_neg(49), A2 => n154, B1 => A_signal(49), 
                           B2 => n145, ZN => n274);
   U129 : NAND2_X1 port map( A1 => n268, A2 => n267, ZN => Y(46));
   U130 : AOI222_X1 port map( A1 => A_shifted(46), A2 => n180, B1 => 
                           zeroSignal(46), B2 => n171, C1 => A_neg_shifted(46),
                           C2 => n161, ZN => n267);
   U131 : AOI22_X1 port map( A1 => A_neg(46), A2 => n154, B1 => A_signal(46), 
                           B2 => n145, ZN => n268);
   U132 : NAND2_X1 port map( A1 => n256, A2 => n255, ZN => Y(40));
   U133 : AOI22_X1 port map( A1 => A_neg(40), A2 => n153, B1 => A_signal(40), 
                           B2 => n144, ZN => n256);
   U134 : AOI222_X1 port map( A1 => A_shifted(40), A2 => n179, B1 => 
                           zeroSignal(40), B2 => n170, C1 => A_neg_shifted(40),
                           C2 => n162, ZN => n255);
   U135 : NAND2_X1 port map( A1 => n216, A2 => n215, ZN => Y(22));
   U136 : AOI222_X1 port map( A1 => A_shifted(22), A2 => n178, B1 => 
                           zeroSignal(22), B2 => n169, C1 => A_neg_shifted(22),
                           C2 => n164, ZN => n215);
   U137 : AOI22_X1 port map( A1 => A_neg(22), A2 => n152, B1 => A_signal(22), 
                           B2 => n143, ZN => n216);
   U138 : NAND2_X1 port map( A1 => n270, A2 => n269, ZN => Y(47));
   U139 : AOI222_X1 port map( A1 => A_shifted(47), A2 => n180, B1 => 
                           zeroSignal(47), B2 => n171, C1 => A_neg_shifted(47),
                           C2 => n161, ZN => n269);
   U140 : AOI22_X1 port map( A1 => A_neg(47), A2 => n154, B1 => A_signal(47), 
                           B2 => n145, ZN => n270);
   U141 : NAND2_X1 port map( A1 => n218, A2 => n217, ZN => Y(23));
   U142 : AOI222_X1 port map( A1 => A_shifted(23), A2 => n178, B1 => 
                           zeroSignal(23), B2 => n169, C1 => A_neg_shifted(23),
                           C2 => n164, ZN => n217);
   U143 : AOI22_X1 port map( A1 => A_neg(23), A2 => n152, B1 => A_signal(23), 
                           B2 => n143, ZN => n218);
   U144 : NAND2_X1 port map( A1 => n220, A2 => n219, ZN => Y(24));
   U145 : AOI222_X1 port map( A1 => A_shifted(24), A2 => n178, B1 => 
                           zeroSignal(24), B2 => n169, C1 => A_neg_shifted(24),
                           C2 => n163, ZN => n219);
   U146 : AOI22_X1 port map( A1 => A_neg(24), A2 => n152, B1 => A_signal(24), 
                           B2 => n143, ZN => n220);
   U147 : NAND2_X1 port map( A1 => n272, A2 => n271, ZN => Y(48));
   U148 : AOI222_X1 port map( A1 => A_shifted(48), A2 => n180, B1 => 
                           zeroSignal(48), B2 => n171, C1 => A_neg_shifted(48),
                           C2 => n161, ZN => n271);
   U149 : AOI22_X1 port map( A1 => A_neg(48), A2 => n154, B1 => A_signal(48), 
                           B2 => n145, ZN => n272);
   U150 : NAND2_X1 port map( A1 => n222, A2 => n221, ZN => Y(25));
   U151 : AOI222_X1 port map( A1 => A_shifted(25), A2 => n178, B1 => 
                           zeroSignal(25), B2 => n169, C1 => A_neg_shifted(25),
                           C2 => n163, ZN => n221);
   U152 : AOI22_X1 port map( A1 => A_neg(25), A2 => n152, B1 => A_signal(25), 
                           B2 => n143, ZN => n222);
   U153 : NAND2_X1 port map( A1 => n278, A2 => n277, ZN => Y(50));
   U154 : AOI22_X1 port map( A1 => A_neg(50), A2 => n154, B1 => A_signal(50), 
                           B2 => n145, ZN => n278);
   U155 : AOI222_X1 port map( A1 => A_shifted(50), A2 => n180, B1 => 
                           zeroSignal(50), B2 => n171, C1 => A_neg_shifted(50),
                           C2 => n161, ZN => n277);
   U156 : NAND2_X1 port map( A1 => n280, A2 => n279, ZN => Y(51));
   U157 : AOI222_X1 port map( A1 => A_shifted(51), A2 => n180, B1 => 
                           zeroSignal(51), B2 => n171, C1 => A_neg_shifted(51),
                           C2 => n161, ZN => n279);
   U158 : AOI22_X1 port map( A1 => A_neg(51), A2 => n154, B1 => A_signal(51), 
                           B2 => n145, ZN => n280);
   U159 : NAND2_X1 port map( A1 => n282, A2 => n281, ZN => Y(52));
   U160 : AOI222_X1 port map( A1 => A_shifted(52), A2 => n180, B1 => 
                           zeroSignal(52), B2 => n171, C1 => A_neg_shifted(52),
                           C2 => n161, ZN => n281);
   U161 : AOI22_X1 port map( A1 => A_neg(52), A2 => n154, B1 => A_signal(52), 
                           B2 => n145, ZN => n282);
   U162 : NAND2_X1 port map( A1 => n284, A2 => n283, ZN => Y(53));
   U163 : AOI22_X1 port map( A1 => A_neg(53), A2 => n155, B1 => A_signal(53), 
                           B2 => n146, ZN => n284);
   U164 : AOI222_X1 port map( A1 => A_shifted(53), A2 => n181, B1 => 
                           zeroSignal(53), B2 => n172, C1 => A_neg_shifted(53),
                           C2 => n161, ZN => n283);
   U165 : NAND2_X1 port map( A1 => n288, A2 => n287, ZN => Y(55));
   U166 : AOI222_X1 port map( A1 => A_shifted(55), A2 => n181, B1 => 
                           zeroSignal(55), B2 => n172, C1 => A_neg_shifted(55),
                           C2 => n161, ZN => n287);
   U167 : AOI22_X1 port map( A1 => A_neg(55), A2 => n155, B1 => A_signal(55), 
                           B2 => n146, ZN => n288);
   U168 : NAND2_X1 port map( A1 => n290, A2 => n289, ZN => Y(56));
   U169 : AOI222_X1 port map( A1 => A_shifted(56), A2 => n181, B1 => 
                           zeroSignal(56), B2 => n172, C1 => A_neg_shifted(56),
                           C2 => n161, ZN => n289);
   U170 : AOI22_X1 port map( A1 => A_neg(56), A2 => n155, B1 => A_signal(56), 
                           B2 => n146, ZN => n290);
   U171 : NAND2_X1 port map( A1 => n286, A2 => n285, ZN => Y(54));
   U172 : AOI222_X1 port map( A1 => A_shifted(54), A2 => n181, B1 => 
                           zeroSignal(54), B2 => n172, C1 => A_neg_shifted(54),
                           C2 => n161, ZN => n285);
   U173 : AOI22_X1 port map( A1 => A_neg(54), A2 => n155, B1 => A_signal(54), 
                           B2 => n146, ZN => n286);
   U174 : NAND2_X1 port map( A1 => n292, A2 => n291, ZN => Y(57));
   U175 : AOI22_X1 port map( A1 => A_neg(57), A2 => n155, B1 => A_signal(57), 
                           B2 => n146, ZN => n292);
   U176 : AOI222_X1 port map( A1 => A_shifted(57), A2 => n181, B1 => 
                           zeroSignal(57), B2 => n172, C1 => A_neg_shifted(57),
                           C2 => n160, ZN => n291);
   U177 : NAND2_X1 port map( A1 => n306, A2 => n305, ZN => Y(63));
   U178 : NAND2_X1 port map( A1 => n304, A2 => n303, ZN => Y(62));
   U179 : AOI222_X1 port map( A1 => A_shifted(62), A2 => n181, B1 => 
                           zeroSignal(62), B2 => n172, C1 => A_neg_shifted(62),
                           C2 => n160, ZN => n303);
   U180 : NAND2_X1 port map( A1 => n296, A2 => n295, ZN => Y(59));
   U181 : AOI222_X1 port map( A1 => A_shifted(59), A2 => n181, B1 => 
                           zeroSignal(59), B2 => n172, C1 => A_neg_shifted(59),
                           C2 => n160, ZN => n295);
   U182 : AOI22_X1 port map( A1 => A_neg(59), A2 => n155, B1 => A_signal(59), 
                           B2 => n146, ZN => n296);
   U183 : NAND2_X1 port map( A1 => n300, A2 => n299, ZN => Y(60));
   U184 : AOI222_X1 port map( A1 => A_shifted(60), A2 => n181, B1 => 
                           zeroSignal(60), B2 => n172, C1 => A_neg_shifted(60),
                           C2 => n160, ZN => n299);
   U185 : NAND2_X1 port map( A1 => n302, A2 => n301, ZN => Y(61));
   U186 : AOI22_X1 port map( A1 => A_neg(61), A2 => n155, B1 => A_signal(61), 
                           B2 => n146, ZN => n302);
   U187 : NAND2_X1 port map( A1 => n294, A2 => n293, ZN => Y(58));
   U188 : AOI22_X1 port map( A1 => A_neg(58), A2 => n155, B1 => A_signal(58), 
                           B2 => n146, ZN => n294);
   U189 : AOI222_X1 port map( A1 => A_shifted(58), A2 => n181, B1 => 
                           zeroSignal(58), B2 => n172, C1 => A_neg_shifted(58),
                           C2 => n160, ZN => n293);
   U190 : NAND2_X1 port map( A1 => n188, A2 => n187, ZN => Y(0));
   U191 : AOI22_X1 port map( A1 => A_neg(0), A2 => n151, B1 => A_signal(0), B2 
                           => n142, ZN => n188);
   U192 : AOI222_X1 port map( A1 => A_shifted(0), A2 => n177, B1 => 
                           zeroSignal(0), B2 => n168, C1 => A_neg_shifted(0), 
                           C2 => n165, ZN => n187);
   U193 : NAND2_X1 port map( A1 => n210, A2 => n209, ZN => Y(1));
   U194 : AOI22_X1 port map( A1 => A_neg(1), A2 => n151, B1 => A_signal(1), B2 
                           => n142, ZN => n210);
   U195 : AOI222_X1 port map( A1 => A_shifted(1), A2 => n177, B1 => 
                           zeroSignal(1), B2 => n168, C1 => A_neg_shifted(1), 
                           C2 => n164, ZN => n209);
   U196 : NAND2_X1 port map( A1 => n232, A2 => n231, ZN => Y(2));
   U197 : AOI22_X1 port map( A1 => A_neg(2), A2 => n152, B1 => A_signal(2), B2 
                           => n143, ZN => n232);
   U198 : AOI222_X1 port map( A1 => A_shifted(2), A2 => n178, B1 => 
                           zeroSignal(2), B2 => n169, C1 => A_neg_shifted(2), 
                           C2 => n163, ZN => n231);
   U199 : NAND2_X1 port map( A1 => n254, A2 => n253, ZN => Y(3));
   U200 : AOI22_X1 port map( A1 => A_neg(3), A2 => n153, B1 => A_signal(3), B2 
                           => n144, ZN => n254);
   U201 : AOI222_X1 port map( A1 => A_shifted(3), A2 => n179, B1 => 
                           zeroSignal(3), B2 => n170, C1 => A_neg_shifted(3), 
                           C2 => n162, ZN => n253);
   U202 : NAND2_X1 port map( A1 => n276, A2 => n275, ZN => Y(4));
   U203 : AOI22_X1 port map( A1 => A_neg(4), A2 => n154, B1 => A_signal(4), B2 
                           => n145, ZN => n276);
   U204 : AOI222_X1 port map( A1 => A_shifted(4), A2 => n180, B1 => 
                           zeroSignal(4), B2 => n171, C1 => A_neg_shifted(4), 
                           C2 => n161, ZN => n275);
   U205 : NAND2_X1 port map( A1 => n298, A2 => n297, ZN => Y(5));
   U206 : AOI22_X1 port map( A1 => A_neg(5), A2 => n155, B1 => A_signal(5), B2 
                           => n146, ZN => n298);
   U207 : AOI222_X1 port map( A1 => A_shifted(5), A2 => n181, B1 => 
                           zeroSignal(5), B2 => n172, C1 => A_neg_shifted(5), 
                           C2 => n160, ZN => n297);
   U208 : NAND2_X1 port map( A1 => n308, A2 => n307, ZN => Y(6));
   U209 : AOI22_X1 port map( A1 => A_neg(6), A2 => n156, B1 => A_signal(6), B2 
                           => n147, ZN => n308);
   U210 : AOI222_X1 port map( A1 => A_shifted(6), A2 => n182, B1 => 
                           zeroSignal(6), B2 => n173, C1 => A_neg_shifted(6), 
                           C2 => n160, ZN => n307);
   U211 : NAND2_X1 port map( A1 => n310, A2 => n309, ZN => Y(7));
   U212 : AOI22_X1 port map( A1 => A_neg(7), A2 => n156, B1 => A_signal(7), B2 
                           => n147, ZN => n310);
   U213 : AOI222_X1 port map( A1 => A_shifted(7), A2 => n182, B1 => 
                           zeroSignal(7), B2 => n173, C1 => A_neg_shifted(7), 
                           C2 => n160, ZN => n309);
   U214 : NAND2_X1 port map( A1 => n312, A2 => n311, ZN => Y(8));
   U215 : AOI22_X1 port map( A1 => A_neg(8), A2 => n156, B1 => A_signal(8), B2 
                           => n147, ZN => n312);
   U216 : AOI222_X1 port map( A1 => A_shifted(8), A2 => n182, B1 => 
                           zeroSignal(8), B2 => n173, C1 => A_neg_shifted(8), 
                           C2 => n160, ZN => n311);
   U217 : NAND2_X1 port map( A1 => n318, A2 => n317, ZN => Y(9));
   U218 : AOI22_X1 port map( A1 => A_neg(9), A2 => n156, B1 => A_signal(9), B2 
                           => n147, ZN => n318);
   U219 : AOI222_X1 port map( A1 => A_shifted(9), A2 => n182, B1 => 
                           zeroSignal(9), B2 => n173, C1 => A_neg_shifted(9), 
                           C2 => n160, ZN => n317);
   U220 : NAND2_X1 port map( A1 => n190, A2 => n189, ZN => Y(10));
   U221 : AOI22_X1 port map( A1 => A_neg(10), A2 => n151, B1 => A_signal(10), 
                           B2 => n142, ZN => n190);
   U222 : AOI222_X1 port map( A1 => A_shifted(10), A2 => n177, B1 => 
                           zeroSignal(10), B2 => n168, C1 => A_neg_shifted(10),
                           C2 => n165, ZN => n189);
   U223 : NAND2_X1 port map( A1 => n192, A2 => n191, ZN => Y(11));
   U224 : AOI22_X1 port map( A1 => A_neg(11), A2 => n151, B1 => A_signal(11), 
                           B2 => n142, ZN => n192);
   U225 : AOI222_X1 port map( A1 => A_shifted(11), A2 => n177, B1 => 
                           zeroSignal(11), B2 => n168, C1 => A_neg_shifted(11),
                           C2 => n165, ZN => n191);
   U226 : NAND2_X1 port map( A1 => n194, A2 => n193, ZN => Y(12));
   U227 : AOI22_X1 port map( A1 => A_neg(12), A2 => n151, B1 => A_signal(12), 
                           B2 => n142, ZN => n194);
   U228 : AOI222_X1 port map( A1 => A_shifted(12), A2 => n177, B1 => 
                           zeroSignal(12), B2 => n168, C1 => A_neg_shifted(12),
                           C2 => n165, ZN => n193);
   U229 : NAND2_X1 port map( A1 => n196, A2 => n195, ZN => Y(13));
   U230 : AOI22_X1 port map( A1 => A_neg(13), A2 => n151, B1 => A_signal(13), 
                           B2 => n142, ZN => n196);
   U231 : AOI222_X1 port map( A1 => A_shifted(13), A2 => n177, B1 => 
                           zeroSignal(13), B2 => n168, C1 => A_neg_shifted(13),
                           C2 => n164, ZN => n195);
   U232 : NAND2_X1 port map( A1 => n198, A2 => n197, ZN => Y(14));
   U233 : AOI22_X1 port map( A1 => A_neg(14), A2 => n151, B1 => A_signal(14), 
                           B2 => n142, ZN => n198);
   U234 : AOI222_X1 port map( A1 => A_shifted(14), A2 => n177, B1 => 
                           zeroSignal(14), B2 => n168, C1 => A_neg_shifted(14),
                           C2 => n164, ZN => n197);
   U235 : NAND2_X1 port map( A1 => n200, A2 => n199, ZN => Y(15));
   U236 : AOI22_X1 port map( A1 => A_neg(15), A2 => n151, B1 => A_signal(15), 
                           B2 => n142, ZN => n200);
   U237 : AOI222_X1 port map( A1 => A_shifted(15), A2 => n177, B1 => 
                           zeroSignal(15), B2 => n168, C1 => A_neg_shifted(15),
                           C2 => n164, ZN => n199);
   U238 : AOI222_X1 port map( A1 => A_shifted(63), A2 => n181, B1 => 
                           zeroSignal(63), B2 => n172, C1 => A_neg_shifted(63),
                           C2 => n160, ZN => n305);
   U239 : AOI22_X1 port map( A1 => A_neg(62), A2 => n155, B1 => A_signal(62), 
                           B2 => n146, ZN => n304);
   U240 : AOI22_X1 port map( A1 => A_neg(63), A2 => n155, B1 => A_signal(63), 
                           B2 => n146, ZN => n306);
   U241 : AOI222_X1 port map( A1 => A_shifted(61), A2 => n181, B1 => 
                           zeroSignal(61), B2 => n172, C1 => A_neg_shifted(61),
                           C2 => n160, ZN => n301);
   U242 : AOI22_X1 port map( A1 => A_neg(60), A2 => n155, B1 => A_signal(60), 
                           B2 => n146, ZN => n300);
   U243 : AOI222_X1 port map( A1 => A_shifted(17), A2 => n177, B1 => 
                           zeroSignal(17), B2 => n168, C1 => A_neg_shifted(17),
                           C2 => n164, ZN => n203);
   U244 : AOI22_X1 port map( A1 => A_neg(16), A2 => n151, B1 => A_signal(16), 
                           B2 => n142, ZN => n202);

end SYN_BEHAVIORAL_2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity MUX51_MuxNbit64_23 is

   port( zeroSignal, A_signal, A_neg, A_shifted, A_neg_shifted : in 
         std_logic_vector (63 downto 0);  Sel : in std_logic_vector (2 downto 
         0);  Y : out std_logic_vector (63 downto 0));

end MUX51_MuxNbit64_23;

architecture SYN_BEHAVIORAL_2 of MUX51_MuxNbit64_23 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, 
      n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, 
      n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, 
      n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, 
      n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, 
      n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, 
      n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, 
      n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, 
      n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, 
      n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, 
      n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, 
      n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, 
      n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, 
      n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, 
      n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, 
      n320 : std_logic;

begin
   
   U1 : AND3_X1 port map( A1 => n319, A2 => n320, A3 => Sel(2), ZN => n141);
   U2 : BUF_X1 port map( A => n141, Z => n166);
   U3 : BUF_X1 port map( A => n185, Z => n184);
   U4 : BUF_X1 port map( A => n159, Z => n158);
   U5 : BUF_X1 port map( A => n150, Z => n149);
   U6 : BUF_X1 port map( A => n141, Z => n167);
   U7 : BUF_X1 port map( A => n185, Z => n183);
   U8 : BUF_X1 port map( A => n159, Z => n157);
   U9 : BUF_X1 port map( A => n150, Z => n148);
   U10 : BUF_X1 port map( A => n176, Z => n175);
   U11 : BUF_X1 port map( A => n176, Z => n174);
   U12 : BUF_X1 port map( A => n158, Z => n151);
   U13 : BUF_X1 port map( A => n184, Z => n177);
   U14 : BUF_X1 port map( A => n149, Z => n142);
   U15 : BUF_X1 port map( A => n166, Z => n164);
   U16 : BUF_X1 port map( A => n184, Z => n178);
   U17 : BUF_X1 port map( A => n158, Z => n152);
   U18 : BUF_X1 port map( A => n149, Z => n143);
   U19 : BUF_X1 port map( A => n166, Z => n163);
   U20 : BUF_X1 port map( A => n184, Z => n179);
   U21 : BUF_X1 port map( A => n158, Z => n153);
   U22 : BUF_X1 port map( A => n149, Z => n144);
   U23 : BUF_X1 port map( A => n167, Z => n162);
   U24 : BUF_X1 port map( A => n183, Z => n180);
   U25 : BUF_X1 port map( A => n157, Z => n154);
   U26 : BUF_X1 port map( A => n148, Z => n145);
   U27 : BUF_X1 port map( A => n167, Z => n161);
   U28 : BUF_X1 port map( A => n183, Z => n181);
   U29 : BUF_X1 port map( A => n157, Z => n155);
   U30 : BUF_X1 port map( A => n148, Z => n146);
   U31 : BUF_X1 port map( A => n167, Z => n160);
   U32 : BUF_X1 port map( A => n175, Z => n169);
   U33 : BUF_X1 port map( A => n175, Z => n170);
   U34 : BUF_X1 port map( A => n174, Z => n171);
   U35 : BUF_X1 port map( A => n175, Z => n168);
   U36 : BUF_X1 port map( A => n174, Z => n172);
   U37 : BUF_X1 port map( A => n166, Z => n165);
   U38 : BUF_X1 port map( A => n157, Z => n156);
   U39 : BUF_X1 port map( A => n148, Z => n147);
   U40 : BUF_X1 port map( A => n174, Z => n173);
   U41 : BUF_X1 port map( A => n183, Z => n182);
   U42 : INV_X1 port map( A => Sel(1), ZN => n320);
   U43 : BUF_X1 port map( A => n314, Z => n159);
   U44 : NOR3_X1 port map( A1 => Sel(0), A2 => Sel(2), A3 => n320, ZN => n314);
   U45 : BUF_X1 port map( A => n316, Z => n185);
   U46 : NOR3_X1 port map( A1 => n319, A2 => Sel(2), A3 => n320, ZN => n316);
   U47 : BUF_X1 port map( A => n313, Z => n150);
   U48 : NOR3_X1 port map( A1 => Sel(1), A2 => Sel(2), A3 => n319, ZN => n313);
   U49 : INV_X1 port map( A => Sel(0), ZN => n319);
   U50 : BUF_X1 port map( A => n315, Z => n176);
   U51 : NOR2_X1 port map( A1 => n165, A2 => n186, ZN => n315);
   U52 : AOI21_X1 port map( B1 => n319, B2 => n320, A => Sel(2), ZN => n186);
   U53 : NAND2_X1 port map( A1 => n208, A2 => n207, ZN => Y(19));
   U54 : AOI22_X1 port map( A1 => A_neg(19), A2 => n151, B1 => A_signal(19), B2
                           => n142, ZN => n208);
   U55 : NAND2_X1 port map( A1 => n206, A2 => n205, ZN => Y(18));
   U56 : AOI222_X1 port map( A1 => A_shifted(18), A2 => n177, B1 => 
                           zeroSignal(18), B2 => n168, C1 => A_neg_shifted(18),
                           C2 => n164, ZN => n205);
   U57 : NAND2_X1 port map( A1 => n212, A2 => n211, ZN => Y(20));
   U58 : AOI22_X1 port map( A1 => A_neg(20), A2 => n152, B1 => A_signal(20), B2
                           => n143, ZN => n212);
   U59 : AOI222_X1 port map( A1 => A_shifted(20), A2 => n178, B1 => 
                           zeroSignal(20), B2 => n169, C1 => A_neg_shifted(20),
                           C2 => n164, ZN => n211);
   U60 : NAND2_X1 port map( A1 => n214, A2 => n213, ZN => Y(21));
   U61 : AOI22_X1 port map( A1 => A_neg(21), A2 => n152, B1 => A_signal(21), B2
                           => n143, ZN => n214);
   U62 : AOI222_X1 port map( A1 => A_shifted(21), A2 => n178, B1 => 
                           zeroSignal(21), B2 => n169, C1 => A_neg_shifted(21),
                           C2 => n164, ZN => n213);
   U63 : NAND2_X1 port map( A1 => n216, A2 => n215, ZN => Y(22));
   U64 : AOI22_X1 port map( A1 => A_neg(22), A2 => n152, B1 => A_signal(22), B2
                           => n143, ZN => n216);
   U65 : AOI222_X1 port map( A1 => A_shifted(22), A2 => n178, B1 => 
                           zeroSignal(22), B2 => n169, C1 => A_neg_shifted(22),
                           C2 => n164, ZN => n215);
   U66 : NAND2_X1 port map( A1 => n228, A2 => n227, ZN => Y(28));
   U67 : AOI222_X1 port map( A1 => A_shifted(28), A2 => n178, B1 => 
                           zeroSignal(28), B2 => n169, C1 => A_neg_shifted(28),
                           C2 => n163, ZN => n227);
   U68 : AOI22_X1 port map( A1 => A_neg(28), A2 => n152, B1 => A_signal(28), B2
                           => n143, ZN => n228);
   U69 : NAND2_X1 port map( A1 => n236, A2 => n235, ZN => Y(31));
   U70 : AOI222_X1 port map( A1 => A_shifted(31), A2 => n179, B1 => 
                           zeroSignal(31), B2 => n170, C1 => A_neg_shifted(31),
                           C2 => n163, ZN => n235);
   U71 : AOI22_X1 port map( A1 => A_neg(31), A2 => n153, B1 => A_signal(31), B2
                           => n144, ZN => n236);
   U72 : NAND2_X1 port map( A1 => n230, A2 => n229, ZN => Y(29));
   U73 : AOI222_X1 port map( A1 => A_shifted(29), A2 => n178, B1 => 
                           zeroSignal(29), B2 => n169, C1 => A_neg_shifted(29),
                           C2 => n163, ZN => n229);
   U74 : AOI22_X1 port map( A1 => A_neg(29), A2 => n152, B1 => A_signal(29), B2
                           => n143, ZN => n230);
   U75 : NAND2_X1 port map( A1 => n234, A2 => n233, ZN => Y(30));
   U76 : AOI222_X1 port map( A1 => A_shifted(30), A2 => n178, B1 => 
                           zeroSignal(30), B2 => n169, C1 => A_neg_shifted(30),
                           C2 => n163, ZN => n233);
   U77 : AOI22_X1 port map( A1 => A_neg(30), A2 => n152, B1 => A_signal(30), B2
                           => n143, ZN => n234);
   U78 : NAND2_X1 port map( A1 => n242, A2 => n241, ZN => Y(34));
   U79 : AOI222_X1 port map( A1 => A_shifted(34), A2 => n179, B1 => 
                           zeroSignal(34), B2 => n170, C1 => A_neg_shifted(34),
                           C2 => n163, ZN => n241);
   U80 : AOI22_X1 port map( A1 => A_neg(34), A2 => n153, B1 => A_signal(34), B2
                           => n144, ZN => n242);
   U81 : NAND2_X1 port map( A1 => n244, A2 => n243, ZN => Y(35));
   U82 : AOI222_X1 port map( A1 => A_shifted(35), A2 => n179, B1 => 
                           zeroSignal(35), B2 => n170, C1 => A_neg_shifted(35),
                           C2 => n162, ZN => n243);
   U83 : AOI22_X1 port map( A1 => A_neg(35), A2 => n153, B1 => A_signal(35), B2
                           => n144, ZN => n244);
   U84 : NAND2_X1 port map( A1 => n240, A2 => n239, ZN => Y(33));
   U85 : AOI222_X1 port map( A1 => A_shifted(33), A2 => n179, B1 => 
                           zeroSignal(33), B2 => n170, C1 => A_neg_shifted(33),
                           C2 => n163, ZN => n239);
   U86 : AOI22_X1 port map( A1 => A_neg(33), A2 => n153, B1 => A_signal(33), B2
                           => n144, ZN => n240);
   U87 : NAND2_X1 port map( A1 => n252, A2 => n251, ZN => Y(39));
   U88 : AOI222_X1 port map( A1 => A_shifted(39), A2 => n179, B1 => 
                           zeroSignal(39), B2 => n170, C1 => A_neg_shifted(39),
                           C2 => n162, ZN => n251);
   U89 : AOI22_X1 port map( A1 => A_neg(39), A2 => n153, B1 => A_signal(39), B2
                           => n144, ZN => n252);
   U90 : NAND2_X1 port map( A1 => n248, A2 => n247, ZN => Y(37));
   U91 : AOI222_X1 port map( A1 => A_shifted(37), A2 => n179, B1 => 
                           zeroSignal(37), B2 => n170, C1 => A_neg_shifted(37),
                           C2 => n162, ZN => n247);
   U92 : AOI22_X1 port map( A1 => A_neg(37), A2 => n153, B1 => A_signal(37), B2
                           => n144, ZN => n248);
   U93 : NAND2_X1 port map( A1 => n250, A2 => n249, ZN => Y(38));
   U94 : AOI222_X1 port map( A1 => A_shifted(38), A2 => n179, B1 => 
                           zeroSignal(38), B2 => n170, C1 => A_neg_shifted(38),
                           C2 => n162, ZN => n249);
   U95 : AOI22_X1 port map( A1 => A_neg(38), A2 => n153, B1 => A_signal(38), B2
                           => n144, ZN => n250);
   U96 : NAND2_X1 port map( A1 => n256, A2 => n255, ZN => Y(40));
   U97 : AOI222_X1 port map( A1 => A_shifted(40), A2 => n179, B1 => 
                           zeroSignal(40), B2 => n170, C1 => A_neg_shifted(40),
                           C2 => n162, ZN => n255);
   U98 : AOI22_X1 port map( A1 => A_neg(40), A2 => n153, B1 => A_signal(40), B2
                           => n144, ZN => n256);
   U99 : NAND2_X1 port map( A1 => n218, A2 => n217, ZN => Y(23));
   U100 : AOI22_X1 port map( A1 => A_neg(23), A2 => n152, B1 => A_signal(23), 
                           B2 => n143, ZN => n218);
   U101 : AOI222_X1 port map( A1 => A_shifted(23), A2 => n178, B1 => 
                           zeroSignal(23), B2 => n169, C1 => A_neg_shifted(23),
                           C2 => n164, ZN => n217);
   U102 : NAND2_X1 port map( A1 => n238, A2 => n237, ZN => Y(32));
   U103 : AOI22_X1 port map( A1 => A_neg(32), A2 => n153, B1 => A_signal(32), 
                           B2 => n144, ZN => n238);
   U104 : AOI222_X1 port map( A1 => A_shifted(32), A2 => n179, B1 => 
                           zeroSignal(32), B2 => n170, C1 => A_neg_shifted(32),
                           C2 => n163, ZN => n237);
   U105 : NAND2_X1 port map( A1 => n258, A2 => n257, ZN => Y(41));
   U106 : AOI222_X1 port map( A1 => A_shifted(41), A2 => n179, B1 => 
                           zeroSignal(41), B2 => n170, C1 => A_neg_shifted(41),
                           C2 => n162, ZN => n257);
   U107 : AOI22_X1 port map( A1 => A_neg(41), A2 => n153, B1 => A_signal(41), 
                           B2 => n144, ZN => n258);
   U108 : NAND2_X1 port map( A1 => n264, A2 => n263, ZN => Y(44));
   U109 : AOI222_X1 port map( A1 => A_shifted(44), A2 => n180, B1 => 
                           zeroSignal(44), B2 => n171, C1 => A_neg_shifted(44),
                           C2 => n162, ZN => n263);
   U110 : AOI22_X1 port map( A1 => A_neg(44), A2 => n154, B1 => A_signal(44), 
                           B2 => n145, ZN => n264);
   U111 : NAND2_X1 port map( A1 => n266, A2 => n265, ZN => Y(45));
   U112 : AOI222_X1 port map( A1 => A_shifted(45), A2 => n180, B1 => 
                           zeroSignal(45), B2 => n171, C1 => A_neg_shifted(45),
                           C2 => n162, ZN => n265);
   U113 : AOI22_X1 port map( A1 => A_neg(45), A2 => n154, B1 => A_signal(45), 
                           B2 => n145, ZN => n266);
   U114 : NAND2_X1 port map( A1 => n246, A2 => n245, ZN => Y(36));
   U115 : AOI22_X1 port map( A1 => A_neg(36), A2 => n153, B1 => A_signal(36), 
                           B2 => n144, ZN => n246);
   U116 : AOI222_X1 port map( A1 => A_shifted(36), A2 => n179, B1 => 
                           zeroSignal(36), B2 => n170, C1 => A_neg_shifted(36),
                           C2 => n162, ZN => n245);
   U117 : NAND2_X1 port map( A1 => n262, A2 => n261, ZN => Y(43));
   U118 : AOI222_X1 port map( A1 => A_shifted(43), A2 => n180, B1 => 
                           zeroSignal(43), B2 => n171, C1 => A_neg_shifted(43),
                           C2 => n162, ZN => n261);
   U119 : AOI22_X1 port map( A1 => A_neg(43), A2 => n154, B1 => A_signal(43), 
                           B2 => n145, ZN => n262);
   U120 : NAND2_X1 port map( A1 => n280, A2 => n279, ZN => Y(51));
   U121 : AOI222_X1 port map( A1 => A_shifted(51), A2 => n180, B1 => 
                           zeroSignal(51), B2 => n171, C1 => A_neg_shifted(51),
                           C2 => n161, ZN => n279);
   U122 : AOI22_X1 port map( A1 => A_neg(51), A2 => n154, B1 => A_signal(51), 
                           B2 => n145, ZN => n280);
   U123 : NAND2_X1 port map( A1 => n268, A2 => n267, ZN => Y(46));
   U124 : AOI222_X1 port map( A1 => A_shifted(46), A2 => n180, B1 => 
                           zeroSignal(46), B2 => n171, C1 => A_neg_shifted(46),
                           C2 => n161, ZN => n267);
   U125 : AOI22_X1 port map( A1 => A_neg(46), A2 => n154, B1 => A_signal(46), 
                           B2 => n145, ZN => n268);
   U126 : NAND2_X1 port map( A1 => n260, A2 => n259, ZN => Y(42));
   U127 : AOI22_X1 port map( A1 => A_neg(42), A2 => n154, B1 => A_signal(42), 
                           B2 => n145, ZN => n260);
   U128 : AOI222_X1 port map( A1 => A_shifted(42), A2 => n180, B1 => 
                           zeroSignal(42), B2 => n171, C1 => A_neg_shifted(42),
                           C2 => n162, ZN => n259);
   U129 : NAND2_X1 port map( A1 => n270, A2 => n269, ZN => Y(47));
   U130 : AOI222_X1 port map( A1 => A_shifted(47), A2 => n180, B1 => 
                           zeroSignal(47), B2 => n171, C1 => A_neg_shifted(47),
                           C2 => n161, ZN => n269);
   U131 : AOI22_X1 port map( A1 => A_neg(47), A2 => n154, B1 => A_signal(47), 
                           B2 => n145, ZN => n270);
   U132 : NAND2_X1 port map( A1 => n274, A2 => n273, ZN => Y(49));
   U133 : AOI222_X1 port map( A1 => A_shifted(49), A2 => n180, B1 => 
                           zeroSignal(49), B2 => n171, C1 => A_neg_shifted(49),
                           C2 => n161, ZN => n273);
   U134 : AOI22_X1 port map( A1 => A_neg(49), A2 => n154, B1 => A_signal(49), 
                           B2 => n145, ZN => n274);
   U135 : NAND2_X1 port map( A1 => n272, A2 => n271, ZN => Y(48));
   U136 : AOI222_X1 port map( A1 => A_shifted(48), A2 => n180, B1 => 
                           zeroSignal(48), B2 => n171, C1 => A_neg_shifted(48),
                           C2 => n161, ZN => n271);
   U137 : AOI22_X1 port map( A1 => A_neg(48), A2 => n154, B1 => A_signal(48), 
                           B2 => n145, ZN => n272);
   U138 : NAND2_X1 port map( A1 => n220, A2 => n219, ZN => Y(24));
   U139 : AOI222_X1 port map( A1 => A_shifted(24), A2 => n178, B1 => 
                           zeroSignal(24), B2 => n169, C1 => A_neg_shifted(24),
                           C2 => n163, ZN => n219);
   U140 : AOI22_X1 port map( A1 => A_neg(24), A2 => n152, B1 => A_signal(24), 
                           B2 => n143, ZN => n220);
   U141 : NAND2_X1 port map( A1 => n222, A2 => n221, ZN => Y(25));
   U142 : AOI222_X1 port map( A1 => A_shifted(25), A2 => n178, B1 => 
                           zeroSignal(25), B2 => n169, C1 => A_neg_shifted(25),
                           C2 => n163, ZN => n221);
   U143 : AOI22_X1 port map( A1 => A_neg(25), A2 => n152, B1 => A_signal(25), 
                           B2 => n143, ZN => n222);
   U144 : NAND2_X1 port map( A1 => n278, A2 => n277, ZN => Y(50));
   U145 : AOI222_X1 port map( A1 => A_shifted(50), A2 => n180, B1 => 
                           zeroSignal(50), B2 => n171, C1 => A_neg_shifted(50),
                           C2 => n161, ZN => n277);
   U146 : AOI22_X1 port map( A1 => A_neg(50), A2 => n154, B1 => A_signal(50), 
                           B2 => n145, ZN => n278);
   U147 : NAND2_X1 port map( A1 => n224, A2 => n223, ZN => Y(26));
   U148 : AOI222_X1 port map( A1 => A_shifted(26), A2 => n178, B1 => 
                           zeroSignal(26), B2 => n169, C1 => A_neg_shifted(26),
                           C2 => n163, ZN => n223);
   U149 : AOI22_X1 port map( A1 => A_neg(26), A2 => n152, B1 => A_signal(26), 
                           B2 => n143, ZN => n224);
   U150 : NAND2_X1 port map( A1 => n226, A2 => n225, ZN => Y(27));
   U151 : AOI222_X1 port map( A1 => A_shifted(27), A2 => n178, B1 => 
                           zeroSignal(27), B2 => n169, C1 => A_neg_shifted(27),
                           C2 => n163, ZN => n225);
   U152 : AOI22_X1 port map( A1 => A_neg(27), A2 => n152, B1 => A_signal(27), 
                           B2 => n143, ZN => n226);
   U153 : NAND2_X1 port map( A1 => n282, A2 => n281, ZN => Y(52));
   U154 : AOI222_X1 port map( A1 => A_shifted(52), A2 => n180, B1 => 
                           zeroSignal(52), B2 => n171, C1 => A_neg_shifted(52),
                           C2 => n161, ZN => n281);
   U155 : AOI22_X1 port map( A1 => A_neg(52), A2 => n154, B1 => A_signal(52), 
                           B2 => n145, ZN => n282);
   U156 : NAND2_X1 port map( A1 => n284, A2 => n283, ZN => Y(53));
   U157 : AOI222_X1 port map( A1 => A_shifted(53), A2 => n181, B1 => 
                           zeroSignal(53), B2 => n172, C1 => A_neg_shifted(53),
                           C2 => n161, ZN => n283);
   U158 : AOI22_X1 port map( A1 => A_neg(53), A2 => n155, B1 => A_signal(53), 
                           B2 => n146, ZN => n284);
   U159 : NAND2_X1 port map( A1 => n286, A2 => n285, ZN => Y(54));
   U160 : AOI222_X1 port map( A1 => A_shifted(54), A2 => n181, B1 => 
                           zeroSignal(54), B2 => n172, C1 => A_neg_shifted(54),
                           C2 => n161, ZN => n285);
   U161 : AOI22_X1 port map( A1 => A_neg(54), A2 => n155, B1 => A_signal(54), 
                           B2 => n146, ZN => n286);
   U162 : NAND2_X1 port map( A1 => n288, A2 => n287, ZN => Y(55));
   U163 : AOI22_X1 port map( A1 => A_neg(55), A2 => n155, B1 => A_signal(55), 
                           B2 => n146, ZN => n288);
   U164 : AOI222_X1 port map( A1 => A_shifted(55), A2 => n181, B1 => 
                           zeroSignal(55), B2 => n172, C1 => A_neg_shifted(55),
                           C2 => n161, ZN => n287);
   U165 : NAND2_X1 port map( A1 => n292, A2 => n291, ZN => Y(57));
   U166 : AOI222_X1 port map( A1 => A_shifted(57), A2 => n181, B1 => 
                           zeroSignal(57), B2 => n172, C1 => A_neg_shifted(57),
                           C2 => n160, ZN => n291);
   U167 : AOI22_X1 port map( A1 => A_neg(57), A2 => n155, B1 => A_signal(57), 
                           B2 => n146, ZN => n292);
   U168 : NAND2_X1 port map( A1 => n290, A2 => n289, ZN => Y(56));
   U169 : AOI222_X1 port map( A1 => A_shifted(56), A2 => n181, B1 => 
                           zeroSignal(56), B2 => n172, C1 => A_neg_shifted(56),
                           C2 => n161, ZN => n289);
   U170 : AOI22_X1 port map( A1 => A_neg(56), A2 => n155, B1 => A_signal(56), 
                           B2 => n146, ZN => n290);
   U171 : NAND2_X1 port map( A1 => n294, A2 => n293, ZN => Y(58));
   U172 : AOI222_X1 port map( A1 => A_shifted(58), A2 => n181, B1 => 
                           zeroSignal(58), B2 => n172, C1 => A_neg_shifted(58),
                           C2 => n160, ZN => n293);
   U173 : AOI22_X1 port map( A1 => A_neg(58), A2 => n155, B1 => A_signal(58), 
                           B2 => n146, ZN => n294);
   U174 : NAND2_X1 port map( A1 => n296, A2 => n295, ZN => Y(59));
   U175 : AOI22_X1 port map( A1 => A_neg(59), A2 => n155, B1 => A_signal(59), 
                           B2 => n146, ZN => n296);
   U176 : AOI222_X1 port map( A1 => A_shifted(59), A2 => n181, B1 => 
                           zeroSignal(59), B2 => n172, C1 => A_neg_shifted(59),
                           C2 => n160, ZN => n295);
   U177 : NAND2_X1 port map( A1 => n304, A2 => n303, ZN => Y(62));
   U178 : AOI222_X1 port map( A1 => A_shifted(62), A2 => n181, B1 => 
                           zeroSignal(62), B2 => n172, C1 => A_neg_shifted(62),
                           C2 => n160, ZN => n303);
   U179 : NAND2_X1 port map( A1 => n302, A2 => n301, ZN => Y(61));
   U180 : AOI222_X1 port map( A1 => A_shifted(61), A2 => n181, B1 => 
                           zeroSignal(61), B2 => n172, C1 => A_neg_shifted(61),
                           C2 => n160, ZN => n301);
   U181 : AOI22_X1 port map( A1 => A_neg(61), A2 => n155, B1 => A_signal(61), 
                           B2 => n146, ZN => n302);
   U182 : NAND2_X1 port map( A1 => n306, A2 => n305, ZN => Y(63));
   U183 : AOI22_X1 port map( A1 => A_neg(63), A2 => n155, B1 => A_signal(63), 
                           B2 => n146, ZN => n306);
   U184 : NAND2_X1 port map( A1 => n300, A2 => n299, ZN => Y(60));
   U185 : AOI22_X1 port map( A1 => A_neg(60), A2 => n155, B1 => A_signal(60), 
                           B2 => n146, ZN => n300);
   U186 : AOI222_X1 port map( A1 => A_shifted(60), A2 => n181, B1 => 
                           zeroSignal(60), B2 => n172, C1 => A_neg_shifted(60),
                           C2 => n160, ZN => n299);
   U187 : NAND2_X1 port map( A1 => n188, A2 => n187, ZN => Y(0));
   U188 : AOI22_X1 port map( A1 => A_neg(0), A2 => n151, B1 => A_signal(0), B2 
                           => n142, ZN => n188);
   U189 : AOI222_X1 port map( A1 => A_shifted(0), A2 => n177, B1 => 
                           zeroSignal(0), B2 => n168, C1 => A_neg_shifted(0), 
                           C2 => n165, ZN => n187);
   U190 : NAND2_X1 port map( A1 => n210, A2 => n209, ZN => Y(1));
   U191 : AOI22_X1 port map( A1 => A_neg(1), A2 => n151, B1 => A_signal(1), B2 
                           => n142, ZN => n210);
   U192 : AOI222_X1 port map( A1 => A_shifted(1), A2 => n177, B1 => 
                           zeroSignal(1), B2 => n168, C1 => A_neg_shifted(1), 
                           C2 => n164, ZN => n209);
   U193 : NAND2_X1 port map( A1 => n232, A2 => n231, ZN => Y(2));
   U194 : AOI22_X1 port map( A1 => A_neg(2), A2 => n152, B1 => A_signal(2), B2 
                           => n143, ZN => n232);
   U195 : AOI222_X1 port map( A1 => A_shifted(2), A2 => n178, B1 => 
                           zeroSignal(2), B2 => n169, C1 => A_neg_shifted(2), 
                           C2 => n163, ZN => n231);
   U196 : NAND2_X1 port map( A1 => n254, A2 => n253, ZN => Y(3));
   U197 : AOI22_X1 port map( A1 => A_neg(3), A2 => n153, B1 => A_signal(3), B2 
                           => n144, ZN => n254);
   U198 : AOI222_X1 port map( A1 => A_shifted(3), A2 => n179, B1 => 
                           zeroSignal(3), B2 => n170, C1 => A_neg_shifted(3), 
                           C2 => n162, ZN => n253);
   U199 : NAND2_X1 port map( A1 => n276, A2 => n275, ZN => Y(4));
   U200 : AOI22_X1 port map( A1 => A_neg(4), A2 => n154, B1 => A_signal(4), B2 
                           => n145, ZN => n276);
   U201 : AOI222_X1 port map( A1 => A_shifted(4), A2 => n180, B1 => 
                           zeroSignal(4), B2 => n171, C1 => A_neg_shifted(4), 
                           C2 => n161, ZN => n275);
   U202 : NAND2_X1 port map( A1 => n298, A2 => n297, ZN => Y(5));
   U203 : AOI22_X1 port map( A1 => A_neg(5), A2 => n155, B1 => A_signal(5), B2 
                           => n146, ZN => n298);
   U204 : AOI222_X1 port map( A1 => A_shifted(5), A2 => n181, B1 => 
                           zeroSignal(5), B2 => n172, C1 => A_neg_shifted(5), 
                           C2 => n160, ZN => n297);
   U205 : NAND2_X1 port map( A1 => n308, A2 => n307, ZN => Y(6));
   U206 : AOI22_X1 port map( A1 => A_neg(6), A2 => n156, B1 => A_signal(6), B2 
                           => n147, ZN => n308);
   U207 : AOI222_X1 port map( A1 => A_shifted(6), A2 => n182, B1 => 
                           zeroSignal(6), B2 => n173, C1 => A_neg_shifted(6), 
                           C2 => n160, ZN => n307);
   U208 : NAND2_X1 port map( A1 => n310, A2 => n309, ZN => Y(7));
   U209 : AOI22_X1 port map( A1 => A_neg(7), A2 => n156, B1 => A_signal(7), B2 
                           => n147, ZN => n310);
   U210 : AOI222_X1 port map( A1 => A_shifted(7), A2 => n182, B1 => 
                           zeroSignal(7), B2 => n173, C1 => A_neg_shifted(7), 
                           C2 => n160, ZN => n309);
   U211 : NAND2_X1 port map( A1 => n312, A2 => n311, ZN => Y(8));
   U212 : AOI22_X1 port map( A1 => A_neg(8), A2 => n156, B1 => A_signal(8), B2 
                           => n147, ZN => n312);
   U213 : AOI222_X1 port map( A1 => A_shifted(8), A2 => n182, B1 => 
                           zeroSignal(8), B2 => n173, C1 => A_neg_shifted(8), 
                           C2 => n160, ZN => n311);
   U214 : NAND2_X1 port map( A1 => n318, A2 => n317, ZN => Y(9));
   U215 : AOI22_X1 port map( A1 => A_neg(9), A2 => n156, B1 => A_signal(9), B2 
                           => n147, ZN => n318);
   U216 : AOI222_X1 port map( A1 => A_shifted(9), A2 => n182, B1 => 
                           zeroSignal(9), B2 => n173, C1 => A_neg_shifted(9), 
                           C2 => n160, ZN => n317);
   U217 : NAND2_X1 port map( A1 => n190, A2 => n189, ZN => Y(10));
   U218 : AOI22_X1 port map( A1 => A_neg(10), A2 => n151, B1 => A_signal(10), 
                           B2 => n142, ZN => n190);
   U219 : AOI222_X1 port map( A1 => A_shifted(10), A2 => n177, B1 => 
                           zeroSignal(10), B2 => n168, C1 => A_neg_shifted(10),
                           C2 => n165, ZN => n189);
   U220 : NAND2_X1 port map( A1 => n192, A2 => n191, ZN => Y(11));
   U221 : AOI22_X1 port map( A1 => A_neg(11), A2 => n151, B1 => A_signal(11), 
                           B2 => n142, ZN => n192);
   U222 : AOI222_X1 port map( A1 => A_shifted(11), A2 => n177, B1 => 
                           zeroSignal(11), B2 => n168, C1 => A_neg_shifted(11),
                           C2 => n165, ZN => n191);
   U223 : NAND2_X1 port map( A1 => n194, A2 => n193, ZN => Y(12));
   U224 : AOI22_X1 port map( A1 => A_neg(12), A2 => n151, B1 => A_signal(12), 
                           B2 => n142, ZN => n194);
   U225 : AOI222_X1 port map( A1 => A_shifted(12), A2 => n177, B1 => 
                           zeroSignal(12), B2 => n168, C1 => A_neg_shifted(12),
                           C2 => n165, ZN => n193);
   U226 : NAND2_X1 port map( A1 => n196, A2 => n195, ZN => Y(13));
   U227 : AOI22_X1 port map( A1 => A_neg(13), A2 => n151, B1 => A_signal(13), 
                           B2 => n142, ZN => n196);
   U228 : AOI222_X1 port map( A1 => A_shifted(13), A2 => n177, B1 => 
                           zeroSignal(13), B2 => n168, C1 => A_neg_shifted(13),
                           C2 => n164, ZN => n195);
   U229 : NAND2_X1 port map( A1 => n198, A2 => n197, ZN => Y(14));
   U230 : AOI22_X1 port map( A1 => A_neg(14), A2 => n151, B1 => A_signal(14), 
                           B2 => n142, ZN => n198);
   U231 : AOI222_X1 port map( A1 => A_shifted(14), A2 => n177, B1 => 
                           zeroSignal(14), B2 => n168, C1 => A_neg_shifted(14),
                           C2 => n164, ZN => n197);
   U232 : NAND2_X1 port map( A1 => n200, A2 => n199, ZN => Y(15));
   U233 : AOI22_X1 port map( A1 => A_neg(15), A2 => n151, B1 => A_signal(15), 
                           B2 => n142, ZN => n200);
   U234 : AOI222_X1 port map( A1 => A_shifted(15), A2 => n177, B1 => 
                           zeroSignal(15), B2 => n168, C1 => A_neg_shifted(15),
                           C2 => n164, ZN => n199);
   U235 : NAND2_X1 port map( A1 => n202, A2 => n201, ZN => Y(16));
   U236 : AOI22_X1 port map( A1 => A_neg(16), A2 => n151, B1 => A_signal(16), 
                           B2 => n142, ZN => n202);
   U237 : AOI222_X1 port map( A1 => A_shifted(16), A2 => n177, B1 => 
                           zeroSignal(16), B2 => n168, C1 => A_neg_shifted(16),
                           C2 => n164, ZN => n201);
   U238 : NAND2_X1 port map( A1 => n204, A2 => n203, ZN => Y(17));
   U239 : AOI22_X1 port map( A1 => A_neg(17), A2 => n151, B1 => A_signal(17), 
                           B2 => n142, ZN => n204);
   U240 : AOI222_X1 port map( A1 => A_shifted(17), A2 => n177, B1 => 
                           zeroSignal(17), B2 => n168, C1 => A_neg_shifted(17),
                           C2 => n164, ZN => n203);
   U241 : AOI222_X1 port map( A1 => A_shifted(63), A2 => n181, B1 => 
                           zeroSignal(63), B2 => n172, C1 => A_neg_shifted(63),
                           C2 => n160, ZN => n305);
   U242 : AOI22_X1 port map( A1 => A_neg(62), A2 => n155, B1 => A_signal(62), 
                           B2 => n146, ZN => n304);
   U243 : AOI222_X1 port map( A1 => A_shifted(19), A2 => n177, B1 => 
                           zeroSignal(19), B2 => n168, C1 => A_neg_shifted(19),
                           C2 => n164, ZN => n207);
   U244 : AOI22_X1 port map( A1 => A_neg(18), A2 => n151, B1 => A_signal(18), 
                           B2 => n142, ZN => n206);

end SYN_BEHAVIORAL_2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity MUX51_MuxNbit64_22 is

   port( zeroSignal, A_signal, A_neg, A_shifted, A_neg_shifted : in 
         std_logic_vector (63 downto 0);  Sel : in std_logic_vector (2 downto 
         0);  Y : out std_logic_vector (63 downto 0));

end MUX51_MuxNbit64_22;

architecture SYN_BEHAVIORAL_2 of MUX51_MuxNbit64_22 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, 
      n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, 
      n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, 
      n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, 
      n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, 
      n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, 
      n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, 
      n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, 
      n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, 
      n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, 
      n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, 
      n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, 
      n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, 
      n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, 
      n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, 
      n320 : std_logic;

begin
   
   U1 : AND3_X1 port map( A1 => n319, A2 => n320, A3 => Sel(2), ZN => n141);
   U2 : BUF_X1 port map( A => n141, Z => n166);
   U3 : BUF_X1 port map( A => n185, Z => n184);
   U4 : BUF_X1 port map( A => n159, Z => n158);
   U5 : BUF_X1 port map( A => n150, Z => n149);
   U6 : BUF_X1 port map( A => n141, Z => n167);
   U7 : BUF_X1 port map( A => n185, Z => n183);
   U8 : BUF_X1 port map( A => n159, Z => n157);
   U9 : BUF_X1 port map( A => n150, Z => n148);
   U10 : BUF_X1 port map( A => n176, Z => n175);
   U11 : BUF_X1 port map( A => n176, Z => n174);
   U12 : BUF_X1 port map( A => n158, Z => n152);
   U13 : BUF_X1 port map( A => n184, Z => n178);
   U14 : BUF_X1 port map( A => n149, Z => n143);
   U15 : BUF_X1 port map( A => n166, Z => n164);
   U16 : BUF_X1 port map( A => n166, Z => n163);
   U17 : BUF_X1 port map( A => n184, Z => n179);
   U18 : BUF_X1 port map( A => n158, Z => n153);
   U19 : BUF_X1 port map( A => n149, Z => n144);
   U20 : BUF_X1 port map( A => n167, Z => n162);
   U21 : BUF_X1 port map( A => n183, Z => n180);
   U22 : BUF_X1 port map( A => n157, Z => n154);
   U23 : BUF_X1 port map( A => n148, Z => n145);
   U24 : BUF_X1 port map( A => n167, Z => n161);
   U25 : BUF_X1 port map( A => n183, Z => n181);
   U26 : BUF_X1 port map( A => n157, Z => n155);
   U27 : BUF_X1 port map( A => n148, Z => n146);
   U28 : BUF_X1 port map( A => n167, Z => n160);
   U29 : BUF_X1 port map( A => n158, Z => n151);
   U30 : BUF_X1 port map( A => n149, Z => n142);
   U31 : BUF_X1 port map( A => n175, Z => n168);
   U32 : BUF_X1 port map( A => n175, Z => n170);
   U33 : BUF_X1 port map( A => n174, Z => n171);
   U34 : BUF_X1 port map( A => n174, Z => n172);
   U35 : BUF_X1 port map( A => n175, Z => n169);
   U36 : BUF_X1 port map( A => n184, Z => n177);
   U37 : BUF_X1 port map( A => n166, Z => n165);
   U38 : BUF_X1 port map( A => n157, Z => n156);
   U39 : BUF_X1 port map( A => n148, Z => n147);
   U40 : BUF_X1 port map( A => n174, Z => n173);
   U41 : BUF_X1 port map( A => n183, Z => n182);
   U42 : INV_X1 port map( A => Sel(1), ZN => n320);
   U43 : BUF_X1 port map( A => n314, Z => n159);
   U44 : NOR3_X1 port map( A1 => Sel(0), A2 => Sel(2), A3 => n320, ZN => n314);
   U45 : BUF_X1 port map( A => n316, Z => n185);
   U46 : NOR3_X1 port map( A1 => n319, A2 => Sel(2), A3 => n320, ZN => n316);
   U47 : INV_X1 port map( A => Sel(0), ZN => n319);
   U48 : BUF_X1 port map( A => n313, Z => n150);
   U49 : NOR3_X1 port map( A1 => Sel(1), A2 => Sel(2), A3 => n319, ZN => n313);
   U50 : BUF_X1 port map( A => n315, Z => n176);
   U51 : NOR2_X1 port map( A1 => n165, A2 => n186, ZN => n315);
   U52 : AOI21_X1 port map( B1 => n319, B2 => n320, A => Sel(2), ZN => n186);
   U53 : NAND2_X1 port map( A1 => n214, A2 => n213, ZN => Y(21));
   U54 : AOI22_X1 port map( A1 => A_neg(21), A2 => n152, B1 => A_signal(21), B2
                           => n143, ZN => n214);
   U55 : NAND2_X1 port map( A1 => n212, A2 => n211, ZN => Y(20));
   U56 : AOI222_X1 port map( A1 => A_shifted(20), A2 => n178, B1 => 
                           zeroSignal(20), B2 => n169, C1 => A_neg_shifted(20),
                           C2 => n164, ZN => n211);
   U57 : NAND2_X1 port map( A1 => n216, A2 => n215, ZN => Y(22));
   U58 : AOI22_X1 port map( A1 => A_neg(22), A2 => n152, B1 => A_signal(22), B2
                           => n143, ZN => n216);
   U59 : AOI222_X1 port map( A1 => A_shifted(22), A2 => n178, B1 => 
                           zeroSignal(22), B2 => n169, C1 => A_neg_shifted(22),
                           C2 => n164, ZN => n215);
   U60 : NAND2_X1 port map( A1 => n218, A2 => n217, ZN => Y(23));
   U61 : AOI22_X1 port map( A1 => A_neg(23), A2 => n152, B1 => A_signal(23), B2
                           => n143, ZN => n218);
   U62 : AOI222_X1 port map( A1 => A_shifted(23), A2 => n178, B1 => 
                           zeroSignal(23), B2 => n169, C1 => A_neg_shifted(23),
                           C2 => n164, ZN => n217);
   U63 : NAND2_X1 port map( A1 => n236, A2 => n235, ZN => Y(31));
   U64 : AOI222_X1 port map( A1 => A_shifted(31), A2 => n179, B1 => 
                           zeroSignal(31), B2 => n170, C1 => A_neg_shifted(31),
                           C2 => n163, ZN => n235);
   U65 : AOI22_X1 port map( A1 => A_neg(31), A2 => n153, B1 => A_signal(31), B2
                           => n144, ZN => n236);
   U66 : NAND2_X1 port map( A1 => n220, A2 => n219, ZN => Y(24));
   U67 : AOI22_X1 port map( A1 => A_neg(24), A2 => n152, B1 => A_signal(24), B2
                           => n143, ZN => n220);
   U68 : AOI222_X1 port map( A1 => A_shifted(24), A2 => n178, B1 => 
                           zeroSignal(24), B2 => n169, C1 => A_neg_shifted(24),
                           C2 => n163, ZN => n219);
   U69 : NAND2_X1 port map( A1 => n234, A2 => n233, ZN => Y(30));
   U70 : AOI222_X1 port map( A1 => A_shifted(30), A2 => n178, B1 => 
                           zeroSignal(30), B2 => n169, C1 => A_neg_shifted(30),
                           C2 => n163, ZN => n233);
   U71 : AOI22_X1 port map( A1 => A_neg(30), A2 => n152, B1 => A_signal(30), B2
                           => n143, ZN => n234);
   U72 : NAND2_X1 port map( A1 => n244, A2 => n243, ZN => Y(35));
   U73 : AOI222_X1 port map( A1 => A_shifted(35), A2 => n179, B1 => 
                           zeroSignal(35), B2 => n170, C1 => A_neg_shifted(35),
                           C2 => n162, ZN => n243);
   U74 : AOI22_X1 port map( A1 => A_neg(35), A2 => n153, B1 => A_signal(35), B2
                           => n144, ZN => n244);
   U75 : NAND2_X1 port map( A1 => n238, A2 => n237, ZN => Y(32));
   U76 : AOI222_X1 port map( A1 => A_shifted(32), A2 => n179, B1 => 
                           zeroSignal(32), B2 => n170, C1 => A_neg_shifted(32),
                           C2 => n163, ZN => n237);
   U77 : AOI22_X1 port map( A1 => A_neg(32), A2 => n153, B1 => A_signal(32), B2
                           => n144, ZN => n238);
   U78 : NAND2_X1 port map( A1 => n240, A2 => n239, ZN => Y(33));
   U79 : AOI222_X1 port map( A1 => A_shifted(33), A2 => n179, B1 => 
                           zeroSignal(33), B2 => n170, C1 => A_neg_shifted(33),
                           C2 => n163, ZN => n239);
   U80 : AOI22_X1 port map( A1 => A_neg(33), A2 => n153, B1 => A_signal(33), B2
                           => n144, ZN => n240);
   U81 : NAND2_X1 port map( A1 => n246, A2 => n245, ZN => Y(36));
   U82 : AOI222_X1 port map( A1 => A_shifted(36), A2 => n179, B1 => 
                           zeroSignal(36), B2 => n170, C1 => A_neg_shifted(36),
                           C2 => n162, ZN => n245);
   U83 : AOI22_X1 port map( A1 => A_neg(36), A2 => n153, B1 => A_signal(36), B2
                           => n144, ZN => n246);
   U84 : NAND2_X1 port map( A1 => n248, A2 => n247, ZN => Y(37));
   U85 : AOI222_X1 port map( A1 => A_shifted(37), A2 => n179, B1 => 
                           zeroSignal(37), B2 => n170, C1 => A_neg_shifted(37),
                           C2 => n162, ZN => n247);
   U86 : AOI22_X1 port map( A1 => A_neg(37), A2 => n153, B1 => A_signal(37), B2
                           => n144, ZN => n248);
   U87 : NAND2_X1 port map( A1 => n252, A2 => n251, ZN => Y(39));
   U88 : AOI222_X1 port map( A1 => A_shifted(39), A2 => n179, B1 => 
                           zeroSignal(39), B2 => n170, C1 => A_neg_shifted(39),
                           C2 => n162, ZN => n251);
   U89 : AOI22_X1 port map( A1 => A_neg(39), A2 => n153, B1 => A_signal(39), B2
                           => n144, ZN => n252);
   U90 : NAND2_X1 port map( A1 => n256, A2 => n255, ZN => Y(40));
   U91 : AOI222_X1 port map( A1 => A_shifted(40), A2 => n179, B1 => 
                           zeroSignal(40), B2 => n170, C1 => A_neg_shifted(40),
                           C2 => n162, ZN => n255);
   U92 : AOI22_X1 port map( A1 => A_neg(40), A2 => n153, B1 => A_signal(40), B2
                           => n144, ZN => n256);
   U93 : NAND2_X1 port map( A1 => n258, A2 => n257, ZN => Y(41));
   U94 : AOI222_X1 port map( A1 => A_shifted(41), A2 => n179, B1 => 
                           zeroSignal(41), B2 => n170, C1 => A_neg_shifted(41),
                           C2 => n162, ZN => n257);
   U95 : AOI22_X1 port map( A1 => A_neg(41), A2 => n153, B1 => A_signal(41), B2
                           => n144, ZN => n258);
   U96 : NAND2_X1 port map( A1 => n242, A2 => n241, ZN => Y(34));
   U97 : AOI22_X1 port map( A1 => A_neg(34), A2 => n153, B1 => A_signal(34), B2
                           => n144, ZN => n242);
   U98 : AOI222_X1 port map( A1 => A_shifted(34), A2 => n179, B1 => 
                           zeroSignal(34), B2 => n170, C1 => A_neg_shifted(34),
                           C2 => n163, ZN => n241);
   U99 : NAND2_X1 port map( A1 => n222, A2 => n221, ZN => Y(25));
   U100 : AOI22_X1 port map( A1 => A_neg(25), A2 => n152, B1 => A_signal(25), 
                           B2 => n143, ZN => n222);
   U101 : AOI222_X1 port map( A1 => A_shifted(25), A2 => n178, B1 => 
                           zeroSignal(25), B2 => n169, C1 => A_neg_shifted(25),
                           C2 => n163, ZN => n221);
   U102 : NAND2_X1 port map( A1 => n260, A2 => n259, ZN => Y(42));
   U103 : AOI222_X1 port map( A1 => A_shifted(42), A2 => n180, B1 => 
                           zeroSignal(42), B2 => n171, C1 => A_neg_shifted(42),
                           C2 => n162, ZN => n259);
   U104 : AOI22_X1 port map( A1 => A_neg(42), A2 => n154, B1 => A_signal(42), 
                           B2 => n145, ZN => n260);
   U105 : NAND2_X1 port map( A1 => n262, A2 => n261, ZN => Y(43));
   U106 : AOI222_X1 port map( A1 => A_shifted(43), A2 => n180, B1 => 
                           zeroSignal(43), B2 => n171, C1 => A_neg_shifted(43),
                           C2 => n162, ZN => n261);
   U107 : AOI22_X1 port map( A1 => A_neg(43), A2 => n154, B1 => A_signal(43), 
                           B2 => n145, ZN => n262);
   U108 : NAND2_X1 port map( A1 => n250, A2 => n249, ZN => Y(38));
   U109 : AOI22_X1 port map( A1 => A_neg(38), A2 => n153, B1 => A_signal(38), 
                           B2 => n144, ZN => n250);
   U110 : AOI222_X1 port map( A1 => A_shifted(38), A2 => n179, B1 => 
                           zeroSignal(38), B2 => n170, C1 => A_neg_shifted(38),
                           C2 => n162, ZN => n249);
   U111 : NAND2_X1 port map( A1 => n266, A2 => n265, ZN => Y(45));
   U112 : AOI222_X1 port map( A1 => A_shifted(45), A2 => n180, B1 => 
                           zeroSignal(45), B2 => n171, C1 => A_neg_shifted(45),
                           C2 => n162, ZN => n265);
   U113 : AOI22_X1 port map( A1 => A_neg(45), A2 => n154, B1 => A_signal(45), 
                           B2 => n145, ZN => n266);
   U114 : NAND2_X1 port map( A1 => n268, A2 => n267, ZN => Y(46));
   U115 : AOI222_X1 port map( A1 => A_shifted(46), A2 => n180, B1 => 
                           zeroSignal(46), B2 => n171, C1 => A_neg_shifted(46),
                           C2 => n161, ZN => n267);
   U116 : AOI22_X1 port map( A1 => A_neg(46), A2 => n154, B1 => A_signal(46), 
                           B2 => n145, ZN => n268);
   U117 : NAND2_X1 port map( A1 => n270, A2 => n269, ZN => Y(47));
   U118 : AOI222_X1 port map( A1 => A_shifted(47), A2 => n180, B1 => 
                           zeroSignal(47), B2 => n171, C1 => A_neg_shifted(47),
                           C2 => n161, ZN => n269);
   U119 : AOI22_X1 port map( A1 => A_neg(47), A2 => n154, B1 => A_signal(47), 
                           B2 => n145, ZN => n270);
   U120 : NAND2_X1 port map( A1 => n284, A2 => n283, ZN => Y(53));
   U121 : AOI222_X1 port map( A1 => A_shifted(53), A2 => n181, B1 => 
                           zeroSignal(53), B2 => n172, C1 => A_neg_shifted(53),
                           C2 => n161, ZN => n283);
   U122 : AOI22_X1 port map( A1 => A_neg(53), A2 => n155, B1 => A_signal(53), 
                           B2 => n146, ZN => n284);
   U123 : NAND2_X1 port map( A1 => n264, A2 => n263, ZN => Y(44));
   U124 : AOI22_X1 port map( A1 => A_neg(44), A2 => n154, B1 => A_signal(44), 
                           B2 => n145, ZN => n264);
   U125 : AOI222_X1 port map( A1 => A_shifted(44), A2 => n180, B1 => 
                           zeroSignal(44), B2 => n171, C1 => A_neg_shifted(44),
                           C2 => n162, ZN => n263);
   U126 : NAND2_X1 port map( A1 => n272, A2 => n271, ZN => Y(48));
   U127 : AOI222_X1 port map( A1 => A_shifted(48), A2 => n180, B1 => 
                           zeroSignal(48), B2 => n171, C1 => A_neg_shifted(48),
                           C2 => n161, ZN => n271);
   U128 : AOI22_X1 port map( A1 => A_neg(48), A2 => n154, B1 => A_signal(48), 
                           B2 => n145, ZN => n272);
   U129 : NAND2_X1 port map( A1 => n274, A2 => n273, ZN => Y(49));
   U130 : AOI222_X1 port map( A1 => A_shifted(49), A2 => n180, B1 => 
                           zeroSignal(49), B2 => n171, C1 => A_neg_shifted(49),
                           C2 => n161, ZN => n273);
   U131 : AOI22_X1 port map( A1 => A_neg(49), A2 => n154, B1 => A_signal(49), 
                           B2 => n145, ZN => n274);
   U132 : NAND2_X1 port map( A1 => n280, A2 => n279, ZN => Y(51));
   U133 : AOI222_X1 port map( A1 => A_shifted(51), A2 => n180, B1 => 
                           zeroSignal(51), B2 => n171, C1 => A_neg_shifted(51),
                           C2 => n161, ZN => n279);
   U134 : AOI22_X1 port map( A1 => A_neg(51), A2 => n154, B1 => A_signal(51), 
                           B2 => n145, ZN => n280);
   U135 : NAND2_X1 port map( A1 => n282, A2 => n281, ZN => Y(52));
   U136 : AOI222_X1 port map( A1 => A_shifted(52), A2 => n180, B1 => 
                           zeroSignal(52), B2 => n171, C1 => A_neg_shifted(52),
                           C2 => n161, ZN => n281);
   U137 : AOI22_X1 port map( A1 => A_neg(52), A2 => n154, B1 => A_signal(52), 
                           B2 => n145, ZN => n282);
   U138 : NAND2_X1 port map( A1 => n278, A2 => n277, ZN => Y(50));
   U139 : AOI222_X1 port map( A1 => A_shifted(50), A2 => n180, B1 => 
                           zeroSignal(50), B2 => n171, C1 => A_neg_shifted(50),
                           C2 => n161, ZN => n277);
   U140 : AOI22_X1 port map( A1 => A_neg(50), A2 => n154, B1 => A_signal(50), 
                           B2 => n145, ZN => n278);
   U141 : NAND2_X1 port map( A1 => n224, A2 => n223, ZN => Y(26));
   U142 : AOI222_X1 port map( A1 => A_shifted(26), A2 => n178, B1 => 
                           zeroSignal(26), B2 => n169, C1 => A_neg_shifted(26),
                           C2 => n163, ZN => n223);
   U143 : AOI22_X1 port map( A1 => A_neg(26), A2 => n152, B1 => A_signal(26), 
                           B2 => n143, ZN => n224);
   U144 : NAND2_X1 port map( A1 => n226, A2 => n225, ZN => Y(27));
   U145 : AOI222_X1 port map( A1 => A_shifted(27), A2 => n178, B1 => 
                           zeroSignal(27), B2 => n169, C1 => A_neg_shifted(27),
                           C2 => n163, ZN => n225);
   U146 : AOI22_X1 port map( A1 => A_neg(27), A2 => n152, B1 => A_signal(27), 
                           B2 => n143, ZN => n226);
   U147 : NAND2_X1 port map( A1 => n228, A2 => n227, ZN => Y(28));
   U148 : AOI222_X1 port map( A1 => A_shifted(28), A2 => n178, B1 => 
                           zeroSignal(28), B2 => n169, C1 => A_neg_shifted(28),
                           C2 => n163, ZN => n227);
   U149 : AOI22_X1 port map( A1 => A_neg(28), A2 => n152, B1 => A_signal(28), 
                           B2 => n143, ZN => n228);
   U150 : NAND2_X1 port map( A1 => n230, A2 => n229, ZN => Y(29));
   U151 : AOI222_X1 port map( A1 => A_shifted(29), A2 => n178, B1 => 
                           zeroSignal(29), B2 => n169, C1 => A_neg_shifted(29),
                           C2 => n163, ZN => n229);
   U152 : AOI22_X1 port map( A1 => A_neg(29), A2 => n152, B1 => A_signal(29), 
                           B2 => n143, ZN => n230);
   U153 : NAND2_X1 port map( A1 => n286, A2 => n285, ZN => Y(54));
   U154 : AOI22_X1 port map( A1 => A_neg(54), A2 => n155, B1 => A_signal(54), 
                           B2 => n146, ZN => n286);
   U155 : AOI222_X1 port map( A1 => A_shifted(54), A2 => n181, B1 => 
                           zeroSignal(54), B2 => n172, C1 => A_neg_shifted(54),
                           C2 => n161, ZN => n285);
   U156 : NAND2_X1 port map( A1 => n288, A2 => n287, ZN => Y(55));
   U157 : AOI222_X1 port map( A1 => A_shifted(55), A2 => n181, B1 => 
                           zeroSignal(55), B2 => n172, C1 => A_neg_shifted(55),
                           C2 => n161, ZN => n287);
   U158 : AOI22_X1 port map( A1 => A_neg(55), A2 => n155, B1 => A_signal(55), 
                           B2 => n146, ZN => n288);
   U159 : NAND2_X1 port map( A1 => n290, A2 => n289, ZN => Y(56));
   U160 : AOI222_X1 port map( A1 => A_shifted(56), A2 => n181, B1 => 
                           zeroSignal(56), B2 => n172, C1 => A_neg_shifted(56),
                           C2 => n161, ZN => n289);
   U161 : AOI22_X1 port map( A1 => A_neg(56), A2 => n155, B1 => A_signal(56), 
                           B2 => n146, ZN => n290);
   U162 : NAND2_X1 port map( A1 => n292, A2 => n291, ZN => Y(57));
   U163 : AOI22_X1 port map( A1 => A_neg(57), A2 => n155, B1 => A_signal(57), 
                           B2 => n146, ZN => n292);
   U164 : AOI222_X1 port map( A1 => A_shifted(57), A2 => n181, B1 => 
                           zeroSignal(57), B2 => n172, C1 => A_neg_shifted(57),
                           C2 => n160, ZN => n291);
   U165 : NAND2_X1 port map( A1 => n296, A2 => n295, ZN => Y(59));
   U166 : AOI222_X1 port map( A1 => A_shifted(59), A2 => n181, B1 => 
                           zeroSignal(59), B2 => n172, C1 => A_neg_shifted(59),
                           C2 => n160, ZN => n295);
   U167 : AOI22_X1 port map( A1 => A_neg(59), A2 => n155, B1 => A_signal(59), 
                           B2 => n146, ZN => n296);
   U168 : NAND2_X1 port map( A1 => n300, A2 => n299, ZN => Y(60));
   U169 : AOI222_X1 port map( A1 => A_shifted(60), A2 => n181, B1 => 
                           zeroSignal(60), B2 => n172, C1 => A_neg_shifted(60),
                           C2 => n160, ZN => n299);
   U170 : AOI22_X1 port map( A1 => A_neg(60), A2 => n155, B1 => A_signal(60), 
                           B2 => n146, ZN => n300);
   U171 : NAND2_X1 port map( A1 => n294, A2 => n293, ZN => Y(58));
   U172 : AOI222_X1 port map( A1 => A_shifted(58), A2 => n181, B1 => 
                           zeroSignal(58), B2 => n172, C1 => A_neg_shifted(58),
                           C2 => n160, ZN => n293);
   U173 : AOI22_X1 port map( A1 => A_neg(58), A2 => n155, B1 => A_signal(58), 
                           B2 => n146, ZN => n294);
   U174 : NAND2_X1 port map( A1 => n302, A2 => n301, ZN => Y(61));
   U175 : AOI22_X1 port map( A1 => A_neg(61), A2 => n155, B1 => A_signal(61), 
                           B2 => n146, ZN => n302);
   U176 : AOI222_X1 port map( A1 => A_shifted(61), A2 => n181, B1 => 
                           zeroSignal(61), B2 => n172, C1 => A_neg_shifted(61),
                           C2 => n160, ZN => n301);
   U177 : NAND2_X1 port map( A1 => n306, A2 => n305, ZN => Y(63));
   U178 : AOI222_X1 port map( A1 => A_shifted(63), A2 => n181, B1 => 
                           zeroSignal(63), B2 => n172, C1 => A_neg_shifted(63),
                           C2 => n160, ZN => n305);
   U179 : AOI22_X1 port map( A1 => A_neg(63), A2 => n155, B1 => A_signal(63), 
                           B2 => n146, ZN => n306);
   U180 : NAND2_X1 port map( A1 => n304, A2 => n303, ZN => Y(62));
   U181 : AOI22_X1 port map( A1 => A_neg(62), A2 => n155, B1 => A_signal(62), 
                           B2 => n146, ZN => n304);
   U182 : AOI222_X1 port map( A1 => A_shifted(62), A2 => n181, B1 => 
                           zeroSignal(62), B2 => n172, C1 => A_neg_shifted(62),
                           C2 => n160, ZN => n303);
   U183 : NAND2_X1 port map( A1 => n188, A2 => n187, ZN => Y(0));
   U184 : AOI22_X1 port map( A1 => A_neg(0), A2 => n151, B1 => A_signal(0), B2 
                           => n142, ZN => n188);
   U185 : AOI222_X1 port map( A1 => A_shifted(0), A2 => n177, B1 => 
                           zeroSignal(0), B2 => n168, C1 => A_neg_shifted(0), 
                           C2 => n165, ZN => n187);
   U186 : NAND2_X1 port map( A1 => n210, A2 => n209, ZN => Y(1));
   U187 : AOI22_X1 port map( A1 => A_neg(1), A2 => n151, B1 => A_signal(1), B2 
                           => n142, ZN => n210);
   U188 : AOI222_X1 port map( A1 => A_shifted(1), A2 => n177, B1 => 
                           zeroSignal(1), B2 => n168, C1 => A_neg_shifted(1), 
                           C2 => n164, ZN => n209);
   U189 : NAND2_X1 port map( A1 => n232, A2 => n231, ZN => Y(2));
   U190 : AOI22_X1 port map( A1 => A_neg(2), A2 => n152, B1 => A_signal(2), B2 
                           => n143, ZN => n232);
   U191 : AOI222_X1 port map( A1 => A_shifted(2), A2 => n178, B1 => 
                           zeroSignal(2), B2 => n169, C1 => A_neg_shifted(2), 
                           C2 => n163, ZN => n231);
   U192 : NAND2_X1 port map( A1 => n254, A2 => n253, ZN => Y(3));
   U193 : AOI22_X1 port map( A1 => A_neg(3), A2 => n153, B1 => A_signal(3), B2 
                           => n144, ZN => n254);
   U194 : AOI222_X1 port map( A1 => A_shifted(3), A2 => n179, B1 => 
                           zeroSignal(3), B2 => n170, C1 => A_neg_shifted(3), 
                           C2 => n162, ZN => n253);
   U195 : NAND2_X1 port map( A1 => n276, A2 => n275, ZN => Y(4));
   U196 : AOI22_X1 port map( A1 => A_neg(4), A2 => n154, B1 => A_signal(4), B2 
                           => n145, ZN => n276);
   U197 : AOI222_X1 port map( A1 => A_shifted(4), A2 => n180, B1 => 
                           zeroSignal(4), B2 => n171, C1 => A_neg_shifted(4), 
                           C2 => n161, ZN => n275);
   U198 : NAND2_X1 port map( A1 => n298, A2 => n297, ZN => Y(5));
   U199 : AOI22_X1 port map( A1 => A_neg(5), A2 => n155, B1 => A_signal(5), B2 
                           => n146, ZN => n298);
   U200 : AOI222_X1 port map( A1 => A_shifted(5), A2 => n181, B1 => 
                           zeroSignal(5), B2 => n172, C1 => A_neg_shifted(5), 
                           C2 => n160, ZN => n297);
   U201 : NAND2_X1 port map( A1 => n308, A2 => n307, ZN => Y(6));
   U202 : AOI22_X1 port map( A1 => A_neg(6), A2 => n156, B1 => A_signal(6), B2 
                           => n147, ZN => n308);
   U203 : AOI222_X1 port map( A1 => A_shifted(6), A2 => n182, B1 => 
                           zeroSignal(6), B2 => n173, C1 => A_neg_shifted(6), 
                           C2 => n160, ZN => n307);
   U204 : NAND2_X1 port map( A1 => n310, A2 => n309, ZN => Y(7));
   U205 : AOI22_X1 port map( A1 => A_neg(7), A2 => n156, B1 => A_signal(7), B2 
                           => n147, ZN => n310);
   U206 : AOI222_X1 port map( A1 => A_shifted(7), A2 => n182, B1 => 
                           zeroSignal(7), B2 => n173, C1 => A_neg_shifted(7), 
                           C2 => n160, ZN => n309);
   U207 : NAND2_X1 port map( A1 => n312, A2 => n311, ZN => Y(8));
   U208 : AOI22_X1 port map( A1 => A_neg(8), A2 => n156, B1 => A_signal(8), B2 
                           => n147, ZN => n312);
   U209 : AOI222_X1 port map( A1 => A_shifted(8), A2 => n182, B1 => 
                           zeroSignal(8), B2 => n173, C1 => A_neg_shifted(8), 
                           C2 => n160, ZN => n311);
   U210 : NAND2_X1 port map( A1 => n318, A2 => n317, ZN => Y(9));
   U211 : AOI22_X1 port map( A1 => A_neg(9), A2 => n156, B1 => A_signal(9), B2 
                           => n147, ZN => n318);
   U212 : AOI222_X1 port map( A1 => A_shifted(9), A2 => n182, B1 => 
                           zeroSignal(9), B2 => n173, C1 => A_neg_shifted(9), 
                           C2 => n160, ZN => n317);
   U213 : NAND2_X1 port map( A1 => n190, A2 => n189, ZN => Y(10));
   U214 : AOI22_X1 port map( A1 => A_neg(10), A2 => n151, B1 => A_signal(10), 
                           B2 => n142, ZN => n190);
   U215 : AOI222_X1 port map( A1 => A_shifted(10), A2 => n177, B1 => 
                           zeroSignal(10), B2 => n168, C1 => A_neg_shifted(10),
                           C2 => n165, ZN => n189);
   U216 : NAND2_X1 port map( A1 => n192, A2 => n191, ZN => Y(11));
   U217 : AOI22_X1 port map( A1 => A_neg(11), A2 => n151, B1 => A_signal(11), 
                           B2 => n142, ZN => n192);
   U218 : AOI222_X1 port map( A1 => A_shifted(11), A2 => n177, B1 => 
                           zeroSignal(11), B2 => n168, C1 => A_neg_shifted(11),
                           C2 => n165, ZN => n191);
   U219 : NAND2_X1 port map( A1 => n194, A2 => n193, ZN => Y(12));
   U220 : AOI22_X1 port map( A1 => A_neg(12), A2 => n151, B1 => A_signal(12), 
                           B2 => n142, ZN => n194);
   U221 : AOI222_X1 port map( A1 => A_shifted(12), A2 => n177, B1 => 
                           zeroSignal(12), B2 => n168, C1 => A_neg_shifted(12),
                           C2 => n165, ZN => n193);
   U222 : NAND2_X1 port map( A1 => n196, A2 => n195, ZN => Y(13));
   U223 : AOI22_X1 port map( A1 => A_neg(13), A2 => n151, B1 => A_signal(13), 
                           B2 => n142, ZN => n196);
   U224 : AOI222_X1 port map( A1 => A_shifted(13), A2 => n177, B1 => 
                           zeroSignal(13), B2 => n168, C1 => A_neg_shifted(13),
                           C2 => n164, ZN => n195);
   U225 : NAND2_X1 port map( A1 => n198, A2 => n197, ZN => Y(14));
   U226 : AOI22_X1 port map( A1 => A_neg(14), A2 => n151, B1 => A_signal(14), 
                           B2 => n142, ZN => n198);
   U227 : AOI222_X1 port map( A1 => A_shifted(14), A2 => n177, B1 => 
                           zeroSignal(14), B2 => n168, C1 => A_neg_shifted(14),
                           C2 => n164, ZN => n197);
   U228 : NAND2_X1 port map( A1 => n200, A2 => n199, ZN => Y(15));
   U229 : AOI22_X1 port map( A1 => A_neg(15), A2 => n151, B1 => A_signal(15), 
                           B2 => n142, ZN => n200);
   U230 : AOI222_X1 port map( A1 => A_shifted(15), A2 => n177, B1 => 
                           zeroSignal(15), B2 => n168, C1 => A_neg_shifted(15),
                           C2 => n164, ZN => n199);
   U231 : NAND2_X1 port map( A1 => n202, A2 => n201, ZN => Y(16));
   U232 : AOI22_X1 port map( A1 => A_neg(16), A2 => n151, B1 => A_signal(16), 
                           B2 => n142, ZN => n202);
   U233 : AOI222_X1 port map( A1 => A_shifted(16), A2 => n177, B1 => 
                           zeroSignal(16), B2 => n168, C1 => A_neg_shifted(16),
                           C2 => n164, ZN => n201);
   U234 : NAND2_X1 port map( A1 => n204, A2 => n203, ZN => Y(17));
   U235 : AOI22_X1 port map( A1 => A_neg(17), A2 => n151, B1 => A_signal(17), 
                           B2 => n142, ZN => n204);
   U236 : AOI222_X1 port map( A1 => A_shifted(17), A2 => n177, B1 => 
                           zeroSignal(17), B2 => n168, C1 => A_neg_shifted(17),
                           C2 => n164, ZN => n203);
   U237 : NAND2_X1 port map( A1 => n206, A2 => n205, ZN => Y(18));
   U238 : AOI22_X1 port map( A1 => A_neg(18), A2 => n151, B1 => A_signal(18), 
                           B2 => n142, ZN => n206);
   U239 : AOI222_X1 port map( A1 => A_shifted(18), A2 => n177, B1 => 
                           zeroSignal(18), B2 => n168, C1 => A_neg_shifted(18),
                           C2 => n164, ZN => n205);
   U240 : NAND2_X1 port map( A1 => n208, A2 => n207, ZN => Y(19));
   U241 : AOI22_X1 port map( A1 => A_neg(19), A2 => n151, B1 => A_signal(19), 
                           B2 => n142, ZN => n208);
   U242 : AOI222_X1 port map( A1 => A_shifted(19), A2 => n177, B1 => 
                           zeroSignal(19), B2 => n168, C1 => A_neg_shifted(19),
                           C2 => n164, ZN => n207);
   U243 : AOI222_X1 port map( A1 => A_shifted(21), A2 => n178, B1 => 
                           zeroSignal(21), B2 => n169, C1 => A_neg_shifted(21),
                           C2 => n164, ZN => n213);
   U244 : AOI22_X1 port map( A1 => A_neg(20), A2 => n152, B1 => A_signal(20), 
                           B2 => n143, ZN => n212);

end SYN_BEHAVIORAL_2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity MUX51_MuxNbit64_21 is

   port( zeroSignal, A_signal, A_neg, A_shifted, A_neg_shifted : in 
         std_logic_vector (63 downto 0);  Sel : in std_logic_vector (2 downto 
         0);  Y : out std_logic_vector (63 downto 0));

end MUX51_MuxNbit64_21;

architecture SYN_BEHAVIORAL_2 of MUX51_MuxNbit64_21 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, 
      n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, 
      n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, 
      n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, 
      n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, 
      n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, 
      n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, 
      n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, 
      n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, 
      n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, 
      n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, 
      n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, 
      n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, 
      n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, 
      n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, 
      n320 : std_logic;

begin
   
   U1 : AND3_X1 port map( A1 => n319, A2 => n320, A3 => Sel(2), ZN => n141);
   U2 : BUF_X1 port map( A => n141, Z => n166);
   U3 : BUF_X1 port map( A => n185, Z => n184);
   U4 : BUF_X1 port map( A => n159, Z => n158);
   U5 : BUF_X1 port map( A => n150, Z => n149);
   U6 : BUF_X1 port map( A => n141, Z => n167);
   U7 : BUF_X1 port map( A => n185, Z => n183);
   U8 : BUF_X1 port map( A => n159, Z => n157);
   U9 : BUF_X1 port map( A => n150, Z => n148);
   U10 : BUF_X1 port map( A => n176, Z => n175);
   U11 : BUF_X1 port map( A => n176, Z => n174);
   U12 : BUF_X1 port map( A => n158, Z => n152);
   U13 : BUF_X1 port map( A => n184, Z => n178);
   U14 : BUF_X1 port map( A => n149, Z => n143);
   U15 : BUF_X1 port map( A => n166, Z => n164);
   U16 : BUF_X1 port map( A => n166, Z => n163);
   U17 : BUF_X1 port map( A => n184, Z => n179);
   U18 : BUF_X1 port map( A => n158, Z => n153);
   U19 : BUF_X1 port map( A => n149, Z => n144);
   U20 : BUF_X1 port map( A => n167, Z => n162);
   U21 : BUF_X1 port map( A => n183, Z => n180);
   U22 : BUF_X1 port map( A => n157, Z => n154);
   U23 : BUF_X1 port map( A => n148, Z => n145);
   U24 : BUF_X1 port map( A => n167, Z => n161);
   U25 : BUF_X1 port map( A => n183, Z => n181);
   U26 : BUF_X1 port map( A => n157, Z => n155);
   U27 : BUF_X1 port map( A => n148, Z => n146);
   U28 : BUF_X1 port map( A => n167, Z => n160);
   U29 : BUF_X1 port map( A => n158, Z => n151);
   U30 : BUF_X1 port map( A => n149, Z => n142);
   U31 : BUF_X1 port map( A => n175, Z => n168);
   U32 : BUF_X1 port map( A => n175, Z => n170);
   U33 : BUF_X1 port map( A => n174, Z => n171);
   U34 : BUF_X1 port map( A => n174, Z => n172);
   U35 : BUF_X1 port map( A => n175, Z => n169);
   U36 : BUF_X1 port map( A => n184, Z => n177);
   U37 : BUF_X1 port map( A => n166, Z => n165);
   U38 : BUF_X1 port map( A => n157, Z => n156);
   U39 : BUF_X1 port map( A => n148, Z => n147);
   U40 : BUF_X1 port map( A => n174, Z => n173);
   U41 : BUF_X1 port map( A => n183, Z => n182);
   U42 : INV_X1 port map( A => Sel(1), ZN => n320);
   U43 : BUF_X1 port map( A => n314, Z => n159);
   U44 : NOR3_X1 port map( A1 => Sel(0), A2 => Sel(2), A3 => n320, ZN => n314);
   U45 : BUF_X1 port map( A => n316, Z => n185);
   U46 : NOR3_X1 port map( A1 => n319, A2 => Sel(2), A3 => n320, ZN => n316);
   U47 : INV_X1 port map( A => Sel(0), ZN => n319);
   U48 : BUF_X1 port map( A => n313, Z => n150);
   U49 : NOR3_X1 port map( A1 => Sel(1), A2 => Sel(2), A3 => n319, ZN => n313);
   U50 : BUF_X1 port map( A => n315, Z => n176);
   U51 : NOR2_X1 port map( A1 => n165, A2 => n186, ZN => n315);
   U52 : AOI21_X1 port map( B1 => n319, B2 => n320, A => Sel(2), ZN => n186);
   U53 : NAND2_X1 port map( A1 => n218, A2 => n217, ZN => Y(23));
   U54 : AOI22_X1 port map( A1 => A_neg(23), A2 => n152, B1 => A_signal(23), B2
                           => n143, ZN => n218);
   U55 : NAND2_X1 port map( A1 => n216, A2 => n215, ZN => Y(22));
   U56 : AOI222_X1 port map( A1 => A_shifted(22), A2 => n178, B1 => 
                           zeroSignal(22), B2 => n169, C1 => A_neg_shifted(22),
                           C2 => n164, ZN => n215);
   U57 : NAND2_X1 port map( A1 => n220, A2 => n219, ZN => Y(24));
   U58 : AOI22_X1 port map( A1 => A_neg(24), A2 => n152, B1 => A_signal(24), B2
                           => n143, ZN => n220);
   U59 : AOI222_X1 port map( A1 => A_shifted(24), A2 => n178, B1 => 
                           zeroSignal(24), B2 => n169, C1 => A_neg_shifted(24),
                           C2 => n163, ZN => n219);
   U60 : NAND2_X1 port map( A1 => n222, A2 => n221, ZN => Y(25));
   U61 : AOI22_X1 port map( A1 => A_neg(25), A2 => n152, B1 => A_signal(25), B2
                           => n143, ZN => n222);
   U62 : AOI222_X1 port map( A1 => A_shifted(25), A2 => n178, B1 => 
                           zeroSignal(25), B2 => n169, C1 => A_neg_shifted(25),
                           C2 => n163, ZN => n221);
   U63 : NAND2_X1 port map( A1 => n224, A2 => n223, ZN => Y(26));
   U64 : AOI22_X1 port map( A1 => A_neg(26), A2 => n152, B1 => A_signal(26), B2
                           => n143, ZN => n224);
   U65 : AOI222_X1 port map( A1 => A_shifted(26), A2 => n178, B1 => 
                           zeroSignal(26), B2 => n169, C1 => A_neg_shifted(26),
                           C2 => n163, ZN => n223);
   U66 : NAND2_X1 port map( A1 => n244, A2 => n243, ZN => Y(35));
   U67 : AOI222_X1 port map( A1 => A_shifted(35), A2 => n179, B1 => 
                           zeroSignal(35), B2 => n170, C1 => A_neg_shifted(35),
                           C2 => n162, ZN => n243);
   U68 : AOI22_X1 port map( A1 => A_neg(35), A2 => n153, B1 => A_signal(35), B2
                           => n144, ZN => n244);
   U69 : NAND2_X1 port map( A1 => n238, A2 => n237, ZN => Y(32));
   U70 : AOI222_X1 port map( A1 => A_shifted(32), A2 => n179, B1 => 
                           zeroSignal(32), B2 => n170, C1 => A_neg_shifted(32),
                           C2 => n163, ZN => n237);
   U71 : AOI22_X1 port map( A1 => A_neg(32), A2 => n153, B1 => A_signal(32), B2
                           => n144, ZN => n238);
   U72 : NAND2_X1 port map( A1 => n242, A2 => n241, ZN => Y(34));
   U73 : AOI222_X1 port map( A1 => A_shifted(34), A2 => n179, B1 => 
                           zeroSignal(34), B2 => n170, C1 => A_neg_shifted(34),
                           C2 => n163, ZN => n241);
   U74 : AOI22_X1 port map( A1 => A_neg(34), A2 => n153, B1 => A_signal(34), B2
                           => n144, ZN => n242);
   U75 : NAND2_X1 port map( A1 => n240, A2 => n239, ZN => Y(33));
   U76 : AOI222_X1 port map( A1 => A_shifted(33), A2 => n179, B1 => 
                           zeroSignal(33), B2 => n170, C1 => A_neg_shifted(33),
                           C2 => n163, ZN => n239);
   U77 : AOI22_X1 port map( A1 => A_neg(33), A2 => n153, B1 => A_signal(33), B2
                           => n144, ZN => n240);
   U78 : NAND2_X1 port map( A1 => n248, A2 => n247, ZN => Y(37));
   U79 : AOI222_X1 port map( A1 => A_shifted(37), A2 => n179, B1 => 
                           zeroSignal(37), B2 => n170, C1 => A_neg_shifted(37),
                           C2 => n162, ZN => n247);
   U80 : AOI22_X1 port map( A1 => A_neg(37), A2 => n153, B1 => A_signal(37), B2
                           => n144, ZN => n248);
   U81 : NAND2_X1 port map( A1 => n250, A2 => n249, ZN => Y(38));
   U82 : AOI222_X1 port map( A1 => A_shifted(38), A2 => n179, B1 => 
                           zeroSignal(38), B2 => n170, C1 => A_neg_shifted(38),
                           C2 => n162, ZN => n249);
   U83 : AOI22_X1 port map( A1 => A_neg(38), A2 => n153, B1 => A_signal(38), B2
                           => n144, ZN => n250);
   U84 : NAND2_X1 port map( A1 => n252, A2 => n251, ZN => Y(39));
   U85 : AOI222_X1 port map( A1 => A_shifted(39), A2 => n179, B1 => 
                           zeroSignal(39), B2 => n170, C1 => A_neg_shifted(39),
                           C2 => n162, ZN => n251);
   U86 : AOI22_X1 port map( A1 => A_neg(39), A2 => n153, B1 => A_signal(39), B2
                           => n144, ZN => n252);
   U87 : NAND2_X1 port map( A1 => n258, A2 => n257, ZN => Y(41));
   U88 : AOI222_X1 port map( A1 => A_shifted(41), A2 => n179, B1 => 
                           zeroSignal(41), B2 => n170, C1 => A_neg_shifted(41),
                           C2 => n162, ZN => n257);
   U89 : AOI22_X1 port map( A1 => A_neg(41), A2 => n153, B1 => A_signal(41), B2
                           => n144, ZN => n258);
   U90 : NAND2_X1 port map( A1 => n246, A2 => n245, ZN => Y(36));
   U91 : AOI22_X1 port map( A1 => A_neg(36), A2 => n153, B1 => A_signal(36), B2
                           => n144, ZN => n246);
   U92 : AOI222_X1 port map( A1 => A_shifted(36), A2 => n179, B1 => 
                           zeroSignal(36), B2 => n170, C1 => A_neg_shifted(36),
                           C2 => n162, ZN => n245);
   U93 : NAND2_X1 port map( A1 => n226, A2 => n225, ZN => Y(27));
   U94 : AOI22_X1 port map( A1 => A_neg(27), A2 => n152, B1 => A_signal(27), B2
                           => n143, ZN => n226);
   U95 : AOI222_X1 port map( A1 => A_shifted(27), A2 => n178, B1 => 
                           zeroSignal(27), B2 => n169, C1 => A_neg_shifted(27),
                           C2 => n163, ZN => n225);
   U96 : NAND2_X1 port map( A1 => n260, A2 => n259, ZN => Y(42));
   U97 : AOI222_X1 port map( A1 => A_shifted(42), A2 => n180, B1 => 
                           zeroSignal(42), B2 => n171, C1 => A_neg_shifted(42),
                           C2 => n162, ZN => n259);
   U98 : AOI22_X1 port map( A1 => A_neg(42), A2 => n154, B1 => A_signal(42), B2
                           => n145, ZN => n260);
   U99 : NAND2_X1 port map( A1 => n264, A2 => n263, ZN => Y(44));
   U100 : AOI222_X1 port map( A1 => A_shifted(44), A2 => n180, B1 => 
                           zeroSignal(44), B2 => n171, C1 => A_neg_shifted(44),
                           C2 => n162, ZN => n263);
   U101 : AOI22_X1 port map( A1 => A_neg(44), A2 => n154, B1 => A_signal(44), 
                           B2 => n145, ZN => n264);
   U102 : NAND2_X1 port map( A1 => n262, A2 => n261, ZN => Y(43));
   U103 : AOI222_X1 port map( A1 => A_shifted(43), A2 => n180, B1 => 
                           zeroSignal(43), B2 => n171, C1 => A_neg_shifted(43),
                           C2 => n162, ZN => n261);
   U104 : AOI22_X1 port map( A1 => A_neg(43), A2 => n154, B1 => A_signal(43), 
                           B2 => n145, ZN => n262);
   U105 : NAND2_X1 port map( A1 => n266, A2 => n265, ZN => Y(45));
   U106 : AOI222_X1 port map( A1 => A_shifted(45), A2 => n180, B1 => 
                           zeroSignal(45), B2 => n171, C1 => A_neg_shifted(45),
                           C2 => n162, ZN => n265);
   U107 : AOI22_X1 port map( A1 => A_neg(45), A2 => n154, B1 => A_signal(45), 
                           B2 => n145, ZN => n266);
   U108 : NAND2_X1 port map( A1 => n256, A2 => n255, ZN => Y(40));
   U109 : AOI22_X1 port map( A1 => A_neg(40), A2 => n153, B1 => A_signal(40), 
                           B2 => n144, ZN => n256);
   U110 : AOI222_X1 port map( A1 => A_shifted(40), A2 => n179, B1 => 
                           zeroSignal(40), B2 => n170, C1 => A_neg_shifted(40),
                           C2 => n162, ZN => n255);
   U111 : NAND2_X1 port map( A1 => n270, A2 => n269, ZN => Y(47));
   U112 : AOI222_X1 port map( A1 => A_shifted(47), A2 => n180, B1 => 
                           zeroSignal(47), B2 => n171, C1 => A_neg_shifted(47),
                           C2 => n161, ZN => n269);
   U113 : AOI22_X1 port map( A1 => A_neg(47), A2 => n154, B1 => A_signal(47), 
                           B2 => n145, ZN => n270);
   U114 : NAND2_X1 port map( A1 => n274, A2 => n273, ZN => Y(49));
   U115 : AOI222_X1 port map( A1 => A_shifted(49), A2 => n180, B1 => 
                           zeroSignal(49), B2 => n171, C1 => A_neg_shifted(49),
                           C2 => n161, ZN => n273);
   U116 : AOI22_X1 port map( A1 => A_neg(49), A2 => n154, B1 => A_signal(49), 
                           B2 => n145, ZN => n274);
   U117 : NAND2_X1 port map( A1 => n272, A2 => n271, ZN => Y(48));
   U118 : AOI222_X1 port map( A1 => A_shifted(48), A2 => n180, B1 => 
                           zeroSignal(48), B2 => n171, C1 => A_neg_shifted(48),
                           C2 => n161, ZN => n271);
   U119 : AOI22_X1 port map( A1 => A_neg(48), A2 => n154, B1 => A_signal(48), 
                           B2 => n145, ZN => n272);
   U120 : NAND2_X1 port map( A1 => n288, A2 => n287, ZN => Y(55));
   U121 : AOI222_X1 port map( A1 => A_shifted(55), A2 => n181, B1 => 
                           zeroSignal(55), B2 => n172, C1 => A_neg_shifted(55),
                           C2 => n161, ZN => n287);
   U122 : AOI22_X1 port map( A1 => A_neg(55), A2 => n155, B1 => A_signal(55), 
                           B2 => n146, ZN => n288);
   U123 : NAND2_X1 port map( A1 => n282, A2 => n281, ZN => Y(52));
   U124 : AOI222_X1 port map( A1 => A_shifted(52), A2 => n180, B1 => 
                           zeroSignal(52), B2 => n171, C1 => A_neg_shifted(52),
                           C2 => n161, ZN => n281);
   U125 : AOI22_X1 port map( A1 => A_neg(52), A2 => n154, B1 => A_signal(52), 
                           B2 => n145, ZN => n282);
   U126 : NAND2_X1 port map( A1 => n278, A2 => n277, ZN => Y(50));
   U127 : AOI222_X1 port map( A1 => A_shifted(50), A2 => n180, B1 => 
                           zeroSignal(50), B2 => n171, C1 => A_neg_shifted(50),
                           C2 => n161, ZN => n277);
   U128 : AOI22_X1 port map( A1 => A_neg(50), A2 => n154, B1 => A_signal(50), 
                           B2 => n145, ZN => n278);
   U129 : NAND2_X1 port map( A1 => n280, A2 => n279, ZN => Y(51));
   U130 : AOI222_X1 port map( A1 => A_shifted(51), A2 => n180, B1 => 
                           zeroSignal(51), B2 => n171, C1 => A_neg_shifted(51),
                           C2 => n161, ZN => n279);
   U131 : AOI22_X1 port map( A1 => A_neg(51), A2 => n154, B1 => A_signal(51), 
                           B2 => n145, ZN => n280);
   U132 : NAND2_X1 port map( A1 => n228, A2 => n227, ZN => Y(28));
   U133 : AOI222_X1 port map( A1 => A_shifted(28), A2 => n178, B1 => 
                           zeroSignal(28), B2 => n169, C1 => A_neg_shifted(28),
                           C2 => n163, ZN => n227);
   U134 : AOI22_X1 port map( A1 => A_neg(28), A2 => n152, B1 => A_signal(28), 
                           B2 => n143, ZN => n228);
   U135 : NAND2_X1 port map( A1 => n284, A2 => n283, ZN => Y(53));
   U136 : AOI222_X1 port map( A1 => A_shifted(53), A2 => n181, B1 => 
                           zeroSignal(53), B2 => n172, C1 => A_neg_shifted(53),
                           C2 => n161, ZN => n283);
   U137 : AOI22_X1 port map( A1 => A_neg(53), A2 => n155, B1 => A_signal(53), 
                           B2 => n146, ZN => n284);
   U138 : NAND2_X1 port map( A1 => n230, A2 => n229, ZN => Y(29));
   U139 : AOI222_X1 port map( A1 => A_shifted(29), A2 => n178, B1 => 
                           zeroSignal(29), B2 => n169, C1 => A_neg_shifted(29),
                           C2 => n163, ZN => n229);
   U140 : AOI22_X1 port map( A1 => A_neg(29), A2 => n152, B1 => A_signal(29), 
                           B2 => n143, ZN => n230);
   U141 : NAND2_X1 port map( A1 => n268, A2 => n267, ZN => Y(46));
   U142 : AOI22_X1 port map( A1 => A_neg(46), A2 => n154, B1 => A_signal(46), 
                           B2 => n145, ZN => n268);
   U143 : AOI222_X1 port map( A1 => A_shifted(46), A2 => n180, B1 => 
                           zeroSignal(46), B2 => n171, C1 => A_neg_shifted(46),
                           C2 => n161, ZN => n267);
   U144 : NAND2_X1 port map( A1 => n286, A2 => n285, ZN => Y(54));
   U145 : AOI222_X1 port map( A1 => A_shifted(54), A2 => n181, B1 => 
                           zeroSignal(54), B2 => n172, C1 => A_neg_shifted(54),
                           C2 => n161, ZN => n285);
   U146 : AOI22_X1 port map( A1 => A_neg(54), A2 => n155, B1 => A_signal(54), 
                           B2 => n146, ZN => n286);
   U147 : NAND2_X1 port map( A1 => n234, A2 => n233, ZN => Y(30));
   U148 : AOI222_X1 port map( A1 => A_shifted(30), A2 => n178, B1 => 
                           zeroSignal(30), B2 => n169, C1 => A_neg_shifted(30),
                           C2 => n163, ZN => n233);
   U149 : AOI22_X1 port map( A1 => A_neg(30), A2 => n152, B1 => A_signal(30), 
                           B2 => n143, ZN => n234);
   U150 : NAND2_X1 port map( A1 => n236, A2 => n235, ZN => Y(31));
   U151 : AOI222_X1 port map( A1 => A_shifted(31), A2 => n179, B1 => 
                           zeroSignal(31), B2 => n170, C1 => A_neg_shifted(31),
                           C2 => n163, ZN => n235);
   U152 : AOI22_X1 port map( A1 => A_neg(31), A2 => n153, B1 => A_signal(31), 
                           B2 => n144, ZN => n236);
   U153 : NAND2_X1 port map( A1 => n290, A2 => n289, ZN => Y(56));
   U154 : AOI222_X1 port map( A1 => A_shifted(56), A2 => n181, B1 => 
                           zeroSignal(56), B2 => n172, C1 => A_neg_shifted(56),
                           C2 => n161, ZN => n289);
   U155 : AOI22_X1 port map( A1 => A_neg(56), A2 => n155, B1 => A_signal(56), 
                           B2 => n146, ZN => n290);
   U156 : NAND2_X1 port map( A1 => n292, A2 => n291, ZN => Y(57));
   U157 : AOI222_X1 port map( A1 => A_shifted(57), A2 => n181, B1 => 
                           zeroSignal(57), B2 => n172, C1 => A_neg_shifted(57),
                           C2 => n160, ZN => n291);
   U158 : AOI22_X1 port map( A1 => A_neg(57), A2 => n155, B1 => A_signal(57), 
                           B2 => n146, ZN => n292);
   U159 : NAND2_X1 port map( A1 => n294, A2 => n293, ZN => Y(58));
   U160 : AOI222_X1 port map( A1 => A_shifted(58), A2 => n181, B1 => 
                           zeroSignal(58), B2 => n172, C1 => A_neg_shifted(58),
                           C2 => n160, ZN => n293);
   U161 : AOI22_X1 port map( A1 => A_neg(58), A2 => n155, B1 => A_signal(58), 
                           B2 => n146, ZN => n294);
   U162 : NAND2_X1 port map( A1 => n296, A2 => n295, ZN => Y(59));
   U163 : AOI22_X1 port map( A1 => A_neg(59), A2 => n155, B1 => A_signal(59), 
                           B2 => n146, ZN => n296);
   U164 : AOI222_X1 port map( A1 => A_shifted(59), A2 => n181, B1 => 
                           zeroSignal(59), B2 => n172, C1 => A_neg_shifted(59),
                           C2 => n160, ZN => n295);
   U165 : NAND2_X1 port map( A1 => n304, A2 => n303, ZN => Y(62));
   U166 : AOI222_X1 port map( A1 => A_shifted(62), A2 => n181, B1 => 
                           zeroSignal(62), B2 => n172, C1 => A_neg_shifted(62),
                           C2 => n160, ZN => n303);
   U167 : AOI22_X1 port map( A1 => A_neg(62), A2 => n155, B1 => A_signal(62), 
                           B2 => n146, ZN => n304);
   U168 : NAND2_X1 port map( A1 => n302, A2 => n301, ZN => Y(61));
   U169 : AOI222_X1 port map( A1 => A_shifted(61), A2 => n181, B1 => 
                           zeroSignal(61), B2 => n172, C1 => A_neg_shifted(61),
                           C2 => n160, ZN => n301);
   U170 : AOI22_X1 port map( A1 => A_neg(61), A2 => n155, B1 => A_signal(61), 
                           B2 => n146, ZN => n302);
   U171 : NAND2_X1 port map( A1 => n300, A2 => n299, ZN => Y(60));
   U172 : AOI222_X1 port map( A1 => A_shifted(60), A2 => n181, B1 => 
                           zeroSignal(60), B2 => n172, C1 => A_neg_shifted(60),
                           C2 => n160, ZN => n299);
   U173 : AOI22_X1 port map( A1 => A_neg(60), A2 => n155, B1 => A_signal(60), 
                           B2 => n146, ZN => n300);
   U174 : NAND2_X1 port map( A1 => n306, A2 => n305, ZN => Y(63));
   U175 : AOI22_X1 port map( A1 => A_neg(63), A2 => n155, B1 => A_signal(63), 
                           B2 => n146, ZN => n306);
   U176 : AOI222_X1 port map( A1 => A_shifted(63), A2 => n181, B1 => 
                           zeroSignal(63), B2 => n172, C1 => A_neg_shifted(63),
                           C2 => n160, ZN => n305);
   U177 : NAND2_X1 port map( A1 => n188, A2 => n187, ZN => Y(0));
   U178 : AOI22_X1 port map( A1 => A_neg(0), A2 => n151, B1 => A_signal(0), B2 
                           => n142, ZN => n188);
   U179 : AOI222_X1 port map( A1 => A_shifted(0), A2 => n177, B1 => 
                           zeroSignal(0), B2 => n168, C1 => A_neg_shifted(0), 
                           C2 => n165, ZN => n187);
   U180 : NAND2_X1 port map( A1 => n210, A2 => n209, ZN => Y(1));
   U181 : AOI22_X1 port map( A1 => A_neg(1), A2 => n151, B1 => A_signal(1), B2 
                           => n142, ZN => n210);
   U182 : AOI222_X1 port map( A1 => A_shifted(1), A2 => n177, B1 => 
                           zeroSignal(1), B2 => n168, C1 => A_neg_shifted(1), 
                           C2 => n164, ZN => n209);
   U183 : NAND2_X1 port map( A1 => n232, A2 => n231, ZN => Y(2));
   U184 : AOI22_X1 port map( A1 => A_neg(2), A2 => n152, B1 => A_signal(2), B2 
                           => n143, ZN => n232);
   U185 : AOI222_X1 port map( A1 => A_shifted(2), A2 => n178, B1 => 
                           zeroSignal(2), B2 => n169, C1 => A_neg_shifted(2), 
                           C2 => n163, ZN => n231);
   U186 : NAND2_X1 port map( A1 => n254, A2 => n253, ZN => Y(3));
   U187 : AOI22_X1 port map( A1 => A_neg(3), A2 => n153, B1 => A_signal(3), B2 
                           => n144, ZN => n254);
   U188 : AOI222_X1 port map( A1 => A_shifted(3), A2 => n179, B1 => 
                           zeroSignal(3), B2 => n170, C1 => A_neg_shifted(3), 
                           C2 => n162, ZN => n253);
   U189 : NAND2_X1 port map( A1 => n276, A2 => n275, ZN => Y(4));
   U190 : AOI22_X1 port map( A1 => A_neg(4), A2 => n154, B1 => A_signal(4), B2 
                           => n145, ZN => n276);
   U191 : AOI222_X1 port map( A1 => A_shifted(4), A2 => n180, B1 => 
                           zeroSignal(4), B2 => n171, C1 => A_neg_shifted(4), 
                           C2 => n161, ZN => n275);
   U192 : NAND2_X1 port map( A1 => n298, A2 => n297, ZN => Y(5));
   U193 : AOI22_X1 port map( A1 => A_neg(5), A2 => n155, B1 => A_signal(5), B2 
                           => n146, ZN => n298);
   U194 : AOI222_X1 port map( A1 => A_shifted(5), A2 => n181, B1 => 
                           zeroSignal(5), B2 => n172, C1 => A_neg_shifted(5), 
                           C2 => n160, ZN => n297);
   U195 : NAND2_X1 port map( A1 => n308, A2 => n307, ZN => Y(6));
   U196 : AOI22_X1 port map( A1 => A_neg(6), A2 => n156, B1 => A_signal(6), B2 
                           => n147, ZN => n308);
   U197 : AOI222_X1 port map( A1 => A_shifted(6), A2 => n182, B1 => 
                           zeroSignal(6), B2 => n173, C1 => A_neg_shifted(6), 
                           C2 => n160, ZN => n307);
   U198 : NAND2_X1 port map( A1 => n310, A2 => n309, ZN => Y(7));
   U199 : AOI22_X1 port map( A1 => A_neg(7), A2 => n156, B1 => A_signal(7), B2 
                           => n147, ZN => n310);
   U200 : AOI222_X1 port map( A1 => A_shifted(7), A2 => n182, B1 => 
                           zeroSignal(7), B2 => n173, C1 => A_neg_shifted(7), 
                           C2 => n160, ZN => n309);
   U201 : NAND2_X1 port map( A1 => n312, A2 => n311, ZN => Y(8));
   U202 : AOI22_X1 port map( A1 => A_neg(8), A2 => n156, B1 => A_signal(8), B2 
                           => n147, ZN => n312);
   U203 : AOI222_X1 port map( A1 => A_shifted(8), A2 => n182, B1 => 
                           zeroSignal(8), B2 => n173, C1 => A_neg_shifted(8), 
                           C2 => n160, ZN => n311);
   U204 : NAND2_X1 port map( A1 => n318, A2 => n317, ZN => Y(9));
   U205 : AOI22_X1 port map( A1 => A_neg(9), A2 => n156, B1 => A_signal(9), B2 
                           => n147, ZN => n318);
   U206 : AOI222_X1 port map( A1 => A_shifted(9), A2 => n182, B1 => 
                           zeroSignal(9), B2 => n173, C1 => A_neg_shifted(9), 
                           C2 => n160, ZN => n317);
   U207 : NAND2_X1 port map( A1 => n190, A2 => n189, ZN => Y(10));
   U208 : AOI22_X1 port map( A1 => A_neg(10), A2 => n151, B1 => A_signal(10), 
                           B2 => n142, ZN => n190);
   U209 : AOI222_X1 port map( A1 => A_shifted(10), A2 => n177, B1 => 
                           zeroSignal(10), B2 => n168, C1 => A_neg_shifted(10),
                           C2 => n165, ZN => n189);
   U210 : NAND2_X1 port map( A1 => n192, A2 => n191, ZN => Y(11));
   U211 : AOI22_X1 port map( A1 => A_neg(11), A2 => n151, B1 => A_signal(11), 
                           B2 => n142, ZN => n192);
   U212 : AOI222_X1 port map( A1 => A_shifted(11), A2 => n177, B1 => 
                           zeroSignal(11), B2 => n168, C1 => A_neg_shifted(11),
                           C2 => n165, ZN => n191);
   U213 : NAND2_X1 port map( A1 => n194, A2 => n193, ZN => Y(12));
   U214 : AOI22_X1 port map( A1 => A_neg(12), A2 => n151, B1 => A_signal(12), 
                           B2 => n142, ZN => n194);
   U215 : AOI222_X1 port map( A1 => A_shifted(12), A2 => n177, B1 => 
                           zeroSignal(12), B2 => n168, C1 => A_neg_shifted(12),
                           C2 => n165, ZN => n193);
   U216 : NAND2_X1 port map( A1 => n196, A2 => n195, ZN => Y(13));
   U217 : AOI22_X1 port map( A1 => A_neg(13), A2 => n151, B1 => A_signal(13), 
                           B2 => n142, ZN => n196);
   U218 : AOI222_X1 port map( A1 => A_shifted(13), A2 => n177, B1 => 
                           zeroSignal(13), B2 => n168, C1 => A_neg_shifted(13),
                           C2 => n164, ZN => n195);
   U219 : NAND2_X1 port map( A1 => n198, A2 => n197, ZN => Y(14));
   U220 : AOI22_X1 port map( A1 => A_neg(14), A2 => n151, B1 => A_signal(14), 
                           B2 => n142, ZN => n198);
   U221 : AOI222_X1 port map( A1 => A_shifted(14), A2 => n177, B1 => 
                           zeroSignal(14), B2 => n168, C1 => A_neg_shifted(14),
                           C2 => n164, ZN => n197);
   U222 : NAND2_X1 port map( A1 => n200, A2 => n199, ZN => Y(15));
   U223 : AOI22_X1 port map( A1 => A_neg(15), A2 => n151, B1 => A_signal(15), 
                           B2 => n142, ZN => n200);
   U224 : AOI222_X1 port map( A1 => A_shifted(15), A2 => n177, B1 => 
                           zeroSignal(15), B2 => n168, C1 => A_neg_shifted(15),
                           C2 => n164, ZN => n199);
   U225 : NAND2_X1 port map( A1 => n202, A2 => n201, ZN => Y(16));
   U226 : AOI22_X1 port map( A1 => A_neg(16), A2 => n151, B1 => A_signal(16), 
                           B2 => n142, ZN => n202);
   U227 : AOI222_X1 port map( A1 => A_shifted(16), A2 => n177, B1 => 
                           zeroSignal(16), B2 => n168, C1 => A_neg_shifted(16),
                           C2 => n164, ZN => n201);
   U228 : NAND2_X1 port map( A1 => n204, A2 => n203, ZN => Y(17));
   U229 : AOI22_X1 port map( A1 => A_neg(17), A2 => n151, B1 => A_signal(17), 
                           B2 => n142, ZN => n204);
   U230 : AOI222_X1 port map( A1 => A_shifted(17), A2 => n177, B1 => 
                           zeroSignal(17), B2 => n168, C1 => A_neg_shifted(17),
                           C2 => n164, ZN => n203);
   U231 : NAND2_X1 port map( A1 => n206, A2 => n205, ZN => Y(18));
   U232 : AOI22_X1 port map( A1 => A_neg(18), A2 => n151, B1 => A_signal(18), 
                           B2 => n142, ZN => n206);
   U233 : AOI222_X1 port map( A1 => A_shifted(18), A2 => n177, B1 => 
                           zeroSignal(18), B2 => n168, C1 => A_neg_shifted(18),
                           C2 => n164, ZN => n205);
   U234 : NAND2_X1 port map( A1 => n208, A2 => n207, ZN => Y(19));
   U235 : AOI22_X1 port map( A1 => A_neg(19), A2 => n151, B1 => A_signal(19), 
                           B2 => n142, ZN => n208);
   U236 : AOI222_X1 port map( A1 => A_shifted(19), A2 => n177, B1 => 
                           zeroSignal(19), B2 => n168, C1 => A_neg_shifted(19),
                           C2 => n164, ZN => n207);
   U237 : NAND2_X1 port map( A1 => n212, A2 => n211, ZN => Y(20));
   U238 : AOI22_X1 port map( A1 => A_neg(20), A2 => n152, B1 => A_signal(20), 
                           B2 => n143, ZN => n212);
   U239 : AOI222_X1 port map( A1 => A_shifted(20), A2 => n178, B1 => 
                           zeroSignal(20), B2 => n169, C1 => A_neg_shifted(20),
                           C2 => n164, ZN => n211);
   U240 : NAND2_X1 port map( A1 => n214, A2 => n213, ZN => Y(21));
   U241 : AOI22_X1 port map( A1 => A_neg(21), A2 => n152, B1 => A_signal(21), 
                           B2 => n143, ZN => n214);
   U242 : AOI222_X1 port map( A1 => A_shifted(21), A2 => n178, B1 => 
                           zeroSignal(21), B2 => n169, C1 => A_neg_shifted(21),
                           C2 => n164, ZN => n213);
   U243 : AOI222_X1 port map( A1 => A_shifted(23), A2 => n178, B1 => 
                           zeroSignal(23), B2 => n169, C1 => A_neg_shifted(23),
                           C2 => n164, ZN => n217);
   U244 : AOI22_X1 port map( A1 => A_neg(22), A2 => n152, B1 => A_signal(22), 
                           B2 => n143, ZN => n216);

end SYN_BEHAVIORAL_2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity MUX51_MuxNbit64_20 is

   port( zeroSignal, A_signal, A_neg, A_shifted, A_neg_shifted : in 
         std_logic_vector (63 downto 0);  Sel : in std_logic_vector (2 downto 
         0);  Y : out std_logic_vector (63 downto 0));

end MUX51_MuxNbit64_20;

architecture SYN_BEHAVIORAL_2 of MUX51_MuxNbit64_20 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, 
      n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, 
      n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, 
      n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, 
      n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, 
      n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, 
      n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, 
      n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, 
      n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, 
      n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, 
      n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, 
      n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, 
      n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, 
      n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, 
      n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, 
      n320 : std_logic;

begin
   
   U1 : AND3_X1 port map( A1 => n319, A2 => n320, A3 => Sel(2), ZN => n141);
   U2 : BUF_X1 port map( A => n141, Z => n166);
   U3 : BUF_X1 port map( A => n185, Z => n184);
   U4 : BUF_X1 port map( A => n159, Z => n158);
   U5 : BUF_X1 port map( A => n150, Z => n149);
   U6 : BUF_X1 port map( A => n141, Z => n167);
   U7 : BUF_X1 port map( A => n185, Z => n183);
   U8 : BUF_X1 port map( A => n159, Z => n157);
   U9 : BUF_X1 port map( A => n150, Z => n148);
   U10 : BUF_X1 port map( A => n176, Z => n175);
   U11 : BUF_X1 port map( A => n176, Z => n174);
   U12 : BUF_X1 port map( A => n158, Z => n152);
   U13 : BUF_X1 port map( A => n184, Z => n178);
   U14 : BUF_X1 port map( A => n149, Z => n143);
   U15 : BUF_X1 port map( A => n166, Z => n163);
   U16 : BUF_X1 port map( A => n184, Z => n179);
   U17 : BUF_X1 port map( A => n158, Z => n153);
   U18 : BUF_X1 port map( A => n149, Z => n144);
   U19 : BUF_X1 port map( A => n167, Z => n162);
   U20 : BUF_X1 port map( A => n183, Z => n180);
   U21 : BUF_X1 port map( A => n157, Z => n154);
   U22 : BUF_X1 port map( A => n148, Z => n145);
   U23 : BUF_X1 port map( A => n167, Z => n161);
   U24 : BUF_X1 port map( A => n183, Z => n181);
   U25 : BUF_X1 port map( A => n157, Z => n155);
   U26 : BUF_X1 port map( A => n148, Z => n146);
   U27 : BUF_X1 port map( A => n167, Z => n160);
   U28 : BUF_X1 port map( A => n158, Z => n151);
   U29 : BUF_X1 port map( A => n149, Z => n142);
   U30 : BUF_X1 port map( A => n175, Z => n168);
   U31 : BUF_X1 port map( A => n175, Z => n170);
   U32 : BUF_X1 port map( A => n174, Z => n171);
   U33 : BUF_X1 port map( A => n174, Z => n172);
   U34 : BUF_X1 port map( A => n166, Z => n164);
   U35 : BUF_X1 port map( A => n175, Z => n169);
   U36 : BUF_X1 port map( A => n184, Z => n177);
   U37 : BUF_X1 port map( A => n166, Z => n165);
   U38 : BUF_X1 port map( A => n157, Z => n156);
   U39 : BUF_X1 port map( A => n148, Z => n147);
   U40 : BUF_X1 port map( A => n174, Z => n173);
   U41 : BUF_X1 port map( A => n183, Z => n182);
   U42 : INV_X1 port map( A => Sel(1), ZN => n320);
   U43 : BUF_X1 port map( A => n314, Z => n159);
   U44 : NOR3_X1 port map( A1 => Sel(0), A2 => Sel(2), A3 => n320, ZN => n314);
   U45 : BUF_X1 port map( A => n316, Z => n185);
   U46 : NOR3_X1 port map( A1 => n319, A2 => Sel(2), A3 => n320, ZN => n316);
   U47 : INV_X1 port map( A => Sel(0), ZN => n319);
   U48 : BUF_X1 port map( A => n313, Z => n150);
   U49 : NOR3_X1 port map( A1 => Sel(1), A2 => Sel(2), A3 => n319, ZN => n313);
   U50 : BUF_X1 port map( A => n315, Z => n176);
   U51 : NOR2_X1 port map( A1 => n165, A2 => n186, ZN => n315);
   U52 : AOI21_X1 port map( B1 => n319, B2 => n320, A => Sel(2), ZN => n186);
   U53 : NAND2_X1 port map( A1 => n222, A2 => n221, ZN => Y(25));
   U54 : AOI22_X1 port map( A1 => A_neg(25), A2 => n152, B1 => A_signal(25), B2
                           => n143, ZN => n222);
   U55 : NAND2_X1 port map( A1 => n220, A2 => n219, ZN => Y(24));
   U56 : AOI222_X1 port map( A1 => A_shifted(24), A2 => n178, B1 => 
                           zeroSignal(24), B2 => n169, C1 => A_neg_shifted(24),
                           C2 => n163, ZN => n219);
   U57 : NAND2_X1 port map( A1 => n224, A2 => n223, ZN => Y(26));
   U58 : AOI22_X1 port map( A1 => A_neg(26), A2 => n152, B1 => A_signal(26), B2
                           => n143, ZN => n224);
   U59 : AOI222_X1 port map( A1 => A_shifted(26), A2 => n178, B1 => 
                           zeroSignal(26), B2 => n169, C1 => A_neg_shifted(26),
                           C2 => n163, ZN => n223);
   U60 : NAND2_X1 port map( A1 => n226, A2 => n225, ZN => Y(27));
   U61 : AOI22_X1 port map( A1 => A_neg(27), A2 => n152, B1 => A_signal(27), B2
                           => n143, ZN => n226);
   U62 : AOI222_X1 port map( A1 => A_shifted(27), A2 => n178, B1 => 
                           zeroSignal(27), B2 => n169, C1 => A_neg_shifted(27),
                           C2 => n163, ZN => n225);
   U63 : NAND2_X1 port map( A1 => n244, A2 => n243, ZN => Y(35));
   U64 : AOI222_X1 port map( A1 => A_shifted(35), A2 => n179, B1 => 
                           zeroSignal(35), B2 => n170, C1 => A_neg_shifted(35),
                           C2 => n162, ZN => n243);
   U65 : AOI22_X1 port map( A1 => A_neg(35), A2 => n153, B1 => A_signal(35), B2
                           => n144, ZN => n244);
   U66 : NAND2_X1 port map( A1 => n228, A2 => n227, ZN => Y(28));
   U67 : AOI22_X1 port map( A1 => A_neg(28), A2 => n152, B1 => A_signal(28), B2
                           => n143, ZN => n228);
   U68 : AOI222_X1 port map( A1 => A_shifted(28), A2 => n178, B1 => 
                           zeroSignal(28), B2 => n169, C1 => A_neg_shifted(28),
                           C2 => n163, ZN => n227);
   U69 : NAND2_X1 port map( A1 => n242, A2 => n241, ZN => Y(34));
   U70 : AOI222_X1 port map( A1 => A_shifted(34), A2 => n179, B1 => 
                           zeroSignal(34), B2 => n170, C1 => A_neg_shifted(34),
                           C2 => n163, ZN => n241);
   U71 : AOI22_X1 port map( A1 => A_neg(34), A2 => n153, B1 => A_signal(34), B2
                           => n144, ZN => n242);
   U72 : NAND2_X1 port map( A1 => n248, A2 => n247, ZN => Y(37));
   U73 : AOI222_X1 port map( A1 => A_shifted(37), A2 => n179, B1 => 
                           zeroSignal(37), B2 => n170, C1 => A_neg_shifted(37),
                           C2 => n162, ZN => n247);
   U74 : AOI22_X1 port map( A1 => A_neg(37), A2 => n153, B1 => A_signal(37), B2
                           => n144, ZN => n248);
   U75 : NAND2_X1 port map( A1 => n246, A2 => n245, ZN => Y(36));
   U76 : AOI222_X1 port map( A1 => A_shifted(36), A2 => n179, B1 => 
                           zeroSignal(36), B2 => n170, C1 => A_neg_shifted(36),
                           C2 => n162, ZN => n245);
   U77 : AOI22_X1 port map( A1 => A_neg(36), A2 => n153, B1 => A_signal(36), B2
                           => n144, ZN => n246);
   U78 : NAND2_X1 port map( A1 => n256, A2 => n255, ZN => Y(40));
   U79 : AOI222_X1 port map( A1 => A_shifted(40), A2 => n179, B1 => 
                           zeroSignal(40), B2 => n170, C1 => A_neg_shifted(40),
                           C2 => n162, ZN => n255);
   U80 : AOI22_X1 port map( A1 => A_neg(40), A2 => n153, B1 => A_signal(40), B2
                           => n144, ZN => n256);
   U81 : NAND2_X1 port map( A1 => n252, A2 => n251, ZN => Y(39));
   U82 : AOI222_X1 port map( A1 => A_shifted(39), A2 => n179, B1 => 
                           zeroSignal(39), B2 => n170, C1 => A_neg_shifted(39),
                           C2 => n162, ZN => n251);
   U83 : AOI22_X1 port map( A1 => A_neg(39), A2 => n153, B1 => A_signal(39), B2
                           => n144, ZN => n252);
   U84 : NAND2_X1 port map( A1 => n258, A2 => n257, ZN => Y(41));
   U85 : AOI222_X1 port map( A1 => A_shifted(41), A2 => n179, B1 => 
                           zeroSignal(41), B2 => n170, C1 => A_neg_shifted(41),
                           C2 => n162, ZN => n257);
   U86 : AOI22_X1 port map( A1 => A_neg(41), A2 => n153, B1 => A_signal(41), B2
                           => n144, ZN => n258);
   U87 : NAND2_X1 port map( A1 => n230, A2 => n229, ZN => Y(29));
   U88 : AOI22_X1 port map( A1 => A_neg(29), A2 => n152, B1 => A_signal(29), B2
                           => n143, ZN => n230);
   U89 : AOI222_X1 port map( A1 => A_shifted(29), A2 => n178, B1 => 
                           zeroSignal(29), B2 => n169, C1 => A_neg_shifted(29),
                           C2 => n163, ZN => n229);
   U90 : NAND2_X1 port map( A1 => n266, A2 => n265, ZN => Y(45));
   U91 : AOI222_X1 port map( A1 => A_shifted(45), A2 => n180, B1 => 
                           zeroSignal(45), B2 => n171, C1 => A_neg_shifted(45),
                           C2 => n162, ZN => n265);
   U92 : AOI22_X1 port map( A1 => A_neg(45), A2 => n154, B1 => A_signal(45), B2
                           => n145, ZN => n266);
   U93 : NAND2_X1 port map( A1 => n262, A2 => n261, ZN => Y(43));
   U94 : AOI222_X1 port map( A1 => A_shifted(43), A2 => n180, B1 => 
                           zeroSignal(43), B2 => n171, C1 => A_neg_shifted(43),
                           C2 => n162, ZN => n261);
   U95 : AOI22_X1 port map( A1 => A_neg(43), A2 => n154, B1 => A_signal(43), B2
                           => n145, ZN => n262);
   U96 : NAND2_X1 port map( A1 => n250, A2 => n249, ZN => Y(38));
   U97 : AOI22_X1 port map( A1 => A_neg(38), A2 => n153, B1 => A_signal(38), B2
                           => n144, ZN => n250);
   U98 : AOI222_X1 port map( A1 => A_shifted(38), A2 => n179, B1 => 
                           zeroSignal(38), B2 => n170, C1 => A_neg_shifted(38),
                           C2 => n162, ZN => n249);
   U99 : NAND2_X1 port map( A1 => n264, A2 => n263, ZN => Y(44));
   U100 : AOI222_X1 port map( A1 => A_shifted(44), A2 => n180, B1 => 
                           zeroSignal(44), B2 => n171, C1 => A_neg_shifted(44),
                           C2 => n162, ZN => n263);
   U101 : AOI22_X1 port map( A1 => A_neg(44), A2 => n154, B1 => A_signal(44), 
                           B2 => n145, ZN => n264);
   U102 : NAND2_X1 port map( A1 => n268, A2 => n267, ZN => Y(46));
   U103 : AOI222_X1 port map( A1 => A_shifted(46), A2 => n180, B1 => 
                           zeroSignal(46), B2 => n171, C1 => A_neg_shifted(46),
                           C2 => n161, ZN => n267);
   U104 : AOI22_X1 port map( A1 => A_neg(46), A2 => n154, B1 => A_signal(46), 
                           B2 => n145, ZN => n268);
   U105 : NAND2_X1 port map( A1 => n270, A2 => n269, ZN => Y(47));
   U106 : AOI222_X1 port map( A1 => A_shifted(47), A2 => n180, B1 => 
                           zeroSignal(47), B2 => n171, C1 => A_neg_shifted(47),
                           C2 => n161, ZN => n269);
   U107 : AOI22_X1 port map( A1 => A_neg(47), A2 => n154, B1 => A_signal(47), 
                           B2 => n145, ZN => n270);
   U108 : NAND2_X1 port map( A1 => n274, A2 => n273, ZN => Y(49));
   U109 : AOI222_X1 port map( A1 => A_shifted(49), A2 => n180, B1 => 
                           zeroSignal(49), B2 => n171, C1 => A_neg_shifted(49),
                           C2 => n161, ZN => n273);
   U110 : AOI22_X1 port map( A1 => A_neg(49), A2 => n154, B1 => A_signal(49), 
                           B2 => n145, ZN => n274);
   U111 : NAND2_X1 port map( A1 => n260, A2 => n259, ZN => Y(42));
   U112 : AOI22_X1 port map( A1 => A_neg(42), A2 => n154, B1 => A_signal(42), 
                           B2 => n145, ZN => n260);
   U113 : AOI222_X1 port map( A1 => A_shifted(42), A2 => n180, B1 => 
                           zeroSignal(42), B2 => n171, C1 => A_neg_shifted(42),
                           C2 => n162, ZN => n259);
   U114 : NAND2_X1 port map( A1 => n280, A2 => n279, ZN => Y(51));
   U115 : AOI222_X1 port map( A1 => A_shifted(51), A2 => n180, B1 => 
                           zeroSignal(51), B2 => n171, C1 => A_neg_shifted(51),
                           C2 => n161, ZN => n279);
   U116 : AOI22_X1 port map( A1 => A_neg(51), A2 => n154, B1 => A_signal(51), 
                           B2 => n145, ZN => n280);
   U117 : NAND2_X1 port map( A1 => n282, A2 => n281, ZN => Y(52));
   U118 : AOI222_X1 port map( A1 => A_shifted(52), A2 => n180, B1 => 
                           zeroSignal(52), B2 => n171, C1 => A_neg_shifted(52),
                           C2 => n161, ZN => n281);
   U119 : AOI22_X1 port map( A1 => A_neg(52), A2 => n154, B1 => A_signal(52), 
                           B2 => n145, ZN => n282);
   U120 : NAND2_X1 port map( A1 => n278, A2 => n277, ZN => Y(50));
   U121 : AOI222_X1 port map( A1 => A_shifted(50), A2 => n180, B1 => 
                           zeroSignal(50), B2 => n171, C1 => A_neg_shifted(50),
                           C2 => n161, ZN => n277);
   U122 : AOI22_X1 port map( A1 => A_neg(50), A2 => n154, B1 => A_signal(50), 
                           B2 => n145, ZN => n278);
   U123 : NAND2_X1 port map( A1 => n292, A2 => n291, ZN => Y(57));
   U124 : AOI222_X1 port map( A1 => A_shifted(57), A2 => n181, B1 => 
                           zeroSignal(57), B2 => n172, C1 => A_neg_shifted(57),
                           C2 => n160, ZN => n291);
   U125 : AOI22_X1 port map( A1 => A_neg(57), A2 => n155, B1 => A_signal(57), 
                           B2 => n146, ZN => n292);
   U126 : NAND2_X1 port map( A1 => n284, A2 => n283, ZN => Y(53));
   U127 : AOI222_X1 port map( A1 => A_shifted(53), A2 => n181, B1 => 
                           zeroSignal(53), B2 => n172, C1 => A_neg_shifted(53),
                           C2 => n161, ZN => n283);
   U128 : AOI22_X1 port map( A1 => A_neg(53), A2 => n155, B1 => A_signal(53), 
                           B2 => n146, ZN => n284);
   U129 : NAND2_X1 port map( A1 => n288, A2 => n287, ZN => Y(55));
   U130 : AOI222_X1 port map( A1 => A_shifted(55), A2 => n181, B1 => 
                           zeroSignal(55), B2 => n172, C1 => A_neg_shifted(55),
                           C2 => n161, ZN => n287);
   U131 : AOI22_X1 port map( A1 => A_neg(55), A2 => n155, B1 => A_signal(55), 
                           B2 => n146, ZN => n288);
   U132 : NAND2_X1 port map( A1 => n236, A2 => n235, ZN => Y(31));
   U133 : AOI222_X1 port map( A1 => A_shifted(31), A2 => n179, B1 => 
                           zeroSignal(31), B2 => n170, C1 => A_neg_shifted(31),
                           C2 => n163, ZN => n235);
   U134 : AOI22_X1 port map( A1 => A_neg(31), A2 => n153, B1 => A_signal(31), 
                           B2 => n144, ZN => n236);
   U135 : NAND2_X1 port map( A1 => n286, A2 => n285, ZN => Y(54));
   U136 : AOI222_X1 port map( A1 => A_shifted(54), A2 => n181, B1 => 
                           zeroSignal(54), B2 => n172, C1 => A_neg_shifted(54),
                           C2 => n161, ZN => n285);
   U137 : AOI22_X1 port map( A1 => A_neg(54), A2 => n155, B1 => A_signal(54), 
                           B2 => n146, ZN => n286);
   U138 : NAND2_X1 port map( A1 => n234, A2 => n233, ZN => Y(30));
   U139 : AOI222_X1 port map( A1 => A_shifted(30), A2 => n178, B1 => 
                           zeroSignal(30), B2 => n169, C1 => A_neg_shifted(30),
                           C2 => n163, ZN => n233);
   U140 : AOI22_X1 port map( A1 => A_neg(30), A2 => n152, B1 => A_signal(30), 
                           B2 => n143, ZN => n234);
   U141 : NAND2_X1 port map( A1 => n272, A2 => n271, ZN => Y(48));
   U142 : AOI22_X1 port map( A1 => A_neg(48), A2 => n154, B1 => A_signal(48), 
                           B2 => n145, ZN => n272);
   U143 : AOI222_X1 port map( A1 => A_shifted(48), A2 => n180, B1 => 
                           zeroSignal(48), B2 => n171, C1 => A_neg_shifted(48),
                           C2 => n161, ZN => n271);
   U144 : NAND2_X1 port map( A1 => n290, A2 => n289, ZN => Y(56));
   U145 : AOI222_X1 port map( A1 => A_shifted(56), A2 => n181, B1 => 
                           zeroSignal(56), B2 => n172, C1 => A_neg_shifted(56),
                           C2 => n161, ZN => n289);
   U146 : AOI22_X1 port map( A1 => A_neg(56), A2 => n155, B1 => A_signal(56), 
                           B2 => n146, ZN => n290);
   U147 : NAND2_X1 port map( A1 => n238, A2 => n237, ZN => Y(32));
   U148 : AOI222_X1 port map( A1 => A_shifted(32), A2 => n179, B1 => 
                           zeroSignal(32), B2 => n170, C1 => A_neg_shifted(32),
                           C2 => n163, ZN => n237);
   U149 : AOI22_X1 port map( A1 => A_neg(32), A2 => n153, B1 => A_signal(32), 
                           B2 => n144, ZN => n238);
   U150 : NAND2_X1 port map( A1 => n240, A2 => n239, ZN => Y(33));
   U151 : AOI222_X1 port map( A1 => A_shifted(33), A2 => n179, B1 => 
                           zeroSignal(33), B2 => n170, C1 => A_neg_shifted(33),
                           C2 => n163, ZN => n239);
   U152 : AOI22_X1 port map( A1 => A_neg(33), A2 => n153, B1 => A_signal(33), 
                           B2 => n144, ZN => n240);
   U153 : NAND2_X1 port map( A1 => n294, A2 => n293, ZN => Y(58));
   U154 : AOI222_X1 port map( A1 => A_shifted(58), A2 => n181, B1 => 
                           zeroSignal(58), B2 => n172, C1 => A_neg_shifted(58),
                           C2 => n160, ZN => n293);
   U155 : AOI22_X1 port map( A1 => A_neg(58), A2 => n155, B1 => A_signal(58), 
                           B2 => n146, ZN => n294);
   U156 : NAND2_X1 port map( A1 => n296, A2 => n295, ZN => Y(59));
   U157 : AOI222_X1 port map( A1 => A_shifted(59), A2 => n181, B1 => 
                           zeroSignal(59), B2 => n172, C1 => A_neg_shifted(59),
                           C2 => n160, ZN => n295);
   U158 : AOI22_X1 port map( A1 => A_neg(59), A2 => n155, B1 => A_signal(59), 
                           B2 => n146, ZN => n296);
   U159 : NAND2_X1 port map( A1 => n300, A2 => n299, ZN => Y(60));
   U160 : AOI222_X1 port map( A1 => A_shifted(60), A2 => n181, B1 => 
                           zeroSignal(60), B2 => n172, C1 => A_neg_shifted(60),
                           C2 => n160, ZN => n299);
   U161 : AOI22_X1 port map( A1 => A_neg(60), A2 => n155, B1 => A_signal(60), 
                           B2 => n146, ZN => n300);
   U162 : NAND2_X1 port map( A1 => n302, A2 => n301, ZN => Y(61));
   U163 : AOI22_X1 port map( A1 => A_neg(61), A2 => n155, B1 => A_signal(61), 
                           B2 => n146, ZN => n302);
   U164 : AOI222_X1 port map( A1 => A_shifted(61), A2 => n181, B1 => 
                           zeroSignal(61), B2 => n172, C1 => A_neg_shifted(61),
                           C2 => n160, ZN => n301);
   U165 : NAND2_X1 port map( A1 => n306, A2 => n305, ZN => Y(63));
   U166 : AOI222_X1 port map( A1 => A_shifted(63), A2 => n181, B1 => 
                           zeroSignal(63), B2 => n172, C1 => A_neg_shifted(63),
                           C2 => n160, ZN => n305);
   U167 : AOI22_X1 port map( A1 => A_neg(63), A2 => n155, B1 => A_signal(63), 
                           B2 => n146, ZN => n306);
   U168 : NAND2_X1 port map( A1 => n304, A2 => n303, ZN => Y(62));
   U169 : AOI222_X1 port map( A1 => A_shifted(62), A2 => n181, B1 => 
                           zeroSignal(62), B2 => n172, C1 => A_neg_shifted(62),
                           C2 => n160, ZN => n303);
   U170 : AOI22_X1 port map( A1 => A_neg(62), A2 => n155, B1 => A_signal(62), 
                           B2 => n146, ZN => n304);
   U171 : NAND2_X1 port map( A1 => n188, A2 => n187, ZN => Y(0));
   U172 : AOI22_X1 port map( A1 => A_neg(0), A2 => n151, B1 => A_signal(0), B2 
                           => n142, ZN => n188);
   U173 : AOI222_X1 port map( A1 => A_shifted(0), A2 => n177, B1 => 
                           zeroSignal(0), B2 => n168, C1 => A_neg_shifted(0), 
                           C2 => n165, ZN => n187);
   U174 : NAND2_X1 port map( A1 => n210, A2 => n209, ZN => Y(1));
   U175 : AOI22_X1 port map( A1 => A_neg(1), A2 => n151, B1 => A_signal(1), B2 
                           => n142, ZN => n210);
   U176 : AOI222_X1 port map( A1 => A_shifted(1), A2 => n177, B1 => 
                           zeroSignal(1), B2 => n168, C1 => A_neg_shifted(1), 
                           C2 => n164, ZN => n209);
   U177 : NAND2_X1 port map( A1 => n232, A2 => n231, ZN => Y(2));
   U178 : AOI22_X1 port map( A1 => A_neg(2), A2 => n152, B1 => A_signal(2), B2 
                           => n143, ZN => n232);
   U179 : AOI222_X1 port map( A1 => A_shifted(2), A2 => n178, B1 => 
                           zeroSignal(2), B2 => n169, C1 => A_neg_shifted(2), 
                           C2 => n163, ZN => n231);
   U180 : NAND2_X1 port map( A1 => n254, A2 => n253, ZN => Y(3));
   U181 : AOI22_X1 port map( A1 => A_neg(3), A2 => n153, B1 => A_signal(3), B2 
                           => n144, ZN => n254);
   U182 : AOI222_X1 port map( A1 => A_shifted(3), A2 => n179, B1 => 
                           zeroSignal(3), B2 => n170, C1 => A_neg_shifted(3), 
                           C2 => n162, ZN => n253);
   U183 : NAND2_X1 port map( A1 => n276, A2 => n275, ZN => Y(4));
   U184 : AOI22_X1 port map( A1 => A_neg(4), A2 => n154, B1 => A_signal(4), B2 
                           => n145, ZN => n276);
   U185 : AOI222_X1 port map( A1 => A_shifted(4), A2 => n180, B1 => 
                           zeroSignal(4), B2 => n171, C1 => A_neg_shifted(4), 
                           C2 => n161, ZN => n275);
   U186 : NAND2_X1 port map( A1 => n298, A2 => n297, ZN => Y(5));
   U187 : AOI22_X1 port map( A1 => A_neg(5), A2 => n155, B1 => A_signal(5), B2 
                           => n146, ZN => n298);
   U188 : AOI222_X1 port map( A1 => A_shifted(5), A2 => n181, B1 => 
                           zeroSignal(5), B2 => n172, C1 => A_neg_shifted(5), 
                           C2 => n160, ZN => n297);
   U189 : NAND2_X1 port map( A1 => n308, A2 => n307, ZN => Y(6));
   U190 : AOI22_X1 port map( A1 => A_neg(6), A2 => n156, B1 => A_signal(6), B2 
                           => n147, ZN => n308);
   U191 : AOI222_X1 port map( A1 => A_shifted(6), A2 => n182, B1 => 
                           zeroSignal(6), B2 => n173, C1 => A_neg_shifted(6), 
                           C2 => n160, ZN => n307);
   U192 : NAND2_X1 port map( A1 => n310, A2 => n309, ZN => Y(7));
   U193 : AOI22_X1 port map( A1 => A_neg(7), A2 => n156, B1 => A_signal(7), B2 
                           => n147, ZN => n310);
   U194 : AOI222_X1 port map( A1 => A_shifted(7), A2 => n182, B1 => 
                           zeroSignal(7), B2 => n173, C1 => A_neg_shifted(7), 
                           C2 => n160, ZN => n309);
   U195 : NAND2_X1 port map( A1 => n312, A2 => n311, ZN => Y(8));
   U196 : AOI22_X1 port map( A1 => A_neg(8), A2 => n156, B1 => A_signal(8), B2 
                           => n147, ZN => n312);
   U197 : AOI222_X1 port map( A1 => A_shifted(8), A2 => n182, B1 => 
                           zeroSignal(8), B2 => n173, C1 => A_neg_shifted(8), 
                           C2 => n160, ZN => n311);
   U198 : NAND2_X1 port map( A1 => n318, A2 => n317, ZN => Y(9));
   U199 : AOI22_X1 port map( A1 => A_neg(9), A2 => n156, B1 => A_signal(9), B2 
                           => n147, ZN => n318);
   U200 : AOI222_X1 port map( A1 => A_shifted(9), A2 => n182, B1 => 
                           zeroSignal(9), B2 => n173, C1 => A_neg_shifted(9), 
                           C2 => n160, ZN => n317);
   U201 : NAND2_X1 port map( A1 => n190, A2 => n189, ZN => Y(10));
   U202 : AOI22_X1 port map( A1 => A_neg(10), A2 => n151, B1 => A_signal(10), 
                           B2 => n142, ZN => n190);
   U203 : AOI222_X1 port map( A1 => A_shifted(10), A2 => n177, B1 => 
                           zeroSignal(10), B2 => n168, C1 => A_neg_shifted(10),
                           C2 => n165, ZN => n189);
   U204 : NAND2_X1 port map( A1 => n192, A2 => n191, ZN => Y(11));
   U205 : AOI22_X1 port map( A1 => A_neg(11), A2 => n151, B1 => A_signal(11), 
                           B2 => n142, ZN => n192);
   U206 : AOI222_X1 port map( A1 => A_shifted(11), A2 => n177, B1 => 
                           zeroSignal(11), B2 => n168, C1 => A_neg_shifted(11),
                           C2 => n165, ZN => n191);
   U207 : NAND2_X1 port map( A1 => n194, A2 => n193, ZN => Y(12));
   U208 : AOI22_X1 port map( A1 => A_neg(12), A2 => n151, B1 => A_signal(12), 
                           B2 => n142, ZN => n194);
   U209 : AOI222_X1 port map( A1 => A_shifted(12), A2 => n177, B1 => 
                           zeroSignal(12), B2 => n168, C1 => A_neg_shifted(12),
                           C2 => n165, ZN => n193);
   U210 : NAND2_X1 port map( A1 => n196, A2 => n195, ZN => Y(13));
   U211 : AOI22_X1 port map( A1 => A_neg(13), A2 => n151, B1 => A_signal(13), 
                           B2 => n142, ZN => n196);
   U212 : AOI222_X1 port map( A1 => A_shifted(13), A2 => n177, B1 => 
                           zeroSignal(13), B2 => n168, C1 => A_neg_shifted(13),
                           C2 => n164, ZN => n195);
   U213 : NAND2_X1 port map( A1 => n198, A2 => n197, ZN => Y(14));
   U214 : AOI22_X1 port map( A1 => A_neg(14), A2 => n151, B1 => A_signal(14), 
                           B2 => n142, ZN => n198);
   U215 : AOI222_X1 port map( A1 => A_shifted(14), A2 => n177, B1 => 
                           zeroSignal(14), B2 => n168, C1 => A_neg_shifted(14),
                           C2 => n164, ZN => n197);
   U216 : NAND2_X1 port map( A1 => n200, A2 => n199, ZN => Y(15));
   U217 : AOI22_X1 port map( A1 => A_neg(15), A2 => n151, B1 => A_signal(15), 
                           B2 => n142, ZN => n200);
   U218 : AOI222_X1 port map( A1 => A_shifted(15), A2 => n177, B1 => 
                           zeroSignal(15), B2 => n168, C1 => A_neg_shifted(15),
                           C2 => n164, ZN => n199);
   U219 : NAND2_X1 port map( A1 => n202, A2 => n201, ZN => Y(16));
   U220 : AOI22_X1 port map( A1 => A_neg(16), A2 => n151, B1 => A_signal(16), 
                           B2 => n142, ZN => n202);
   U221 : AOI222_X1 port map( A1 => A_shifted(16), A2 => n177, B1 => 
                           zeroSignal(16), B2 => n168, C1 => A_neg_shifted(16),
                           C2 => n164, ZN => n201);
   U222 : NAND2_X1 port map( A1 => n204, A2 => n203, ZN => Y(17));
   U223 : AOI22_X1 port map( A1 => A_neg(17), A2 => n151, B1 => A_signal(17), 
                           B2 => n142, ZN => n204);
   U224 : AOI222_X1 port map( A1 => A_shifted(17), A2 => n177, B1 => 
                           zeroSignal(17), B2 => n168, C1 => A_neg_shifted(17),
                           C2 => n164, ZN => n203);
   U225 : NAND2_X1 port map( A1 => n206, A2 => n205, ZN => Y(18));
   U226 : AOI22_X1 port map( A1 => A_neg(18), A2 => n151, B1 => A_signal(18), 
                           B2 => n142, ZN => n206);
   U227 : AOI222_X1 port map( A1 => A_shifted(18), A2 => n177, B1 => 
                           zeroSignal(18), B2 => n168, C1 => A_neg_shifted(18),
                           C2 => n164, ZN => n205);
   U228 : NAND2_X1 port map( A1 => n208, A2 => n207, ZN => Y(19));
   U229 : AOI22_X1 port map( A1 => A_neg(19), A2 => n151, B1 => A_signal(19), 
                           B2 => n142, ZN => n208);
   U230 : AOI222_X1 port map( A1 => A_shifted(19), A2 => n177, B1 => 
                           zeroSignal(19), B2 => n168, C1 => A_neg_shifted(19),
                           C2 => n164, ZN => n207);
   U231 : NAND2_X1 port map( A1 => n212, A2 => n211, ZN => Y(20));
   U232 : AOI22_X1 port map( A1 => A_neg(20), A2 => n152, B1 => A_signal(20), 
                           B2 => n143, ZN => n212);
   U233 : AOI222_X1 port map( A1 => A_shifted(20), A2 => n178, B1 => 
                           zeroSignal(20), B2 => n169, C1 => A_neg_shifted(20),
                           C2 => n164, ZN => n211);
   U234 : NAND2_X1 port map( A1 => n214, A2 => n213, ZN => Y(21));
   U235 : AOI22_X1 port map( A1 => A_neg(21), A2 => n152, B1 => A_signal(21), 
                           B2 => n143, ZN => n214);
   U236 : AOI222_X1 port map( A1 => A_shifted(21), A2 => n178, B1 => 
                           zeroSignal(21), B2 => n169, C1 => A_neg_shifted(21),
                           C2 => n164, ZN => n213);
   U237 : NAND2_X1 port map( A1 => n216, A2 => n215, ZN => Y(22));
   U238 : AOI22_X1 port map( A1 => A_neg(22), A2 => n152, B1 => A_signal(22), 
                           B2 => n143, ZN => n216);
   U239 : AOI222_X1 port map( A1 => A_shifted(22), A2 => n178, B1 => 
                           zeroSignal(22), B2 => n169, C1 => A_neg_shifted(22),
                           C2 => n164, ZN => n215);
   U240 : NAND2_X1 port map( A1 => n218, A2 => n217, ZN => Y(23));
   U241 : AOI22_X1 port map( A1 => A_neg(23), A2 => n152, B1 => A_signal(23), 
                           B2 => n143, ZN => n218);
   U242 : AOI222_X1 port map( A1 => A_shifted(23), A2 => n178, B1 => 
                           zeroSignal(23), B2 => n169, C1 => A_neg_shifted(23),
                           C2 => n164, ZN => n217);
   U243 : AOI222_X1 port map( A1 => A_shifted(25), A2 => n178, B1 => 
                           zeroSignal(25), B2 => n169, C1 => A_neg_shifted(25),
                           C2 => n163, ZN => n221);
   U244 : AOI22_X1 port map( A1 => A_neg(24), A2 => n152, B1 => A_signal(24), 
                           B2 => n143, ZN => n220);

end SYN_BEHAVIORAL_2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity MUX51_MuxNbit64_19 is

   port( zeroSignal, A_signal, A_neg, A_shifted, A_neg_shifted : in 
         std_logic_vector (63 downto 0);  Sel : in std_logic_vector (2 downto 
         0);  Y : out std_logic_vector (63 downto 0));

end MUX51_MuxNbit64_19;

architecture SYN_BEHAVIORAL_2 of MUX51_MuxNbit64_19 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, 
      n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, 
      n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, 
      n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, 
      n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, 
      n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, 
      n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, 
      n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, 
      n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, 
      n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, 
      n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, 
      n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, 
      n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, 
      n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, 
      n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, 
      n320 : std_logic;

begin
   
   U1 : AND3_X1 port map( A1 => n319, A2 => n320, A3 => Sel(2), ZN => n141);
   U2 : BUF_X1 port map( A => n141, Z => n166);
   U3 : BUF_X1 port map( A => n185, Z => n184);
   U4 : BUF_X1 port map( A => n159, Z => n158);
   U5 : BUF_X1 port map( A => n150, Z => n149);
   U6 : BUF_X1 port map( A => n141, Z => n167);
   U7 : BUF_X1 port map( A => n185, Z => n183);
   U8 : BUF_X1 port map( A => n159, Z => n157);
   U9 : BUF_X1 port map( A => n150, Z => n148);
   U10 : BUF_X1 port map( A => n176, Z => n175);
   U11 : BUF_X1 port map( A => n176, Z => n174);
   U12 : BUF_X1 port map( A => n158, Z => n152);
   U13 : BUF_X1 port map( A => n184, Z => n178);
   U14 : BUF_X1 port map( A => n149, Z => n143);
   U15 : BUF_X1 port map( A => n166, Z => n163);
   U16 : BUF_X1 port map( A => n184, Z => n179);
   U17 : BUF_X1 port map( A => n158, Z => n153);
   U18 : BUF_X1 port map( A => n149, Z => n144);
   U19 : BUF_X1 port map( A => n167, Z => n162);
   U20 : BUF_X1 port map( A => n183, Z => n180);
   U21 : BUF_X1 port map( A => n157, Z => n154);
   U22 : BUF_X1 port map( A => n148, Z => n145);
   U23 : BUF_X1 port map( A => n167, Z => n161);
   U24 : BUF_X1 port map( A => n183, Z => n181);
   U25 : BUF_X1 port map( A => n157, Z => n155);
   U26 : BUF_X1 port map( A => n148, Z => n146);
   U27 : BUF_X1 port map( A => n167, Z => n160);
   U28 : BUF_X1 port map( A => n158, Z => n151);
   U29 : BUF_X1 port map( A => n149, Z => n142);
   U30 : BUF_X1 port map( A => n175, Z => n168);
   U31 : BUF_X1 port map( A => n175, Z => n170);
   U32 : BUF_X1 port map( A => n174, Z => n171);
   U33 : BUF_X1 port map( A => n174, Z => n172);
   U34 : BUF_X1 port map( A => n166, Z => n164);
   U35 : BUF_X1 port map( A => n175, Z => n169);
   U36 : BUF_X1 port map( A => n184, Z => n177);
   U37 : BUF_X1 port map( A => n166, Z => n165);
   U38 : BUF_X1 port map( A => n157, Z => n156);
   U39 : BUF_X1 port map( A => n148, Z => n147);
   U40 : BUF_X1 port map( A => n174, Z => n173);
   U41 : BUF_X1 port map( A => n183, Z => n182);
   U42 : INV_X1 port map( A => Sel(1), ZN => n320);
   U43 : BUF_X1 port map( A => n314, Z => n159);
   U44 : NOR3_X1 port map( A1 => Sel(0), A2 => Sel(2), A3 => n320, ZN => n314);
   U45 : BUF_X1 port map( A => n316, Z => n185);
   U46 : NOR3_X1 port map( A1 => n319, A2 => Sel(2), A3 => n320, ZN => n316);
   U47 : INV_X1 port map( A => Sel(0), ZN => n319);
   U48 : BUF_X1 port map( A => n313, Z => n150);
   U49 : NOR3_X1 port map( A1 => Sel(1), A2 => Sel(2), A3 => n319, ZN => n313);
   U50 : BUF_X1 port map( A => n315, Z => n176);
   U51 : NOR2_X1 port map( A1 => n165, A2 => n186, ZN => n315);
   U52 : AOI21_X1 port map( B1 => n319, B2 => n320, A => Sel(2), ZN => n186);
   U53 : NAND2_X1 port map( A1 => n226, A2 => n225, ZN => Y(27));
   U54 : AOI22_X1 port map( A1 => A_neg(27), A2 => n152, B1 => A_signal(27), B2
                           => n143, ZN => n226);
   U55 : NAND2_X1 port map( A1 => n224, A2 => n223, ZN => Y(26));
   U56 : AOI222_X1 port map( A1 => A_shifted(26), A2 => n178, B1 => 
                           zeroSignal(26), B2 => n169, C1 => A_neg_shifted(26),
                           C2 => n163, ZN => n223);
   U57 : NAND2_X1 port map( A1 => n228, A2 => n227, ZN => Y(28));
   U58 : AOI22_X1 port map( A1 => A_neg(28), A2 => n152, B1 => A_signal(28), B2
                           => n143, ZN => n228);
   U59 : AOI222_X1 port map( A1 => A_shifted(28), A2 => n178, B1 => 
                           zeroSignal(28), B2 => n169, C1 => A_neg_shifted(28),
                           C2 => n163, ZN => n227);
   U60 : NAND2_X1 port map( A1 => n230, A2 => n229, ZN => Y(29));
   U61 : AOI22_X1 port map( A1 => A_neg(29), A2 => n152, B1 => A_signal(29), B2
                           => n143, ZN => n230);
   U62 : AOI222_X1 port map( A1 => A_shifted(29), A2 => n178, B1 => 
                           zeroSignal(29), B2 => n169, C1 => A_neg_shifted(29),
                           C2 => n163, ZN => n229);
   U63 : NAND2_X1 port map( A1 => n234, A2 => n233, ZN => Y(30));
   U64 : AOI22_X1 port map( A1 => A_neg(30), A2 => n152, B1 => A_signal(30), B2
                           => n143, ZN => n234);
   U65 : AOI222_X1 port map( A1 => A_shifted(30), A2 => n178, B1 => 
                           zeroSignal(30), B2 => n169, C1 => A_neg_shifted(30),
                           C2 => n163, ZN => n233);
   U66 : NAND2_X1 port map( A1 => n248, A2 => n247, ZN => Y(37));
   U67 : AOI222_X1 port map( A1 => A_shifted(37), A2 => n179, B1 => 
                           zeroSignal(37), B2 => n170, C1 => A_neg_shifted(37),
                           C2 => n162, ZN => n247);
   U68 : AOI22_X1 port map( A1 => A_neg(37), A2 => n153, B1 => A_signal(37), B2
                           => n144, ZN => n248);
   U69 : NAND2_X1 port map( A1 => n246, A2 => n245, ZN => Y(36));
   U70 : AOI222_X1 port map( A1 => A_shifted(36), A2 => n179, B1 => 
                           zeroSignal(36), B2 => n170, C1 => A_neg_shifted(36),
                           C2 => n162, ZN => n245);
   U71 : AOI22_X1 port map( A1 => A_neg(36), A2 => n153, B1 => A_signal(36), B2
                           => n144, ZN => n246);
   U72 : NAND2_X1 port map( A1 => n250, A2 => n249, ZN => Y(38));
   U73 : AOI222_X1 port map( A1 => A_shifted(38), A2 => n179, B1 => 
                           zeroSignal(38), B2 => n170, C1 => A_neg_shifted(38),
                           C2 => n162, ZN => n249);
   U74 : AOI22_X1 port map( A1 => A_neg(38), A2 => n153, B1 => A_signal(38), B2
                           => n144, ZN => n250);
   U75 : NAND2_X1 port map( A1 => n252, A2 => n251, ZN => Y(39));
   U76 : AOI222_X1 port map( A1 => A_shifted(39), A2 => n179, B1 => 
                           zeroSignal(39), B2 => n170, C1 => A_neg_shifted(39),
                           C2 => n162, ZN => n251);
   U77 : AOI22_X1 port map( A1 => A_neg(39), A2 => n153, B1 => A_signal(39), B2
                           => n144, ZN => n252);
   U78 : NAND2_X1 port map( A1 => n258, A2 => n257, ZN => Y(41));
   U79 : AOI222_X1 port map( A1 => A_shifted(41), A2 => n179, B1 => 
                           zeroSignal(41), B2 => n170, C1 => A_neg_shifted(41),
                           C2 => n162, ZN => n257);
   U80 : AOI22_X1 port map( A1 => A_neg(41), A2 => n153, B1 => A_signal(41), B2
                           => n144, ZN => n258);
   U81 : NAND2_X1 port map( A1 => n260, A2 => n259, ZN => Y(42));
   U82 : AOI222_X1 port map( A1 => A_shifted(42), A2 => n180, B1 => 
                           zeroSignal(42), B2 => n171, C1 => A_neg_shifted(42),
                           C2 => n162, ZN => n259);
   U83 : AOI22_X1 port map( A1 => A_neg(42), A2 => n154, B1 => A_signal(42), B2
                           => n145, ZN => n260);
   U84 : NAND2_X1 port map( A1 => n236, A2 => n235, ZN => Y(31));
   U85 : AOI22_X1 port map( A1 => A_neg(31), A2 => n153, B1 => A_signal(31), B2
                           => n144, ZN => n236);
   U86 : AOI222_X1 port map( A1 => A_shifted(31), A2 => n179, B1 => 
                           zeroSignal(31), B2 => n170, C1 => A_neg_shifted(31),
                           C2 => n163, ZN => n235);
   U87 : NAND2_X1 port map( A1 => n262, A2 => n261, ZN => Y(43));
   U88 : AOI222_X1 port map( A1 => A_shifted(43), A2 => n180, B1 => 
                           zeroSignal(43), B2 => n171, C1 => A_neg_shifted(43),
                           C2 => n162, ZN => n261);
   U89 : AOI22_X1 port map( A1 => A_neg(43), A2 => n154, B1 => A_signal(43), B2
                           => n145, ZN => n262);
   U90 : NAND2_X1 port map( A1 => n256, A2 => n255, ZN => Y(40));
   U91 : AOI22_X1 port map( A1 => A_neg(40), A2 => n153, B1 => A_signal(40), B2
                           => n144, ZN => n256);
   U92 : AOI222_X1 port map( A1 => A_shifted(40), A2 => n179, B1 => 
                           zeroSignal(40), B2 => n170, C1 => A_neg_shifted(40),
                           C2 => n162, ZN => n255);
   U93 : NAND2_X1 port map( A1 => n266, A2 => n265, ZN => Y(45));
   U94 : AOI222_X1 port map( A1 => A_shifted(45), A2 => n180, B1 => 
                           zeroSignal(45), B2 => n171, C1 => A_neg_shifted(45),
                           C2 => n162, ZN => n265);
   U95 : AOI22_X1 port map( A1 => A_neg(45), A2 => n154, B1 => A_signal(45), B2
                           => n145, ZN => n266);
   U96 : NAND2_X1 port map( A1 => n270, A2 => n269, ZN => Y(47));
   U97 : AOI222_X1 port map( A1 => A_shifted(47), A2 => n180, B1 => 
                           zeroSignal(47), B2 => n171, C1 => A_neg_shifted(47),
                           C2 => n161, ZN => n269);
   U98 : AOI22_X1 port map( A1 => A_neg(47), A2 => n154, B1 => A_signal(47), B2
                           => n145, ZN => n270);
   U99 : NAND2_X1 port map( A1 => n268, A2 => n267, ZN => Y(46));
   U100 : AOI222_X1 port map( A1 => A_shifted(46), A2 => n180, B1 => 
                           zeroSignal(46), B2 => n171, C1 => A_neg_shifted(46),
                           C2 => n161, ZN => n267);
   U101 : AOI22_X1 port map( A1 => A_neg(46), A2 => n154, B1 => A_signal(46), 
                           B2 => n145, ZN => n268);
   U102 : NAND2_X1 port map( A1 => n272, A2 => n271, ZN => Y(48));
   U103 : AOI222_X1 port map( A1 => A_shifted(48), A2 => n180, B1 => 
                           zeroSignal(48), B2 => n171, C1 => A_neg_shifted(48),
                           C2 => n161, ZN => n271);
   U104 : AOI22_X1 port map( A1 => A_neg(48), A2 => n154, B1 => A_signal(48), 
                           B2 => n145, ZN => n272);
   U105 : NAND2_X1 port map( A1 => n274, A2 => n273, ZN => Y(49));
   U106 : AOI222_X1 port map( A1 => A_shifted(49), A2 => n180, B1 => 
                           zeroSignal(49), B2 => n171, C1 => A_neg_shifted(49),
                           C2 => n161, ZN => n273);
   U107 : AOI22_X1 port map( A1 => A_neg(49), A2 => n154, B1 => A_signal(49), 
                           B2 => n145, ZN => n274);
   U108 : NAND2_X1 port map( A1 => n282, A2 => n281, ZN => Y(52));
   U109 : AOI222_X1 port map( A1 => A_shifted(52), A2 => n180, B1 => 
                           zeroSignal(52), B2 => n171, C1 => A_neg_shifted(52),
                           C2 => n161, ZN => n281);
   U110 : AOI22_X1 port map( A1 => A_neg(52), A2 => n154, B1 => A_signal(52), 
                           B2 => n145, ZN => n282);
   U111 : NAND2_X1 port map( A1 => n264, A2 => n263, ZN => Y(44));
   U112 : AOI22_X1 port map( A1 => A_neg(44), A2 => n154, B1 => A_signal(44), 
                           B2 => n145, ZN => n264);
   U113 : AOI222_X1 port map( A1 => A_shifted(44), A2 => n180, B1 => 
                           zeroSignal(44), B2 => n171, C1 => A_neg_shifted(44),
                           C2 => n162, ZN => n263);
   U114 : NAND2_X1 port map( A1 => n280, A2 => n279, ZN => Y(51));
   U115 : AOI222_X1 port map( A1 => A_shifted(51), A2 => n180, B1 => 
                           zeroSignal(51), B2 => n171, C1 => A_neg_shifted(51),
                           C2 => n161, ZN => n279);
   U116 : AOI22_X1 port map( A1 => A_neg(51), A2 => n154, B1 => A_signal(51), 
                           B2 => n145, ZN => n280);
   U117 : NAND2_X1 port map( A1 => n284, A2 => n283, ZN => Y(53));
   U118 : AOI222_X1 port map( A1 => A_shifted(53), A2 => n181, B1 => 
                           zeroSignal(53), B2 => n172, C1 => A_neg_shifted(53),
                           C2 => n161, ZN => n283);
   U119 : AOI22_X1 port map( A1 => A_neg(53), A2 => n155, B1 => A_signal(53), 
                           B2 => n146, ZN => n284);
   U120 : NAND2_X1 port map( A1 => n296, A2 => n295, ZN => Y(59));
   U121 : AOI222_X1 port map( A1 => A_shifted(59), A2 => n181, B1 => 
                           zeroSignal(59), B2 => n172, C1 => A_neg_shifted(59),
                           C2 => n160, ZN => n295);
   U122 : AOI22_X1 port map( A1 => A_neg(59), A2 => n155, B1 => A_signal(59), 
                           B2 => n146, ZN => n296);
   U123 : NAND2_X1 port map( A1 => n286, A2 => n285, ZN => Y(54));
   U124 : AOI222_X1 port map( A1 => A_shifted(54), A2 => n181, B1 => 
                           zeroSignal(54), B2 => n172, C1 => A_neg_shifted(54),
                           C2 => n161, ZN => n285);
   U125 : AOI22_X1 port map( A1 => A_neg(54), A2 => n155, B1 => A_signal(54), 
                           B2 => n146, ZN => n286);
   U126 : NAND2_X1 port map( A1 => n288, A2 => n287, ZN => Y(55));
   U127 : AOI222_X1 port map( A1 => A_shifted(55), A2 => n181, B1 => 
                           zeroSignal(55), B2 => n172, C1 => A_neg_shifted(55),
                           C2 => n161, ZN => n287);
   U128 : AOI22_X1 port map( A1 => A_neg(55), A2 => n155, B1 => A_signal(55), 
                           B2 => n146, ZN => n288);
   U129 : NAND2_X1 port map( A1 => n292, A2 => n291, ZN => Y(57));
   U130 : AOI222_X1 port map( A1 => A_shifted(57), A2 => n181, B1 => 
                           zeroSignal(57), B2 => n172, C1 => A_neg_shifted(57),
                           C2 => n160, ZN => n291);
   U131 : AOI22_X1 port map( A1 => A_neg(57), A2 => n155, B1 => A_signal(57), 
                           B2 => n146, ZN => n292);
   U132 : NAND2_X1 port map( A1 => n278, A2 => n277, ZN => Y(50));
   U133 : AOI22_X1 port map( A1 => A_neg(50), A2 => n154, B1 => A_signal(50), 
                           B2 => n145, ZN => n278);
   U134 : AOI222_X1 port map( A1 => A_shifted(50), A2 => n180, B1 => 
                           zeroSignal(50), B2 => n171, C1 => A_neg_shifted(50),
                           C2 => n161, ZN => n277);
   U135 : NAND2_X1 port map( A1 => n290, A2 => n289, ZN => Y(56));
   U136 : AOI222_X1 port map( A1 => A_shifted(56), A2 => n181, B1 => 
                           zeroSignal(56), B2 => n172, C1 => A_neg_shifted(56),
                           C2 => n161, ZN => n289);
   U137 : AOI22_X1 port map( A1 => A_neg(56), A2 => n155, B1 => A_signal(56), 
                           B2 => n146, ZN => n290);
   U138 : NAND2_X1 port map( A1 => n238, A2 => n237, ZN => Y(32));
   U139 : AOI222_X1 port map( A1 => A_shifted(32), A2 => n179, B1 => 
                           zeroSignal(32), B2 => n170, C1 => A_neg_shifted(32),
                           C2 => n163, ZN => n237);
   U140 : AOI22_X1 port map( A1 => A_neg(32), A2 => n153, B1 => A_signal(32), 
                           B2 => n144, ZN => n238);
   U141 : NAND2_X1 port map( A1 => n294, A2 => n293, ZN => Y(58));
   U142 : AOI222_X1 port map( A1 => A_shifted(58), A2 => n181, B1 => 
                           zeroSignal(58), B2 => n172, C1 => A_neg_shifted(58),
                           C2 => n160, ZN => n293);
   U143 : AOI22_X1 port map( A1 => A_neg(58), A2 => n155, B1 => A_signal(58), 
                           B2 => n146, ZN => n294);
   U144 : NAND2_X1 port map( A1 => n242, A2 => n241, ZN => Y(34));
   U145 : AOI222_X1 port map( A1 => A_shifted(34), A2 => n179, B1 => 
                           zeroSignal(34), B2 => n170, C1 => A_neg_shifted(34),
                           C2 => n163, ZN => n241);
   U146 : AOI22_X1 port map( A1 => A_neg(34), A2 => n153, B1 => A_signal(34), 
                           B2 => n144, ZN => n242);
   U147 : NAND2_X1 port map( A1 => n240, A2 => n239, ZN => Y(33));
   U148 : AOI222_X1 port map( A1 => A_shifted(33), A2 => n179, B1 => 
                           zeroSignal(33), B2 => n170, C1 => A_neg_shifted(33),
                           C2 => n163, ZN => n239);
   U149 : AOI22_X1 port map( A1 => A_neg(33), A2 => n153, B1 => A_signal(33), 
                           B2 => n144, ZN => n240);
   U150 : NAND2_X1 port map( A1 => n244, A2 => n243, ZN => Y(35));
   U151 : AOI222_X1 port map( A1 => A_shifted(35), A2 => n179, B1 => 
                           zeroSignal(35), B2 => n170, C1 => A_neg_shifted(35),
                           C2 => n162, ZN => n243);
   U152 : AOI22_X1 port map( A1 => A_neg(35), A2 => n153, B1 => A_signal(35), 
                           B2 => n144, ZN => n244);
   U153 : NAND2_X1 port map( A1 => n300, A2 => n299, ZN => Y(60));
   U154 : AOI222_X1 port map( A1 => A_shifted(60), A2 => n181, B1 => 
                           zeroSignal(60), B2 => n172, C1 => A_neg_shifted(60),
                           C2 => n160, ZN => n299);
   U155 : AOI22_X1 port map( A1 => A_neg(60), A2 => n155, B1 => A_signal(60), 
                           B2 => n146, ZN => n300);
   U156 : NAND2_X1 port map( A1 => n302, A2 => n301, ZN => Y(61));
   U157 : AOI222_X1 port map( A1 => A_shifted(61), A2 => n181, B1 => 
                           zeroSignal(61), B2 => n172, C1 => A_neg_shifted(61),
                           C2 => n160, ZN => n301);
   U158 : AOI22_X1 port map( A1 => A_neg(61), A2 => n155, B1 => A_signal(61), 
                           B2 => n146, ZN => n302);
   U159 : NAND2_X1 port map( A1 => n304, A2 => n303, ZN => Y(62));
   U160 : AOI222_X1 port map( A1 => A_shifted(62), A2 => n181, B1 => 
                           zeroSignal(62), B2 => n172, C1 => A_neg_shifted(62),
                           C2 => n160, ZN => n303);
   U161 : AOI22_X1 port map( A1 => A_neg(62), A2 => n155, B1 => A_signal(62), 
                           B2 => n146, ZN => n304);
   U162 : NAND2_X1 port map( A1 => n306, A2 => n305, ZN => Y(63));
   U163 : AOI22_X1 port map( A1 => A_neg(63), A2 => n155, B1 => A_signal(63), 
                           B2 => n146, ZN => n306);
   U164 : AOI222_X1 port map( A1 => A_shifted(63), A2 => n181, B1 => 
                           zeroSignal(63), B2 => n172, C1 => A_neg_shifted(63),
                           C2 => n160, ZN => n305);
   U165 : NAND2_X1 port map( A1 => n188, A2 => n187, ZN => Y(0));
   U166 : AOI22_X1 port map( A1 => A_neg(0), A2 => n151, B1 => A_signal(0), B2 
                           => n142, ZN => n188);
   U167 : AOI222_X1 port map( A1 => A_shifted(0), A2 => n177, B1 => 
                           zeroSignal(0), B2 => n168, C1 => A_neg_shifted(0), 
                           C2 => n165, ZN => n187);
   U168 : NAND2_X1 port map( A1 => n210, A2 => n209, ZN => Y(1));
   U169 : AOI22_X1 port map( A1 => A_neg(1), A2 => n151, B1 => A_signal(1), B2 
                           => n142, ZN => n210);
   U170 : AOI222_X1 port map( A1 => A_shifted(1), A2 => n177, B1 => 
                           zeroSignal(1), B2 => n168, C1 => A_neg_shifted(1), 
                           C2 => n164, ZN => n209);
   U171 : NAND2_X1 port map( A1 => n232, A2 => n231, ZN => Y(2));
   U172 : AOI22_X1 port map( A1 => A_neg(2), A2 => n152, B1 => A_signal(2), B2 
                           => n143, ZN => n232);
   U173 : AOI222_X1 port map( A1 => A_shifted(2), A2 => n178, B1 => 
                           zeroSignal(2), B2 => n169, C1 => A_neg_shifted(2), 
                           C2 => n163, ZN => n231);
   U174 : NAND2_X1 port map( A1 => n254, A2 => n253, ZN => Y(3));
   U175 : AOI22_X1 port map( A1 => A_neg(3), A2 => n153, B1 => A_signal(3), B2 
                           => n144, ZN => n254);
   U176 : AOI222_X1 port map( A1 => A_shifted(3), A2 => n179, B1 => 
                           zeroSignal(3), B2 => n170, C1 => A_neg_shifted(3), 
                           C2 => n162, ZN => n253);
   U177 : NAND2_X1 port map( A1 => n276, A2 => n275, ZN => Y(4));
   U178 : AOI22_X1 port map( A1 => A_neg(4), A2 => n154, B1 => A_signal(4), B2 
                           => n145, ZN => n276);
   U179 : AOI222_X1 port map( A1 => A_shifted(4), A2 => n180, B1 => 
                           zeroSignal(4), B2 => n171, C1 => A_neg_shifted(4), 
                           C2 => n161, ZN => n275);
   U180 : NAND2_X1 port map( A1 => n298, A2 => n297, ZN => Y(5));
   U181 : AOI22_X1 port map( A1 => A_neg(5), A2 => n155, B1 => A_signal(5), B2 
                           => n146, ZN => n298);
   U182 : AOI222_X1 port map( A1 => A_shifted(5), A2 => n181, B1 => 
                           zeroSignal(5), B2 => n172, C1 => A_neg_shifted(5), 
                           C2 => n160, ZN => n297);
   U183 : NAND2_X1 port map( A1 => n308, A2 => n307, ZN => Y(6));
   U184 : AOI22_X1 port map( A1 => A_neg(6), A2 => n156, B1 => A_signal(6), B2 
                           => n147, ZN => n308);
   U185 : AOI222_X1 port map( A1 => A_shifted(6), A2 => n182, B1 => 
                           zeroSignal(6), B2 => n173, C1 => A_neg_shifted(6), 
                           C2 => n160, ZN => n307);
   U186 : NAND2_X1 port map( A1 => n310, A2 => n309, ZN => Y(7));
   U187 : AOI22_X1 port map( A1 => A_neg(7), A2 => n156, B1 => A_signal(7), B2 
                           => n147, ZN => n310);
   U188 : AOI222_X1 port map( A1 => A_shifted(7), A2 => n182, B1 => 
                           zeroSignal(7), B2 => n173, C1 => A_neg_shifted(7), 
                           C2 => n160, ZN => n309);
   U189 : NAND2_X1 port map( A1 => n312, A2 => n311, ZN => Y(8));
   U190 : AOI22_X1 port map( A1 => A_neg(8), A2 => n156, B1 => A_signal(8), B2 
                           => n147, ZN => n312);
   U191 : AOI222_X1 port map( A1 => A_shifted(8), A2 => n182, B1 => 
                           zeroSignal(8), B2 => n173, C1 => A_neg_shifted(8), 
                           C2 => n160, ZN => n311);
   U192 : NAND2_X1 port map( A1 => n318, A2 => n317, ZN => Y(9));
   U193 : AOI22_X1 port map( A1 => A_neg(9), A2 => n156, B1 => A_signal(9), B2 
                           => n147, ZN => n318);
   U194 : AOI222_X1 port map( A1 => A_shifted(9), A2 => n182, B1 => 
                           zeroSignal(9), B2 => n173, C1 => A_neg_shifted(9), 
                           C2 => n160, ZN => n317);
   U195 : NAND2_X1 port map( A1 => n190, A2 => n189, ZN => Y(10));
   U196 : AOI22_X1 port map( A1 => A_neg(10), A2 => n151, B1 => A_signal(10), 
                           B2 => n142, ZN => n190);
   U197 : AOI222_X1 port map( A1 => A_shifted(10), A2 => n177, B1 => 
                           zeroSignal(10), B2 => n168, C1 => A_neg_shifted(10),
                           C2 => n165, ZN => n189);
   U198 : NAND2_X1 port map( A1 => n192, A2 => n191, ZN => Y(11));
   U199 : AOI22_X1 port map( A1 => A_neg(11), A2 => n151, B1 => A_signal(11), 
                           B2 => n142, ZN => n192);
   U200 : AOI222_X1 port map( A1 => A_shifted(11), A2 => n177, B1 => 
                           zeroSignal(11), B2 => n168, C1 => A_neg_shifted(11),
                           C2 => n165, ZN => n191);
   U201 : NAND2_X1 port map( A1 => n194, A2 => n193, ZN => Y(12));
   U202 : AOI22_X1 port map( A1 => A_neg(12), A2 => n151, B1 => A_signal(12), 
                           B2 => n142, ZN => n194);
   U203 : AOI222_X1 port map( A1 => A_shifted(12), A2 => n177, B1 => 
                           zeroSignal(12), B2 => n168, C1 => A_neg_shifted(12),
                           C2 => n165, ZN => n193);
   U204 : NAND2_X1 port map( A1 => n196, A2 => n195, ZN => Y(13));
   U205 : AOI22_X1 port map( A1 => A_neg(13), A2 => n151, B1 => A_signal(13), 
                           B2 => n142, ZN => n196);
   U206 : AOI222_X1 port map( A1 => A_shifted(13), A2 => n177, B1 => 
                           zeroSignal(13), B2 => n168, C1 => A_neg_shifted(13),
                           C2 => n164, ZN => n195);
   U207 : NAND2_X1 port map( A1 => n198, A2 => n197, ZN => Y(14));
   U208 : AOI22_X1 port map( A1 => A_neg(14), A2 => n151, B1 => A_signal(14), 
                           B2 => n142, ZN => n198);
   U209 : AOI222_X1 port map( A1 => A_shifted(14), A2 => n177, B1 => 
                           zeroSignal(14), B2 => n168, C1 => A_neg_shifted(14),
                           C2 => n164, ZN => n197);
   U210 : NAND2_X1 port map( A1 => n200, A2 => n199, ZN => Y(15));
   U211 : AOI22_X1 port map( A1 => A_neg(15), A2 => n151, B1 => A_signal(15), 
                           B2 => n142, ZN => n200);
   U212 : AOI222_X1 port map( A1 => A_shifted(15), A2 => n177, B1 => 
                           zeroSignal(15), B2 => n168, C1 => A_neg_shifted(15),
                           C2 => n164, ZN => n199);
   U213 : NAND2_X1 port map( A1 => n202, A2 => n201, ZN => Y(16));
   U214 : AOI22_X1 port map( A1 => A_neg(16), A2 => n151, B1 => A_signal(16), 
                           B2 => n142, ZN => n202);
   U215 : AOI222_X1 port map( A1 => A_shifted(16), A2 => n177, B1 => 
                           zeroSignal(16), B2 => n168, C1 => A_neg_shifted(16),
                           C2 => n164, ZN => n201);
   U216 : NAND2_X1 port map( A1 => n204, A2 => n203, ZN => Y(17));
   U217 : AOI22_X1 port map( A1 => A_neg(17), A2 => n151, B1 => A_signal(17), 
                           B2 => n142, ZN => n204);
   U218 : AOI222_X1 port map( A1 => A_shifted(17), A2 => n177, B1 => 
                           zeroSignal(17), B2 => n168, C1 => A_neg_shifted(17),
                           C2 => n164, ZN => n203);
   U219 : NAND2_X1 port map( A1 => n206, A2 => n205, ZN => Y(18));
   U220 : AOI22_X1 port map( A1 => A_neg(18), A2 => n151, B1 => A_signal(18), 
                           B2 => n142, ZN => n206);
   U221 : AOI222_X1 port map( A1 => A_shifted(18), A2 => n177, B1 => 
                           zeroSignal(18), B2 => n168, C1 => A_neg_shifted(18),
                           C2 => n164, ZN => n205);
   U222 : NAND2_X1 port map( A1 => n208, A2 => n207, ZN => Y(19));
   U223 : AOI22_X1 port map( A1 => A_neg(19), A2 => n151, B1 => A_signal(19), 
                           B2 => n142, ZN => n208);
   U224 : AOI222_X1 port map( A1 => A_shifted(19), A2 => n177, B1 => 
                           zeroSignal(19), B2 => n168, C1 => A_neg_shifted(19),
                           C2 => n164, ZN => n207);
   U225 : NAND2_X1 port map( A1 => n212, A2 => n211, ZN => Y(20));
   U226 : AOI22_X1 port map( A1 => A_neg(20), A2 => n152, B1 => A_signal(20), 
                           B2 => n143, ZN => n212);
   U227 : AOI222_X1 port map( A1 => A_shifted(20), A2 => n178, B1 => 
                           zeroSignal(20), B2 => n169, C1 => A_neg_shifted(20),
                           C2 => n164, ZN => n211);
   U228 : NAND2_X1 port map( A1 => n214, A2 => n213, ZN => Y(21));
   U229 : AOI22_X1 port map( A1 => A_neg(21), A2 => n152, B1 => A_signal(21), 
                           B2 => n143, ZN => n214);
   U230 : AOI222_X1 port map( A1 => A_shifted(21), A2 => n178, B1 => 
                           zeroSignal(21), B2 => n169, C1 => A_neg_shifted(21),
                           C2 => n164, ZN => n213);
   U231 : NAND2_X1 port map( A1 => n216, A2 => n215, ZN => Y(22));
   U232 : AOI22_X1 port map( A1 => A_neg(22), A2 => n152, B1 => A_signal(22), 
                           B2 => n143, ZN => n216);
   U233 : AOI222_X1 port map( A1 => A_shifted(22), A2 => n178, B1 => 
                           zeroSignal(22), B2 => n169, C1 => A_neg_shifted(22),
                           C2 => n164, ZN => n215);
   U234 : NAND2_X1 port map( A1 => n218, A2 => n217, ZN => Y(23));
   U235 : AOI22_X1 port map( A1 => A_neg(23), A2 => n152, B1 => A_signal(23), 
                           B2 => n143, ZN => n218);
   U236 : AOI222_X1 port map( A1 => A_shifted(23), A2 => n178, B1 => 
                           zeroSignal(23), B2 => n169, C1 => A_neg_shifted(23),
                           C2 => n164, ZN => n217);
   U237 : NAND2_X1 port map( A1 => n220, A2 => n219, ZN => Y(24));
   U238 : AOI22_X1 port map( A1 => A_neg(24), A2 => n152, B1 => A_signal(24), 
                           B2 => n143, ZN => n220);
   U239 : AOI222_X1 port map( A1 => A_shifted(24), A2 => n178, B1 => 
                           zeroSignal(24), B2 => n169, C1 => A_neg_shifted(24),
                           C2 => n163, ZN => n219);
   U240 : NAND2_X1 port map( A1 => n222, A2 => n221, ZN => Y(25));
   U241 : AOI22_X1 port map( A1 => A_neg(25), A2 => n152, B1 => A_signal(25), 
                           B2 => n143, ZN => n222);
   U242 : AOI222_X1 port map( A1 => A_shifted(25), A2 => n178, B1 => 
                           zeroSignal(25), B2 => n169, C1 => A_neg_shifted(25),
                           C2 => n163, ZN => n221);
   U243 : AOI222_X1 port map( A1 => A_shifted(27), A2 => n178, B1 => 
                           zeroSignal(27), B2 => n169, C1 => A_neg_shifted(27),
                           C2 => n163, ZN => n225);
   U244 : AOI22_X1 port map( A1 => A_neg(26), A2 => n152, B1 => A_signal(26), 
                           B2 => n143, ZN => n224);

end SYN_BEHAVIORAL_2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity MUX51_MuxNbit64_18 is

   port( zeroSignal, A_signal, A_neg, A_shifted, A_neg_shifted : in 
         std_logic_vector (63 downto 0);  Sel : in std_logic_vector (2 downto 
         0);  Y : out std_logic_vector (63 downto 0));

end MUX51_MuxNbit64_18;

architecture SYN_BEHAVIORAL_2 of MUX51_MuxNbit64_18 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, 
      n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, 
      n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, 
      n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, 
      n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, 
      n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, 
      n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, 
      n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, 
      n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, 
      n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, 
      n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, 
      n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, 
      n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, 
      n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, 
      n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, 
      n320 : std_logic;

begin
   
   U1 : AND3_X1 port map( A1 => n319, A2 => n320, A3 => Sel(2), ZN => n141);
   U2 : BUF_X1 port map( A => n141, Z => n166);
   U3 : BUF_X1 port map( A => n185, Z => n184);
   U4 : BUF_X1 port map( A => n159, Z => n158);
   U5 : BUF_X1 port map( A => n150, Z => n149);
   U6 : BUF_X1 port map( A => n141, Z => n167);
   U7 : BUF_X1 port map( A => n185, Z => n183);
   U8 : BUF_X1 port map( A => n159, Z => n157);
   U9 : BUF_X1 port map( A => n150, Z => n148);
   U10 : BUF_X1 port map( A => n176, Z => n175);
   U11 : BUF_X1 port map( A => n176, Z => n174);
   U12 : BUF_X1 port map( A => n158, Z => n152);
   U13 : BUF_X1 port map( A => n184, Z => n178);
   U14 : BUF_X1 port map( A => n149, Z => n143);
   U15 : BUF_X1 port map( A => n166, Z => n163);
   U16 : BUF_X1 port map( A => n184, Z => n179);
   U17 : BUF_X1 port map( A => n158, Z => n153);
   U18 : BUF_X1 port map( A => n149, Z => n144);
   U19 : BUF_X1 port map( A => n167, Z => n162);
   U20 : BUF_X1 port map( A => n183, Z => n180);
   U21 : BUF_X1 port map( A => n157, Z => n154);
   U22 : BUF_X1 port map( A => n148, Z => n145);
   U23 : BUF_X1 port map( A => n167, Z => n161);
   U24 : BUF_X1 port map( A => n183, Z => n181);
   U25 : BUF_X1 port map( A => n157, Z => n155);
   U26 : BUF_X1 port map( A => n148, Z => n146);
   U27 : BUF_X1 port map( A => n167, Z => n160);
   U28 : BUF_X1 port map( A => n158, Z => n151);
   U29 : BUF_X1 port map( A => n149, Z => n142);
   U30 : BUF_X1 port map( A => n175, Z => n168);
   U31 : BUF_X1 port map( A => n175, Z => n170);
   U32 : BUF_X1 port map( A => n174, Z => n171);
   U33 : BUF_X1 port map( A => n174, Z => n172);
   U34 : BUF_X1 port map( A => n166, Z => n164);
   U35 : BUF_X1 port map( A => n175, Z => n169);
   U36 : BUF_X1 port map( A => n184, Z => n177);
   U37 : BUF_X1 port map( A => n166, Z => n165);
   U38 : BUF_X1 port map( A => n157, Z => n156);
   U39 : BUF_X1 port map( A => n148, Z => n147);
   U40 : BUF_X1 port map( A => n174, Z => n173);
   U41 : BUF_X1 port map( A => n183, Z => n182);
   U42 : INV_X1 port map( A => Sel(1), ZN => n320);
   U43 : BUF_X1 port map( A => n314, Z => n159);
   U44 : NOR3_X1 port map( A1 => Sel(0), A2 => Sel(2), A3 => n320, ZN => n314);
   U45 : BUF_X1 port map( A => n316, Z => n185);
   U46 : NOR3_X1 port map( A1 => n319, A2 => Sel(2), A3 => n320, ZN => n316);
   U47 : INV_X1 port map( A => Sel(0), ZN => n319);
   U48 : BUF_X1 port map( A => n313, Z => n150);
   U49 : NOR3_X1 port map( A1 => Sel(1), A2 => Sel(2), A3 => n319, ZN => n313);
   U50 : BUF_X1 port map( A => n315, Z => n176);
   U51 : NOR2_X1 port map( A1 => n165, A2 => n186, ZN => n315);
   U52 : AOI21_X1 port map( B1 => n319, B2 => n320, A => Sel(2), ZN => n186);
   U53 : NAND2_X1 port map( A1 => n230, A2 => n229, ZN => Y(29));
   U54 : AOI22_X1 port map( A1 => A_neg(29), A2 => n152, B1 => A_signal(29), B2
                           => n143, ZN => n230);
   U55 : NAND2_X1 port map( A1 => n228, A2 => n227, ZN => Y(28));
   U56 : AOI222_X1 port map( A1 => A_shifted(28), A2 => n178, B1 => 
                           zeroSignal(28), B2 => n169, C1 => A_neg_shifted(28),
                           C2 => n163, ZN => n227);
   U57 : NAND2_X1 port map( A1 => n234, A2 => n233, ZN => Y(30));
   U58 : AOI22_X1 port map( A1 => A_neg(30), A2 => n152, B1 => A_signal(30), B2
                           => n143, ZN => n234);
   U59 : AOI222_X1 port map( A1 => A_shifted(30), A2 => n178, B1 => 
                           zeroSignal(30), B2 => n169, C1 => A_neg_shifted(30),
                           C2 => n163, ZN => n233);
   U60 : NAND2_X1 port map( A1 => n236, A2 => n235, ZN => Y(31));
   U61 : AOI22_X1 port map( A1 => A_neg(31), A2 => n153, B1 => A_signal(31), B2
                           => n144, ZN => n236);
   U62 : AOI222_X1 port map( A1 => A_shifted(31), A2 => n179, B1 => 
                           zeroSignal(31), B2 => n170, C1 => A_neg_shifted(31),
                           C2 => n163, ZN => n235);
   U63 : NAND2_X1 port map( A1 => n238, A2 => n237, ZN => Y(32));
   U64 : AOI22_X1 port map( A1 => A_neg(32), A2 => n153, B1 => A_signal(32), B2
                           => n144, ZN => n238);
   U65 : AOI222_X1 port map( A1 => A_shifted(32), A2 => n179, B1 => 
                           zeroSignal(32), B2 => n170, C1 => A_neg_shifted(32),
                           C2 => n163, ZN => n237);
   U66 : NAND2_X1 port map( A1 => n250, A2 => n249, ZN => Y(38));
   U67 : AOI222_X1 port map( A1 => A_shifted(38), A2 => n179, B1 => 
                           zeroSignal(38), B2 => n170, C1 => A_neg_shifted(38),
                           C2 => n162, ZN => n249);
   U68 : AOI22_X1 port map( A1 => A_neg(38), A2 => n153, B1 => A_signal(38), B2
                           => n144, ZN => n250);
   U69 : NAND2_X1 port map( A1 => n252, A2 => n251, ZN => Y(39));
   U70 : AOI222_X1 port map( A1 => A_shifted(39), A2 => n179, B1 => 
                           zeroSignal(39), B2 => n170, C1 => A_neg_shifted(39),
                           C2 => n162, ZN => n251);
   U71 : AOI22_X1 port map( A1 => A_neg(39), A2 => n153, B1 => A_signal(39), B2
                           => n144, ZN => n252);
   U72 : NAND2_X1 port map( A1 => n256, A2 => n255, ZN => Y(40));
   U73 : AOI222_X1 port map( A1 => A_shifted(40), A2 => n179, B1 => 
                           zeroSignal(40), B2 => n170, C1 => A_neg_shifted(40),
                           C2 => n162, ZN => n255);
   U74 : AOI22_X1 port map( A1 => A_neg(40), A2 => n153, B1 => A_signal(40), B2
                           => n144, ZN => n256);
   U75 : NAND2_X1 port map( A1 => n258, A2 => n257, ZN => Y(41));
   U76 : AOI222_X1 port map( A1 => A_shifted(41), A2 => n179, B1 => 
                           zeroSignal(41), B2 => n170, C1 => A_neg_shifted(41),
                           C2 => n162, ZN => n257);
   U77 : AOI22_X1 port map( A1 => A_neg(41), A2 => n153, B1 => A_signal(41), B2
                           => n144, ZN => n258);
   U78 : NAND2_X1 port map( A1 => n264, A2 => n263, ZN => Y(44));
   U79 : AOI222_X1 port map( A1 => A_shifted(44), A2 => n180, B1 => 
                           zeroSignal(44), B2 => n171, C1 => A_neg_shifted(44),
                           C2 => n162, ZN => n263);
   U80 : AOI22_X1 port map( A1 => A_neg(44), A2 => n154, B1 => A_signal(44), B2
                           => n145, ZN => n264);
   U81 : NAND2_X1 port map( A1 => n262, A2 => n261, ZN => Y(43));
   U82 : AOI222_X1 port map( A1 => A_shifted(43), A2 => n180, B1 => 
                           zeroSignal(43), B2 => n171, C1 => A_neg_shifted(43),
                           C2 => n162, ZN => n261);
   U83 : AOI22_X1 port map( A1 => A_neg(43), A2 => n154, B1 => A_signal(43), B2
                           => n145, ZN => n262);
   U84 : NAND2_X1 port map( A1 => n266, A2 => n265, ZN => Y(45));
   U85 : AOI222_X1 port map( A1 => A_shifted(45), A2 => n180, B1 => 
                           zeroSignal(45), B2 => n171, C1 => A_neg_shifted(45),
                           C2 => n162, ZN => n265);
   U86 : AOI22_X1 port map( A1 => A_neg(45), A2 => n154, B1 => A_signal(45), B2
                           => n145, ZN => n266);
   U87 : NAND2_X1 port map( A1 => n240, A2 => n239, ZN => Y(33));
   U88 : AOI22_X1 port map( A1 => A_neg(33), A2 => n153, B1 => A_signal(33), B2
                           => n144, ZN => n240);
   U89 : AOI222_X1 port map( A1 => A_shifted(33), A2 => n179, B1 => 
                           zeroSignal(33), B2 => n170, C1 => A_neg_shifted(33),
                           C2 => n163, ZN => n239);
   U90 : NAND2_X1 port map( A1 => n260, A2 => n259, ZN => Y(42));
   U91 : AOI22_X1 port map( A1 => A_neg(42), A2 => n154, B1 => A_signal(42), B2
                           => n145, ZN => n260);
   U92 : AOI222_X1 port map( A1 => A_shifted(42), A2 => n180, B1 => 
                           zeroSignal(42), B2 => n171, C1 => A_neg_shifted(42),
                           C2 => n162, ZN => n259);
   U93 : NAND2_X1 port map( A1 => n270, A2 => n269, ZN => Y(47));
   U94 : AOI222_X1 port map( A1 => A_shifted(47), A2 => n180, B1 => 
                           zeroSignal(47), B2 => n171, C1 => A_neg_shifted(47),
                           C2 => n161, ZN => n269);
   U95 : AOI22_X1 port map( A1 => A_neg(47), A2 => n154, B1 => A_signal(47), B2
                           => n145, ZN => n270);
   U96 : NAND2_X1 port map( A1 => n274, A2 => n273, ZN => Y(49));
   U97 : AOI222_X1 port map( A1 => A_shifted(49), A2 => n180, B1 => 
                           zeroSignal(49), B2 => n171, C1 => A_neg_shifted(49),
                           C2 => n161, ZN => n273);
   U98 : AOI22_X1 port map( A1 => A_neg(49), A2 => n154, B1 => A_signal(49), B2
                           => n145, ZN => n274);
   U99 : NAND2_X1 port map( A1 => n272, A2 => n271, ZN => Y(48));
   U100 : AOI222_X1 port map( A1 => A_shifted(48), A2 => n180, B1 => 
                           zeroSignal(48), B2 => n171, C1 => A_neg_shifted(48),
                           C2 => n161, ZN => n271);
   U101 : AOI22_X1 port map( A1 => A_neg(48), A2 => n154, B1 => A_signal(48), 
                           B2 => n145, ZN => n272);
   U102 : NAND2_X1 port map( A1 => n278, A2 => n277, ZN => Y(50));
   U103 : AOI222_X1 port map( A1 => A_shifted(50), A2 => n180, B1 => 
                           zeroSignal(50), B2 => n171, C1 => A_neg_shifted(50),
                           C2 => n161, ZN => n277);
   U104 : AOI22_X1 port map( A1 => A_neg(50), A2 => n154, B1 => A_signal(50), 
                           B2 => n145, ZN => n278);
   U105 : NAND2_X1 port map( A1 => n268, A2 => n267, ZN => Y(46));
   U106 : AOI22_X1 port map( A1 => A_neg(46), A2 => n154, B1 => A_signal(46), 
                           B2 => n145, ZN => n268);
   U107 : AOI222_X1 port map( A1 => A_shifted(46), A2 => n180, B1 => 
                           zeroSignal(46), B2 => n171, C1 => A_neg_shifted(46),
                           C2 => n161, ZN => n267);
   U108 : NAND2_X1 port map( A1 => n280, A2 => n279, ZN => Y(51));
   U109 : AOI222_X1 port map( A1 => A_shifted(51), A2 => n180, B1 => 
                           zeroSignal(51), B2 => n171, C1 => A_neg_shifted(51),
                           C2 => n161, ZN => n279);
   U110 : AOI22_X1 port map( A1 => A_neg(51), A2 => n154, B1 => A_signal(51), 
                           B2 => n145, ZN => n280);
   U111 : NAND2_X1 port map( A1 => n284, A2 => n283, ZN => Y(53));
   U112 : AOI222_X1 port map( A1 => A_shifted(53), A2 => n181, B1 => 
                           zeroSignal(53), B2 => n172, C1 => A_neg_shifted(53),
                           C2 => n161, ZN => n283);
   U113 : AOI22_X1 port map( A1 => A_neg(53), A2 => n155, B1 => A_signal(53), 
                           B2 => n146, ZN => n284);
   U114 : NAND2_X1 port map( A1 => n288, A2 => n287, ZN => Y(55));
   U115 : AOI222_X1 port map( A1 => A_shifted(55), A2 => n181, B1 => 
                           zeroSignal(55), B2 => n172, C1 => A_neg_shifted(55),
                           C2 => n161, ZN => n287);
   U116 : AOI22_X1 port map( A1 => A_neg(55), A2 => n155, B1 => A_signal(55), 
                           B2 => n146, ZN => n288);
   U117 : NAND2_X1 port map( A1 => n302, A2 => n301, ZN => Y(61));
   U118 : AOI222_X1 port map( A1 => A_shifted(61), A2 => n181, B1 => 
                           zeroSignal(61), B2 => n172, C1 => A_neg_shifted(61),
                           C2 => n160, ZN => n301);
   U119 : AOI22_X1 port map( A1 => A_neg(61), A2 => n155, B1 => A_signal(61), 
                           B2 => n146, ZN => n302);
   U120 : NAND2_X1 port map( A1 => n286, A2 => n285, ZN => Y(54));
   U121 : AOI222_X1 port map( A1 => A_shifted(54), A2 => n181, B1 => 
                           zeroSignal(54), B2 => n172, C1 => A_neg_shifted(54),
                           C2 => n161, ZN => n285);
   U122 : AOI22_X1 port map( A1 => A_neg(54), A2 => n155, B1 => A_signal(54), 
                           B2 => n146, ZN => n286);
   U123 : NAND2_X1 port map( A1 => n290, A2 => n289, ZN => Y(56));
   U124 : AOI222_X1 port map( A1 => A_shifted(56), A2 => n181, B1 => 
                           zeroSignal(56), B2 => n172, C1 => A_neg_shifted(56),
                           C2 => n161, ZN => n289);
   U125 : AOI22_X1 port map( A1 => A_neg(56), A2 => n155, B1 => A_signal(56), 
                           B2 => n146, ZN => n290);
   U126 : NAND2_X1 port map( A1 => n282, A2 => n281, ZN => Y(52));
   U127 : AOI22_X1 port map( A1 => A_neg(52), A2 => n154, B1 => A_signal(52), 
                           B2 => n145, ZN => n282);
   U128 : AOI222_X1 port map( A1 => A_shifted(52), A2 => n180, B1 => 
                           zeroSignal(52), B2 => n171, C1 => A_neg_shifted(52),
                           C2 => n161, ZN => n281);
   U129 : NAND2_X1 port map( A1 => n292, A2 => n291, ZN => Y(57));
   U130 : AOI222_X1 port map( A1 => A_shifted(57), A2 => n181, B1 => 
                           zeroSignal(57), B2 => n172, C1 => A_neg_shifted(57),
                           C2 => n160, ZN => n291);
   U131 : AOI22_X1 port map( A1 => A_neg(57), A2 => n155, B1 => A_signal(57), 
                           B2 => n146, ZN => n292);
   U132 : NAND2_X1 port map( A1 => n296, A2 => n295, ZN => Y(59));
   U133 : AOI222_X1 port map( A1 => A_shifted(59), A2 => n181, B1 => 
                           zeroSignal(59), B2 => n172, C1 => A_neg_shifted(59),
                           C2 => n160, ZN => n295);
   U134 : AOI22_X1 port map( A1 => A_neg(59), A2 => n155, B1 => A_signal(59), 
                           B2 => n146, ZN => n296);
   U135 : NAND2_X1 port map( A1 => n294, A2 => n293, ZN => Y(58));
   U136 : AOI222_X1 port map( A1 => A_shifted(58), A2 => n181, B1 => 
                           zeroSignal(58), B2 => n172, C1 => A_neg_shifted(58),
                           C2 => n160, ZN => n293);
   U137 : AOI22_X1 port map( A1 => A_neg(58), A2 => n155, B1 => A_signal(58), 
                           B2 => n146, ZN => n294);
   U138 : NAND2_X1 port map( A1 => n242, A2 => n241, ZN => Y(34));
   U139 : AOI222_X1 port map( A1 => A_shifted(34), A2 => n179, B1 => 
                           zeroSignal(34), B2 => n170, C1 => A_neg_shifted(34),
                           C2 => n163, ZN => n241);
   U140 : AOI22_X1 port map( A1 => A_neg(34), A2 => n153, B1 => A_signal(34), 
                           B2 => n144, ZN => n242);
   U141 : NAND2_X1 port map( A1 => n300, A2 => n299, ZN => Y(60));
   U142 : AOI222_X1 port map( A1 => A_shifted(60), A2 => n181, B1 => 
                           zeroSignal(60), B2 => n172, C1 => A_neg_shifted(60),
                           C2 => n160, ZN => n299);
   U143 : AOI22_X1 port map( A1 => A_neg(60), A2 => n155, B1 => A_signal(60), 
                           B2 => n146, ZN => n300);
   U144 : NAND2_X1 port map( A1 => n244, A2 => n243, ZN => Y(35));
   U145 : AOI222_X1 port map( A1 => A_shifted(35), A2 => n179, B1 => 
                           zeroSignal(35), B2 => n170, C1 => A_neg_shifted(35),
                           C2 => n162, ZN => n243);
   U146 : AOI22_X1 port map( A1 => A_neg(35), A2 => n153, B1 => A_signal(35), 
                           B2 => n144, ZN => n244);
   U147 : NAND2_X1 port map( A1 => n304, A2 => n303, ZN => Y(62));
   U148 : AOI222_X1 port map( A1 => A_shifted(62), A2 => n181, B1 => 
                           zeroSignal(62), B2 => n172, C1 => A_neg_shifted(62),
                           C2 => n160, ZN => n303);
   U149 : AOI22_X1 port map( A1 => A_neg(62), A2 => n155, B1 => A_signal(62), 
                           B2 => n146, ZN => n304);
   U150 : NAND2_X1 port map( A1 => n248, A2 => n247, ZN => Y(37));
   U151 : AOI222_X1 port map( A1 => A_shifted(37), A2 => n179, B1 => 
                           zeroSignal(37), B2 => n170, C1 => A_neg_shifted(37),
                           C2 => n162, ZN => n247);
   U152 : AOI22_X1 port map( A1 => A_neg(37), A2 => n153, B1 => A_signal(37), 
                           B2 => n144, ZN => n248);
   U153 : NAND2_X1 port map( A1 => n246, A2 => n245, ZN => Y(36));
   U154 : AOI222_X1 port map( A1 => A_shifted(36), A2 => n179, B1 => 
                           zeroSignal(36), B2 => n170, C1 => A_neg_shifted(36),
                           C2 => n162, ZN => n245);
   U155 : AOI22_X1 port map( A1 => A_neg(36), A2 => n153, B1 => A_signal(36), 
                           B2 => n144, ZN => n246);
   U156 : NAND2_X1 port map( A1 => n306, A2 => n305, ZN => Y(63));
   U157 : AOI222_X1 port map( A1 => A_shifted(63), A2 => n181, B1 => 
                           zeroSignal(63), B2 => n172, C1 => A_neg_shifted(63),
                           C2 => n160, ZN => n305);
   U158 : AOI22_X1 port map( A1 => A_neg(63), A2 => n155, B1 => A_signal(63), 
                           B2 => n146, ZN => n306);
   U159 : NAND2_X1 port map( A1 => n188, A2 => n187, ZN => Y(0));
   U160 : AOI22_X1 port map( A1 => A_neg(0), A2 => n151, B1 => A_signal(0), B2 
                           => n142, ZN => n188);
   U161 : AOI222_X1 port map( A1 => A_shifted(0), A2 => n177, B1 => 
                           zeroSignal(0), B2 => n168, C1 => A_neg_shifted(0), 
                           C2 => n165, ZN => n187);
   U162 : NAND2_X1 port map( A1 => n210, A2 => n209, ZN => Y(1));
   U163 : AOI22_X1 port map( A1 => A_neg(1), A2 => n151, B1 => A_signal(1), B2 
                           => n142, ZN => n210);
   U164 : AOI222_X1 port map( A1 => A_shifted(1), A2 => n177, B1 => 
                           zeroSignal(1), B2 => n168, C1 => A_neg_shifted(1), 
                           C2 => n164, ZN => n209);
   U165 : NAND2_X1 port map( A1 => n232, A2 => n231, ZN => Y(2));
   U166 : AOI22_X1 port map( A1 => A_neg(2), A2 => n152, B1 => A_signal(2), B2 
                           => n143, ZN => n232);
   U167 : AOI222_X1 port map( A1 => A_shifted(2), A2 => n178, B1 => 
                           zeroSignal(2), B2 => n169, C1 => A_neg_shifted(2), 
                           C2 => n163, ZN => n231);
   U168 : NAND2_X1 port map( A1 => n254, A2 => n253, ZN => Y(3));
   U169 : AOI22_X1 port map( A1 => A_neg(3), A2 => n153, B1 => A_signal(3), B2 
                           => n144, ZN => n254);
   U170 : AOI222_X1 port map( A1 => A_shifted(3), A2 => n179, B1 => 
                           zeroSignal(3), B2 => n170, C1 => A_neg_shifted(3), 
                           C2 => n162, ZN => n253);
   U171 : NAND2_X1 port map( A1 => n276, A2 => n275, ZN => Y(4));
   U172 : AOI22_X1 port map( A1 => A_neg(4), A2 => n154, B1 => A_signal(4), B2 
                           => n145, ZN => n276);
   U173 : AOI222_X1 port map( A1 => A_shifted(4), A2 => n180, B1 => 
                           zeroSignal(4), B2 => n171, C1 => A_neg_shifted(4), 
                           C2 => n161, ZN => n275);
   U174 : NAND2_X1 port map( A1 => n298, A2 => n297, ZN => Y(5));
   U175 : AOI22_X1 port map( A1 => A_neg(5), A2 => n155, B1 => A_signal(5), B2 
                           => n146, ZN => n298);
   U176 : AOI222_X1 port map( A1 => A_shifted(5), A2 => n181, B1 => 
                           zeroSignal(5), B2 => n172, C1 => A_neg_shifted(5), 
                           C2 => n160, ZN => n297);
   U177 : NAND2_X1 port map( A1 => n308, A2 => n307, ZN => Y(6));
   U178 : AOI22_X1 port map( A1 => A_neg(6), A2 => n156, B1 => A_signal(6), B2 
                           => n147, ZN => n308);
   U179 : AOI222_X1 port map( A1 => A_shifted(6), A2 => n182, B1 => 
                           zeroSignal(6), B2 => n173, C1 => A_neg_shifted(6), 
                           C2 => n160, ZN => n307);
   U180 : NAND2_X1 port map( A1 => n310, A2 => n309, ZN => Y(7));
   U181 : AOI22_X1 port map( A1 => A_neg(7), A2 => n156, B1 => A_signal(7), B2 
                           => n147, ZN => n310);
   U182 : AOI222_X1 port map( A1 => A_shifted(7), A2 => n182, B1 => 
                           zeroSignal(7), B2 => n173, C1 => A_neg_shifted(7), 
                           C2 => n160, ZN => n309);
   U183 : NAND2_X1 port map( A1 => n312, A2 => n311, ZN => Y(8));
   U184 : AOI22_X1 port map( A1 => A_neg(8), A2 => n156, B1 => A_signal(8), B2 
                           => n147, ZN => n312);
   U185 : AOI222_X1 port map( A1 => A_shifted(8), A2 => n182, B1 => 
                           zeroSignal(8), B2 => n173, C1 => A_neg_shifted(8), 
                           C2 => n160, ZN => n311);
   U186 : NAND2_X1 port map( A1 => n318, A2 => n317, ZN => Y(9));
   U187 : AOI22_X1 port map( A1 => A_neg(9), A2 => n156, B1 => A_signal(9), B2 
                           => n147, ZN => n318);
   U188 : AOI222_X1 port map( A1 => A_shifted(9), A2 => n182, B1 => 
                           zeroSignal(9), B2 => n173, C1 => A_neg_shifted(9), 
                           C2 => n160, ZN => n317);
   U189 : NAND2_X1 port map( A1 => n190, A2 => n189, ZN => Y(10));
   U190 : AOI22_X1 port map( A1 => A_neg(10), A2 => n151, B1 => A_signal(10), 
                           B2 => n142, ZN => n190);
   U191 : AOI222_X1 port map( A1 => A_shifted(10), A2 => n177, B1 => 
                           zeroSignal(10), B2 => n168, C1 => A_neg_shifted(10),
                           C2 => n165, ZN => n189);
   U192 : NAND2_X1 port map( A1 => n192, A2 => n191, ZN => Y(11));
   U193 : AOI22_X1 port map( A1 => A_neg(11), A2 => n151, B1 => A_signal(11), 
                           B2 => n142, ZN => n192);
   U194 : AOI222_X1 port map( A1 => A_shifted(11), A2 => n177, B1 => 
                           zeroSignal(11), B2 => n168, C1 => A_neg_shifted(11),
                           C2 => n165, ZN => n191);
   U195 : NAND2_X1 port map( A1 => n194, A2 => n193, ZN => Y(12));
   U196 : AOI22_X1 port map( A1 => A_neg(12), A2 => n151, B1 => A_signal(12), 
                           B2 => n142, ZN => n194);
   U197 : AOI222_X1 port map( A1 => A_shifted(12), A2 => n177, B1 => 
                           zeroSignal(12), B2 => n168, C1 => A_neg_shifted(12),
                           C2 => n165, ZN => n193);
   U198 : NAND2_X1 port map( A1 => n196, A2 => n195, ZN => Y(13));
   U199 : AOI22_X1 port map( A1 => A_neg(13), A2 => n151, B1 => A_signal(13), 
                           B2 => n142, ZN => n196);
   U200 : AOI222_X1 port map( A1 => A_shifted(13), A2 => n177, B1 => 
                           zeroSignal(13), B2 => n168, C1 => A_neg_shifted(13),
                           C2 => n164, ZN => n195);
   U201 : NAND2_X1 port map( A1 => n198, A2 => n197, ZN => Y(14));
   U202 : AOI22_X1 port map( A1 => A_neg(14), A2 => n151, B1 => A_signal(14), 
                           B2 => n142, ZN => n198);
   U203 : AOI222_X1 port map( A1 => A_shifted(14), A2 => n177, B1 => 
                           zeroSignal(14), B2 => n168, C1 => A_neg_shifted(14),
                           C2 => n164, ZN => n197);
   U204 : NAND2_X1 port map( A1 => n200, A2 => n199, ZN => Y(15));
   U205 : AOI22_X1 port map( A1 => A_neg(15), A2 => n151, B1 => A_signal(15), 
                           B2 => n142, ZN => n200);
   U206 : AOI222_X1 port map( A1 => A_shifted(15), A2 => n177, B1 => 
                           zeroSignal(15), B2 => n168, C1 => A_neg_shifted(15),
                           C2 => n164, ZN => n199);
   U207 : NAND2_X1 port map( A1 => n202, A2 => n201, ZN => Y(16));
   U208 : AOI22_X1 port map( A1 => A_neg(16), A2 => n151, B1 => A_signal(16), 
                           B2 => n142, ZN => n202);
   U209 : AOI222_X1 port map( A1 => A_shifted(16), A2 => n177, B1 => 
                           zeroSignal(16), B2 => n168, C1 => A_neg_shifted(16),
                           C2 => n164, ZN => n201);
   U210 : NAND2_X1 port map( A1 => n204, A2 => n203, ZN => Y(17));
   U211 : AOI22_X1 port map( A1 => A_neg(17), A2 => n151, B1 => A_signal(17), 
                           B2 => n142, ZN => n204);
   U212 : AOI222_X1 port map( A1 => A_shifted(17), A2 => n177, B1 => 
                           zeroSignal(17), B2 => n168, C1 => A_neg_shifted(17),
                           C2 => n164, ZN => n203);
   U213 : NAND2_X1 port map( A1 => n206, A2 => n205, ZN => Y(18));
   U214 : AOI22_X1 port map( A1 => A_neg(18), A2 => n151, B1 => A_signal(18), 
                           B2 => n142, ZN => n206);
   U215 : AOI222_X1 port map( A1 => A_shifted(18), A2 => n177, B1 => 
                           zeroSignal(18), B2 => n168, C1 => A_neg_shifted(18),
                           C2 => n164, ZN => n205);
   U216 : NAND2_X1 port map( A1 => n208, A2 => n207, ZN => Y(19));
   U217 : AOI22_X1 port map( A1 => A_neg(19), A2 => n151, B1 => A_signal(19), 
                           B2 => n142, ZN => n208);
   U218 : AOI222_X1 port map( A1 => A_shifted(19), A2 => n177, B1 => 
                           zeroSignal(19), B2 => n168, C1 => A_neg_shifted(19),
                           C2 => n164, ZN => n207);
   U219 : NAND2_X1 port map( A1 => n212, A2 => n211, ZN => Y(20));
   U220 : AOI22_X1 port map( A1 => A_neg(20), A2 => n152, B1 => A_signal(20), 
                           B2 => n143, ZN => n212);
   U221 : AOI222_X1 port map( A1 => A_shifted(20), A2 => n178, B1 => 
                           zeroSignal(20), B2 => n169, C1 => A_neg_shifted(20),
                           C2 => n164, ZN => n211);
   U222 : NAND2_X1 port map( A1 => n214, A2 => n213, ZN => Y(21));
   U223 : AOI22_X1 port map( A1 => A_neg(21), A2 => n152, B1 => A_signal(21), 
                           B2 => n143, ZN => n214);
   U224 : AOI222_X1 port map( A1 => A_shifted(21), A2 => n178, B1 => 
                           zeroSignal(21), B2 => n169, C1 => A_neg_shifted(21),
                           C2 => n164, ZN => n213);
   U225 : NAND2_X1 port map( A1 => n216, A2 => n215, ZN => Y(22));
   U226 : AOI22_X1 port map( A1 => A_neg(22), A2 => n152, B1 => A_signal(22), 
                           B2 => n143, ZN => n216);
   U227 : AOI222_X1 port map( A1 => A_shifted(22), A2 => n178, B1 => 
                           zeroSignal(22), B2 => n169, C1 => A_neg_shifted(22),
                           C2 => n164, ZN => n215);
   U228 : NAND2_X1 port map( A1 => n218, A2 => n217, ZN => Y(23));
   U229 : AOI22_X1 port map( A1 => A_neg(23), A2 => n152, B1 => A_signal(23), 
                           B2 => n143, ZN => n218);
   U230 : AOI222_X1 port map( A1 => A_shifted(23), A2 => n178, B1 => 
                           zeroSignal(23), B2 => n169, C1 => A_neg_shifted(23),
                           C2 => n164, ZN => n217);
   U231 : NAND2_X1 port map( A1 => n220, A2 => n219, ZN => Y(24));
   U232 : AOI22_X1 port map( A1 => A_neg(24), A2 => n152, B1 => A_signal(24), 
                           B2 => n143, ZN => n220);
   U233 : AOI222_X1 port map( A1 => A_shifted(24), A2 => n178, B1 => 
                           zeroSignal(24), B2 => n169, C1 => A_neg_shifted(24),
                           C2 => n163, ZN => n219);
   U234 : NAND2_X1 port map( A1 => n222, A2 => n221, ZN => Y(25));
   U235 : AOI22_X1 port map( A1 => A_neg(25), A2 => n152, B1 => A_signal(25), 
                           B2 => n143, ZN => n222);
   U236 : AOI222_X1 port map( A1 => A_shifted(25), A2 => n178, B1 => 
                           zeroSignal(25), B2 => n169, C1 => A_neg_shifted(25),
                           C2 => n163, ZN => n221);
   U237 : NAND2_X1 port map( A1 => n224, A2 => n223, ZN => Y(26));
   U238 : AOI22_X1 port map( A1 => A_neg(26), A2 => n152, B1 => A_signal(26), 
                           B2 => n143, ZN => n224);
   U239 : AOI222_X1 port map( A1 => A_shifted(26), A2 => n178, B1 => 
                           zeroSignal(26), B2 => n169, C1 => A_neg_shifted(26),
                           C2 => n163, ZN => n223);
   U240 : NAND2_X1 port map( A1 => n226, A2 => n225, ZN => Y(27));
   U241 : AOI22_X1 port map( A1 => A_neg(27), A2 => n152, B1 => A_signal(27), 
                           B2 => n143, ZN => n226);
   U242 : AOI222_X1 port map( A1 => A_shifted(27), A2 => n178, B1 => 
                           zeroSignal(27), B2 => n169, C1 => A_neg_shifted(27),
                           C2 => n163, ZN => n225);
   U243 : AOI222_X1 port map( A1 => A_shifted(29), A2 => n178, B1 => 
                           zeroSignal(29), B2 => n169, C1 => A_neg_shifted(29),
                           C2 => n163, ZN => n229);
   U244 : AOI22_X1 port map( A1 => A_neg(28), A2 => n152, B1 => A_signal(28), 
                           B2 => n143, ZN => n228);

end SYN_BEHAVIORAL_2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity MUX51_MuxNbit64_17 is

   port( zeroSignal, A_signal, A_neg, A_shifted, A_neg_shifted : in 
         std_logic_vector (63 downto 0);  Sel : in std_logic_vector (2 downto 
         0);  Y : out std_logic_vector (63 downto 0));

end MUX51_MuxNbit64_17;

architecture SYN_BEHAVIORAL_2 of MUX51_MuxNbit64_17 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, 
      n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, 
      n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, 
      n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, 
      n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, 
      n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, 
      n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, 
      n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, 
      n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, 
      n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, 
      n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, 
      n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, 
      n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, 
      n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, 
      n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, 
      n320 : std_logic;

begin
   
   U1 : AND3_X1 port map( A1 => n319, A2 => n320, A3 => Sel(2), ZN => n141);
   U2 : BUF_X1 port map( A => n141, Z => n166);
   U3 : BUF_X1 port map( A => n185, Z => n184);
   U4 : BUF_X1 port map( A => n159, Z => n158);
   U5 : BUF_X1 port map( A => n150, Z => n149);
   U6 : BUF_X1 port map( A => n141, Z => n167);
   U7 : BUF_X1 port map( A => n185, Z => n183);
   U8 : BUF_X1 port map( A => n159, Z => n157);
   U9 : BUF_X1 port map( A => n150, Z => n148);
   U10 : BUF_X1 port map( A => n176, Z => n175);
   U11 : BUF_X1 port map( A => n176, Z => n174);
   U12 : BUF_X1 port map( A => n158, Z => n153);
   U13 : BUF_X1 port map( A => n184, Z => n179);
   U14 : BUF_X1 port map( A => n149, Z => n144);
   U15 : BUF_X1 port map( A => n166, Z => n163);
   U16 : BUF_X1 port map( A => n149, Z => n143);
   U17 : BUF_X1 port map( A => n158, Z => n152);
   U18 : BUF_X1 port map( A => n167, Z => n162);
   U19 : BUF_X1 port map( A => n183, Z => n180);
   U20 : BUF_X1 port map( A => n157, Z => n154);
   U21 : BUF_X1 port map( A => n148, Z => n145);
   U22 : BUF_X1 port map( A => n167, Z => n161);
   U23 : BUF_X1 port map( A => n183, Z => n181);
   U24 : BUF_X1 port map( A => n157, Z => n155);
   U25 : BUF_X1 port map( A => n148, Z => n146);
   U26 : BUF_X1 port map( A => n167, Z => n160);
   U27 : BUF_X1 port map( A => n158, Z => n151);
   U28 : BUF_X1 port map( A => n149, Z => n142);
   U29 : BUF_X1 port map( A => n175, Z => n168);
   U30 : BUF_X1 port map( A => n175, Z => n169);
   U31 : BUF_X1 port map( A => n174, Z => n171);
   U32 : BUF_X1 port map( A => n174, Z => n172);
   U33 : BUF_X1 port map( A => n166, Z => n164);
   U34 : BUF_X1 port map( A => n175, Z => n170);
   U35 : BUF_X1 port map( A => n184, Z => n177);
   U36 : BUF_X1 port map( A => n184, Z => n178);
   U37 : BUF_X1 port map( A => n166, Z => n165);
   U38 : BUF_X1 port map( A => n157, Z => n156);
   U39 : BUF_X1 port map( A => n148, Z => n147);
   U40 : BUF_X1 port map( A => n174, Z => n173);
   U41 : BUF_X1 port map( A => n183, Z => n182);
   U42 : INV_X1 port map( A => Sel(1), ZN => n320);
   U43 : BUF_X1 port map( A => n314, Z => n159);
   U44 : NOR3_X1 port map( A1 => Sel(0), A2 => Sel(2), A3 => n320, ZN => n314);
   U45 : BUF_X1 port map( A => n316, Z => n185);
   U46 : NOR3_X1 port map( A1 => n319, A2 => Sel(2), A3 => n320, ZN => n316);
   U47 : INV_X1 port map( A => Sel(0), ZN => n319);
   U48 : BUF_X1 port map( A => n313, Z => n150);
   U49 : NOR3_X1 port map( A1 => Sel(1), A2 => Sel(2), A3 => n319, ZN => n313);
   U50 : BUF_X1 port map( A => n315, Z => n176);
   U51 : NOR2_X1 port map( A1 => n165, A2 => n186, ZN => n315);
   U52 : AOI21_X1 port map( B1 => n319, B2 => n320, A => Sel(2), ZN => n186);
   U53 : NAND2_X1 port map( A1 => n236, A2 => n235, ZN => Y(31));
   U54 : AOI22_X1 port map( A1 => A_neg(31), A2 => n153, B1 => A_signal(31), B2
                           => n144, ZN => n236);
   U55 : NAND2_X1 port map( A1 => n238, A2 => n237, ZN => Y(32));
   U56 : AOI22_X1 port map( A1 => A_neg(32), A2 => n153, B1 => A_signal(32), B2
                           => n144, ZN => n238);
   U57 : AOI222_X1 port map( A1 => A_shifted(32), A2 => n179, B1 => 
                           zeroSignal(32), B2 => n170, C1 => A_neg_shifted(32),
                           C2 => n163, ZN => n237);
   U58 : NAND2_X1 port map( A1 => n234, A2 => n233, ZN => Y(30));
   U59 : AOI222_X1 port map( A1 => A_shifted(30), A2 => n178, B1 => 
                           zeroSignal(30), B2 => n169, C1 => A_neg_shifted(30),
                           C2 => n163, ZN => n233);
   U60 : NAND2_X1 port map( A1 => n240, A2 => n239, ZN => Y(33));
   U61 : AOI22_X1 port map( A1 => A_neg(33), A2 => n153, B1 => A_signal(33), B2
                           => n144, ZN => n240);
   U62 : AOI222_X1 port map( A1 => A_shifted(33), A2 => n179, B1 => 
                           zeroSignal(33), B2 => n170, C1 => A_neg_shifted(33),
                           C2 => n163, ZN => n239);
   U63 : NAND2_X1 port map( A1 => n242, A2 => n241, ZN => Y(34));
   U64 : AOI22_X1 port map( A1 => A_neg(34), A2 => n153, B1 => A_signal(34), B2
                           => n144, ZN => n242);
   U65 : AOI222_X1 port map( A1 => A_shifted(34), A2 => n179, B1 => 
                           zeroSignal(34), B2 => n170, C1 => A_neg_shifted(34),
                           C2 => n163, ZN => n241);
   U66 : NAND2_X1 port map( A1 => n256, A2 => n255, ZN => Y(40));
   U67 : AOI222_X1 port map( A1 => A_shifted(40), A2 => n179, B1 => 
                           zeroSignal(40), B2 => n170, C1 => A_neg_shifted(40),
                           C2 => n162, ZN => n255);
   U68 : AOI22_X1 port map( A1 => A_neg(40), A2 => n153, B1 => A_signal(40), B2
                           => n144, ZN => n256);
   U69 : NAND2_X1 port map( A1 => n258, A2 => n257, ZN => Y(41));
   U70 : AOI222_X1 port map( A1 => A_shifted(41), A2 => n179, B1 => 
                           zeroSignal(41), B2 => n170, C1 => A_neg_shifted(41),
                           C2 => n162, ZN => n257);
   U71 : AOI22_X1 port map( A1 => A_neg(41), A2 => n153, B1 => A_signal(41), B2
                           => n144, ZN => n258);
   U72 : NAND2_X1 port map( A1 => n260, A2 => n259, ZN => Y(42));
   U73 : AOI222_X1 port map( A1 => A_shifted(42), A2 => n180, B1 => 
                           zeroSignal(42), B2 => n171, C1 => A_neg_shifted(42),
                           C2 => n162, ZN => n259);
   U74 : AOI22_X1 port map( A1 => A_neg(42), A2 => n154, B1 => A_signal(42), B2
                           => n145, ZN => n260);
   U75 : NAND2_X1 port map( A1 => n262, A2 => n261, ZN => Y(43));
   U76 : AOI222_X1 port map( A1 => A_shifted(43), A2 => n180, B1 => 
                           zeroSignal(43), B2 => n171, C1 => A_neg_shifted(43),
                           C2 => n162, ZN => n261);
   U77 : AOI22_X1 port map( A1 => A_neg(43), A2 => n154, B1 => A_signal(43), B2
                           => n145, ZN => n262);
   U78 : NAND2_X1 port map( A1 => n268, A2 => n267, ZN => Y(46));
   U79 : AOI222_X1 port map( A1 => A_shifted(46), A2 => n180, B1 => 
                           zeroSignal(46), B2 => n171, C1 => A_neg_shifted(46),
                           C2 => n161, ZN => n267);
   U80 : AOI22_X1 port map( A1 => A_neg(46), A2 => n154, B1 => A_signal(46), B2
                           => n145, ZN => n268);
   U81 : NAND2_X1 port map( A1 => n266, A2 => n265, ZN => Y(45));
   U82 : AOI222_X1 port map( A1 => A_shifted(45), A2 => n180, B1 => 
                           zeroSignal(45), B2 => n171, C1 => A_neg_shifted(45),
                           C2 => n162, ZN => n265);
   U83 : AOI22_X1 port map( A1 => A_neg(45), A2 => n154, B1 => A_signal(45), B2
                           => n145, ZN => n266);
   U84 : NAND2_X1 port map( A1 => n270, A2 => n269, ZN => Y(47));
   U85 : AOI222_X1 port map( A1 => A_shifted(47), A2 => n180, B1 => 
                           zeroSignal(47), B2 => n171, C1 => A_neg_shifted(47),
                           C2 => n161, ZN => n269);
   U86 : AOI22_X1 port map( A1 => A_neg(47), A2 => n154, B1 => A_signal(47), B2
                           => n145, ZN => n270);
   U87 : NAND2_X1 port map( A1 => n264, A2 => n263, ZN => Y(44));
   U88 : AOI22_X1 port map( A1 => A_neg(44), A2 => n154, B1 => A_signal(44), B2
                           => n145, ZN => n264);
   U89 : AOI222_X1 port map( A1 => A_shifted(44), A2 => n180, B1 => 
                           zeroSignal(44), B2 => n171, C1 => A_neg_shifted(44),
                           C2 => n162, ZN => n263);
   U90 : NAND2_X1 port map( A1 => n274, A2 => n273, ZN => Y(49));
   U91 : AOI222_X1 port map( A1 => A_shifted(49), A2 => n180, B1 => 
                           zeroSignal(49), B2 => n171, C1 => A_neg_shifted(49),
                           C2 => n161, ZN => n273);
   U92 : AOI22_X1 port map( A1 => A_neg(49), A2 => n154, B1 => A_signal(49), B2
                           => n145, ZN => n274);
   U93 : NAND2_X1 port map( A1 => n244, A2 => n243, ZN => Y(35));
   U94 : AOI22_X1 port map( A1 => A_neg(35), A2 => n153, B1 => A_signal(35), B2
                           => n144, ZN => n244);
   U95 : AOI222_X1 port map( A1 => A_shifted(35), A2 => n179, B1 => 
                           zeroSignal(35), B2 => n170, C1 => A_neg_shifted(35),
                           C2 => n162, ZN => n243);
   U96 : NAND2_X1 port map( A1 => n280, A2 => n279, ZN => Y(51));
   U97 : AOI222_X1 port map( A1 => A_shifted(51), A2 => n180, B1 => 
                           zeroSignal(51), B2 => n171, C1 => A_neg_shifted(51),
                           C2 => n161, ZN => n279);
   U98 : AOI22_X1 port map( A1 => A_neg(51), A2 => n154, B1 => A_signal(51), B2
                           => n145, ZN => n280);
   U99 : NAND2_X1 port map( A1 => n278, A2 => n277, ZN => Y(50));
   U100 : AOI222_X1 port map( A1 => A_shifted(50), A2 => n180, B1 => 
                           zeroSignal(50), B2 => n171, C1 => A_neg_shifted(50),
                           C2 => n161, ZN => n277);
   U101 : AOI22_X1 port map( A1 => A_neg(50), A2 => n154, B1 => A_signal(50), 
                           B2 => n145, ZN => n278);
   U102 : NAND2_X1 port map( A1 => n306, A2 => n305, ZN => Y(63));
   U103 : AOI222_X1 port map( A1 => A_shifted(63), A2 => n181, B1 => 
                           zeroSignal(63), B2 => n172, C1 => A_neg_shifted(63),
                           C2 => n160, ZN => n305);
   U104 : AOI22_X1 port map( A1 => A_neg(63), A2 => n155, B1 => A_signal(63), 
                           B2 => n146, ZN => n306);
   U105 : NAND2_X1 port map( A1 => n282, A2 => n281, ZN => Y(52));
   U106 : AOI222_X1 port map( A1 => A_shifted(52), A2 => n180, B1 => 
                           zeroSignal(52), B2 => n171, C1 => A_neg_shifted(52),
                           C2 => n161, ZN => n281);
   U107 : AOI22_X1 port map( A1 => A_neg(52), A2 => n154, B1 => A_signal(52), 
                           B2 => n145, ZN => n282);
   U108 : NAND2_X1 port map( A1 => n272, A2 => n271, ZN => Y(48));
   U109 : AOI22_X1 port map( A1 => A_neg(48), A2 => n154, B1 => A_signal(48), 
                           B2 => n145, ZN => n272);
   U110 : AOI222_X1 port map( A1 => A_shifted(48), A2 => n180, B1 => 
                           zeroSignal(48), B2 => n171, C1 => A_neg_shifted(48),
                           C2 => n161, ZN => n271);
   U111 : NAND2_X1 port map( A1 => n284, A2 => n283, ZN => Y(53));
   U112 : AOI222_X1 port map( A1 => A_shifted(53), A2 => n181, B1 => 
                           zeroSignal(53), B2 => n172, C1 => A_neg_shifted(53),
                           C2 => n161, ZN => n283);
   U113 : AOI22_X1 port map( A1 => A_neg(53), A2 => n155, B1 => A_signal(53), 
                           B2 => n146, ZN => n284);
   U114 : NAND2_X1 port map( A1 => n288, A2 => n287, ZN => Y(55));
   U115 : AOI222_X1 port map( A1 => A_shifted(55), A2 => n181, B1 => 
                           zeroSignal(55), B2 => n172, C1 => A_neg_shifted(55),
                           C2 => n161, ZN => n287);
   U116 : AOI22_X1 port map( A1 => A_neg(55), A2 => n155, B1 => A_signal(55), 
                           B2 => n146, ZN => n288);
   U117 : NAND2_X1 port map( A1 => n292, A2 => n291, ZN => Y(57));
   U118 : AOI222_X1 port map( A1 => A_shifted(57), A2 => n181, B1 => 
                           zeroSignal(57), B2 => n172, C1 => A_neg_shifted(57),
                           C2 => n160, ZN => n291);
   U119 : AOI22_X1 port map( A1 => A_neg(57), A2 => n155, B1 => A_signal(57), 
                           B2 => n146, ZN => n292);
   U120 : NAND2_X1 port map( A1 => n290, A2 => n289, ZN => Y(56));
   U121 : AOI222_X1 port map( A1 => A_shifted(56), A2 => n181, B1 => 
                           zeroSignal(56), B2 => n172, C1 => A_neg_shifted(56),
                           C2 => n161, ZN => n289);
   U122 : AOI22_X1 port map( A1 => A_neg(56), A2 => n155, B1 => A_signal(56), 
                           B2 => n146, ZN => n290);
   U123 : NAND2_X1 port map( A1 => n304, A2 => n303, ZN => Y(62));
   U124 : AOI222_X1 port map( A1 => A_shifted(62), A2 => n181, B1 => 
                           zeroSignal(62), B2 => n172, C1 => A_neg_shifted(62),
                           C2 => n160, ZN => n303);
   U125 : AOI22_X1 port map( A1 => A_neg(62), A2 => n155, B1 => A_signal(62), 
                           B2 => n146, ZN => n304);
   U126 : NAND2_X1 port map( A1 => n294, A2 => n293, ZN => Y(58));
   U127 : AOI222_X1 port map( A1 => A_shifted(58), A2 => n181, B1 => 
                           zeroSignal(58), B2 => n172, C1 => A_neg_shifted(58),
                           C2 => n160, ZN => n293);
   U128 : AOI22_X1 port map( A1 => A_neg(58), A2 => n155, B1 => A_signal(58), 
                           B2 => n146, ZN => n294);
   U129 : NAND2_X1 port map( A1 => n302, A2 => n301, ZN => Y(61));
   U130 : AOI222_X1 port map( A1 => A_shifted(61), A2 => n181, B1 => 
                           zeroSignal(61), B2 => n172, C1 => A_neg_shifted(61),
                           C2 => n160, ZN => n301);
   U131 : AOI22_X1 port map( A1 => A_neg(61), A2 => n155, B1 => A_signal(61), 
                           B2 => n146, ZN => n302);
   U132 : NAND2_X1 port map( A1 => n286, A2 => n285, ZN => Y(54));
   U133 : AOI22_X1 port map( A1 => A_neg(54), A2 => n155, B1 => A_signal(54), 
                           B2 => n146, ZN => n286);
   U134 : AOI222_X1 port map( A1 => A_shifted(54), A2 => n181, B1 => 
                           zeroSignal(54), B2 => n172, C1 => A_neg_shifted(54),
                           C2 => n161, ZN => n285);
   U135 : NAND2_X1 port map( A1 => n296, A2 => n295, ZN => Y(59));
   U136 : AOI222_X1 port map( A1 => A_shifted(59), A2 => n181, B1 => 
                           zeroSignal(59), B2 => n172, C1 => A_neg_shifted(59),
                           C2 => n160, ZN => n295);
   U137 : AOI22_X1 port map( A1 => A_neg(59), A2 => n155, B1 => A_signal(59), 
                           B2 => n146, ZN => n296);
   U138 : NAND2_X1 port map( A1 => n300, A2 => n299, ZN => Y(60));
   U139 : AOI222_X1 port map( A1 => A_shifted(60), A2 => n181, B1 => 
                           zeroSignal(60), B2 => n172, C1 => A_neg_shifted(60),
                           C2 => n160, ZN => n299);
   U140 : AOI22_X1 port map( A1 => A_neg(60), A2 => n155, B1 => A_signal(60), 
                           B2 => n146, ZN => n300);
   U141 : NAND2_X1 port map( A1 => n246, A2 => n245, ZN => Y(36));
   U142 : AOI222_X1 port map( A1 => A_shifted(36), A2 => n179, B1 => 
                           zeroSignal(36), B2 => n170, C1 => A_neg_shifted(36),
                           C2 => n162, ZN => n245);
   U143 : AOI22_X1 port map( A1 => A_neg(36), A2 => n153, B1 => A_signal(36), 
                           B2 => n144, ZN => n246);
   U144 : NAND2_X1 port map( A1 => n248, A2 => n247, ZN => Y(37));
   U145 : AOI222_X1 port map( A1 => A_shifted(37), A2 => n179, B1 => 
                           zeroSignal(37), B2 => n170, C1 => A_neg_shifted(37),
                           C2 => n162, ZN => n247);
   U146 : AOI22_X1 port map( A1 => A_neg(37), A2 => n153, B1 => A_signal(37), 
                           B2 => n144, ZN => n248);
   U147 : NAND2_X1 port map( A1 => n250, A2 => n249, ZN => Y(38));
   U148 : AOI222_X1 port map( A1 => A_shifted(38), A2 => n179, B1 => 
                           zeroSignal(38), B2 => n170, C1 => A_neg_shifted(38),
                           C2 => n162, ZN => n249);
   U149 : AOI22_X1 port map( A1 => A_neg(38), A2 => n153, B1 => A_signal(38), 
                           B2 => n144, ZN => n250);
   U150 : NAND2_X1 port map( A1 => n252, A2 => n251, ZN => Y(39));
   U151 : AOI222_X1 port map( A1 => A_shifted(39), A2 => n179, B1 => 
                           zeroSignal(39), B2 => n170, C1 => A_neg_shifted(39),
                           C2 => n162, ZN => n251);
   U152 : AOI22_X1 port map( A1 => A_neg(39), A2 => n153, B1 => A_signal(39), 
                           B2 => n144, ZN => n252);
   U153 : NAND2_X1 port map( A1 => n188, A2 => n187, ZN => Y(0));
   U154 : AOI22_X1 port map( A1 => A_neg(0), A2 => n151, B1 => A_signal(0), B2 
                           => n142, ZN => n188);
   U155 : AOI222_X1 port map( A1 => A_shifted(0), A2 => n177, B1 => 
                           zeroSignal(0), B2 => n168, C1 => A_neg_shifted(0), 
                           C2 => n165, ZN => n187);
   U156 : NAND2_X1 port map( A1 => n210, A2 => n209, ZN => Y(1));
   U157 : AOI22_X1 port map( A1 => A_neg(1), A2 => n151, B1 => A_signal(1), B2 
                           => n142, ZN => n210);
   U158 : AOI222_X1 port map( A1 => A_shifted(1), A2 => n177, B1 => 
                           zeroSignal(1), B2 => n168, C1 => A_neg_shifted(1), 
                           C2 => n164, ZN => n209);
   U159 : NAND2_X1 port map( A1 => n232, A2 => n231, ZN => Y(2));
   U160 : AOI22_X1 port map( A1 => A_neg(2), A2 => n152, B1 => A_signal(2), B2 
                           => n143, ZN => n232);
   U161 : AOI222_X1 port map( A1 => A_shifted(2), A2 => n178, B1 => 
                           zeroSignal(2), B2 => n169, C1 => A_neg_shifted(2), 
                           C2 => n163, ZN => n231);
   U162 : NAND2_X1 port map( A1 => n254, A2 => n253, ZN => Y(3));
   U163 : AOI22_X1 port map( A1 => A_neg(3), A2 => n153, B1 => A_signal(3), B2 
                           => n144, ZN => n254);
   U164 : AOI222_X1 port map( A1 => A_shifted(3), A2 => n179, B1 => 
                           zeroSignal(3), B2 => n170, C1 => A_neg_shifted(3), 
                           C2 => n162, ZN => n253);
   U165 : NAND2_X1 port map( A1 => n276, A2 => n275, ZN => Y(4));
   U166 : AOI22_X1 port map( A1 => A_neg(4), A2 => n154, B1 => A_signal(4), B2 
                           => n145, ZN => n276);
   U167 : AOI222_X1 port map( A1 => A_shifted(4), A2 => n180, B1 => 
                           zeroSignal(4), B2 => n171, C1 => A_neg_shifted(4), 
                           C2 => n161, ZN => n275);
   U168 : NAND2_X1 port map( A1 => n298, A2 => n297, ZN => Y(5));
   U169 : AOI22_X1 port map( A1 => A_neg(5), A2 => n155, B1 => A_signal(5), B2 
                           => n146, ZN => n298);
   U170 : AOI222_X1 port map( A1 => A_shifted(5), A2 => n181, B1 => 
                           zeroSignal(5), B2 => n172, C1 => A_neg_shifted(5), 
                           C2 => n160, ZN => n297);
   U171 : NAND2_X1 port map( A1 => n308, A2 => n307, ZN => Y(6));
   U172 : AOI22_X1 port map( A1 => A_neg(6), A2 => n156, B1 => A_signal(6), B2 
                           => n147, ZN => n308);
   U173 : AOI222_X1 port map( A1 => A_shifted(6), A2 => n182, B1 => 
                           zeroSignal(6), B2 => n173, C1 => A_neg_shifted(6), 
                           C2 => n160, ZN => n307);
   U174 : NAND2_X1 port map( A1 => n310, A2 => n309, ZN => Y(7));
   U175 : AOI22_X1 port map( A1 => A_neg(7), A2 => n156, B1 => A_signal(7), B2 
                           => n147, ZN => n310);
   U176 : AOI222_X1 port map( A1 => A_shifted(7), A2 => n182, B1 => 
                           zeroSignal(7), B2 => n173, C1 => A_neg_shifted(7), 
                           C2 => n160, ZN => n309);
   U177 : NAND2_X1 port map( A1 => n312, A2 => n311, ZN => Y(8));
   U178 : AOI22_X1 port map( A1 => A_neg(8), A2 => n156, B1 => A_signal(8), B2 
                           => n147, ZN => n312);
   U179 : AOI222_X1 port map( A1 => A_shifted(8), A2 => n182, B1 => 
                           zeroSignal(8), B2 => n173, C1 => A_neg_shifted(8), 
                           C2 => n160, ZN => n311);
   U180 : NAND2_X1 port map( A1 => n318, A2 => n317, ZN => Y(9));
   U181 : AOI22_X1 port map( A1 => A_neg(9), A2 => n156, B1 => A_signal(9), B2 
                           => n147, ZN => n318);
   U182 : AOI222_X1 port map( A1 => A_shifted(9), A2 => n182, B1 => 
                           zeroSignal(9), B2 => n173, C1 => A_neg_shifted(9), 
                           C2 => n160, ZN => n317);
   U183 : NAND2_X1 port map( A1 => n190, A2 => n189, ZN => Y(10));
   U184 : AOI22_X1 port map( A1 => A_neg(10), A2 => n151, B1 => A_signal(10), 
                           B2 => n142, ZN => n190);
   U185 : AOI222_X1 port map( A1 => A_shifted(10), A2 => n177, B1 => 
                           zeroSignal(10), B2 => n168, C1 => A_neg_shifted(10),
                           C2 => n165, ZN => n189);
   U186 : NAND2_X1 port map( A1 => n192, A2 => n191, ZN => Y(11));
   U187 : AOI22_X1 port map( A1 => A_neg(11), A2 => n151, B1 => A_signal(11), 
                           B2 => n142, ZN => n192);
   U188 : AOI222_X1 port map( A1 => A_shifted(11), A2 => n177, B1 => 
                           zeroSignal(11), B2 => n168, C1 => A_neg_shifted(11),
                           C2 => n165, ZN => n191);
   U189 : NAND2_X1 port map( A1 => n194, A2 => n193, ZN => Y(12));
   U190 : AOI22_X1 port map( A1 => A_neg(12), A2 => n151, B1 => A_signal(12), 
                           B2 => n142, ZN => n194);
   U191 : AOI222_X1 port map( A1 => A_shifted(12), A2 => n177, B1 => 
                           zeroSignal(12), B2 => n168, C1 => A_neg_shifted(12),
                           C2 => n165, ZN => n193);
   U192 : NAND2_X1 port map( A1 => n196, A2 => n195, ZN => Y(13));
   U193 : AOI22_X1 port map( A1 => A_neg(13), A2 => n151, B1 => A_signal(13), 
                           B2 => n142, ZN => n196);
   U194 : AOI222_X1 port map( A1 => A_shifted(13), A2 => n177, B1 => 
                           zeroSignal(13), B2 => n168, C1 => A_neg_shifted(13),
                           C2 => n164, ZN => n195);
   U195 : NAND2_X1 port map( A1 => n198, A2 => n197, ZN => Y(14));
   U196 : AOI22_X1 port map( A1 => A_neg(14), A2 => n151, B1 => A_signal(14), 
                           B2 => n142, ZN => n198);
   U197 : AOI222_X1 port map( A1 => A_shifted(14), A2 => n177, B1 => 
                           zeroSignal(14), B2 => n168, C1 => A_neg_shifted(14),
                           C2 => n164, ZN => n197);
   U198 : NAND2_X1 port map( A1 => n200, A2 => n199, ZN => Y(15));
   U199 : AOI22_X1 port map( A1 => A_neg(15), A2 => n151, B1 => A_signal(15), 
                           B2 => n142, ZN => n200);
   U200 : AOI222_X1 port map( A1 => A_shifted(15), A2 => n177, B1 => 
                           zeroSignal(15), B2 => n168, C1 => A_neg_shifted(15),
                           C2 => n164, ZN => n199);
   U201 : NAND2_X1 port map( A1 => n202, A2 => n201, ZN => Y(16));
   U202 : AOI22_X1 port map( A1 => A_neg(16), A2 => n151, B1 => A_signal(16), 
                           B2 => n142, ZN => n202);
   U203 : AOI222_X1 port map( A1 => A_shifted(16), A2 => n177, B1 => 
                           zeroSignal(16), B2 => n168, C1 => A_neg_shifted(16),
                           C2 => n164, ZN => n201);
   U204 : NAND2_X1 port map( A1 => n204, A2 => n203, ZN => Y(17));
   U205 : AOI22_X1 port map( A1 => A_neg(17), A2 => n151, B1 => A_signal(17), 
                           B2 => n142, ZN => n204);
   U206 : AOI222_X1 port map( A1 => A_shifted(17), A2 => n177, B1 => 
                           zeroSignal(17), B2 => n168, C1 => A_neg_shifted(17),
                           C2 => n164, ZN => n203);
   U207 : NAND2_X1 port map( A1 => n206, A2 => n205, ZN => Y(18));
   U208 : AOI22_X1 port map( A1 => A_neg(18), A2 => n151, B1 => A_signal(18), 
                           B2 => n142, ZN => n206);
   U209 : AOI222_X1 port map( A1 => A_shifted(18), A2 => n177, B1 => 
                           zeroSignal(18), B2 => n168, C1 => A_neg_shifted(18),
                           C2 => n164, ZN => n205);
   U210 : NAND2_X1 port map( A1 => n208, A2 => n207, ZN => Y(19));
   U211 : AOI22_X1 port map( A1 => A_neg(19), A2 => n151, B1 => A_signal(19), 
                           B2 => n142, ZN => n208);
   U212 : AOI222_X1 port map( A1 => A_shifted(19), A2 => n177, B1 => 
                           zeroSignal(19), B2 => n168, C1 => A_neg_shifted(19),
                           C2 => n164, ZN => n207);
   U213 : NAND2_X1 port map( A1 => n212, A2 => n211, ZN => Y(20));
   U214 : AOI22_X1 port map( A1 => A_neg(20), A2 => n152, B1 => A_signal(20), 
                           B2 => n143, ZN => n212);
   U215 : AOI222_X1 port map( A1 => A_shifted(20), A2 => n178, B1 => 
                           zeroSignal(20), B2 => n169, C1 => A_neg_shifted(20),
                           C2 => n164, ZN => n211);
   U216 : NAND2_X1 port map( A1 => n214, A2 => n213, ZN => Y(21));
   U217 : AOI22_X1 port map( A1 => A_neg(21), A2 => n152, B1 => A_signal(21), 
                           B2 => n143, ZN => n214);
   U218 : AOI222_X1 port map( A1 => A_shifted(21), A2 => n178, B1 => 
                           zeroSignal(21), B2 => n169, C1 => A_neg_shifted(21),
                           C2 => n164, ZN => n213);
   U219 : NAND2_X1 port map( A1 => n216, A2 => n215, ZN => Y(22));
   U220 : AOI22_X1 port map( A1 => A_neg(22), A2 => n152, B1 => A_signal(22), 
                           B2 => n143, ZN => n216);
   U221 : AOI222_X1 port map( A1 => A_shifted(22), A2 => n178, B1 => 
                           zeroSignal(22), B2 => n169, C1 => A_neg_shifted(22),
                           C2 => n164, ZN => n215);
   U222 : NAND2_X1 port map( A1 => n218, A2 => n217, ZN => Y(23));
   U223 : AOI22_X1 port map( A1 => A_neg(23), A2 => n152, B1 => A_signal(23), 
                           B2 => n143, ZN => n218);
   U224 : AOI222_X1 port map( A1 => A_shifted(23), A2 => n178, B1 => 
                           zeroSignal(23), B2 => n169, C1 => A_neg_shifted(23),
                           C2 => n164, ZN => n217);
   U225 : NAND2_X1 port map( A1 => n220, A2 => n219, ZN => Y(24));
   U226 : AOI22_X1 port map( A1 => A_neg(24), A2 => n152, B1 => A_signal(24), 
                           B2 => n143, ZN => n220);
   U227 : AOI222_X1 port map( A1 => A_shifted(24), A2 => n178, B1 => 
                           zeroSignal(24), B2 => n169, C1 => A_neg_shifted(24),
                           C2 => n163, ZN => n219);
   U228 : NAND2_X1 port map( A1 => n222, A2 => n221, ZN => Y(25));
   U229 : AOI22_X1 port map( A1 => A_neg(25), A2 => n152, B1 => A_signal(25), 
                           B2 => n143, ZN => n222);
   U230 : AOI222_X1 port map( A1 => A_shifted(25), A2 => n178, B1 => 
                           zeroSignal(25), B2 => n169, C1 => A_neg_shifted(25),
                           C2 => n163, ZN => n221);
   U231 : NAND2_X1 port map( A1 => n224, A2 => n223, ZN => Y(26));
   U232 : AOI22_X1 port map( A1 => A_neg(26), A2 => n152, B1 => A_signal(26), 
                           B2 => n143, ZN => n224);
   U233 : AOI222_X1 port map( A1 => A_shifted(26), A2 => n178, B1 => 
                           zeroSignal(26), B2 => n169, C1 => A_neg_shifted(26),
                           C2 => n163, ZN => n223);
   U234 : NAND2_X1 port map( A1 => n226, A2 => n225, ZN => Y(27));
   U235 : AOI22_X1 port map( A1 => A_neg(27), A2 => n152, B1 => A_signal(27), 
                           B2 => n143, ZN => n226);
   U236 : AOI222_X1 port map( A1 => A_shifted(27), A2 => n178, B1 => 
                           zeroSignal(27), B2 => n169, C1 => A_neg_shifted(27),
                           C2 => n163, ZN => n225);
   U237 : NAND2_X1 port map( A1 => n228, A2 => n227, ZN => Y(28));
   U238 : AOI22_X1 port map( A1 => A_neg(28), A2 => n152, B1 => A_signal(28), 
                           B2 => n143, ZN => n228);
   U239 : AOI222_X1 port map( A1 => A_shifted(28), A2 => n178, B1 => 
                           zeroSignal(28), B2 => n169, C1 => A_neg_shifted(28),
                           C2 => n163, ZN => n227);
   U240 : NAND2_X1 port map( A1 => n230, A2 => n229, ZN => Y(29));
   U241 : AOI22_X1 port map( A1 => A_neg(29), A2 => n152, B1 => A_signal(29), 
                           B2 => n143, ZN => n230);
   U242 : AOI222_X1 port map( A1 => A_shifted(29), A2 => n178, B1 => 
                           zeroSignal(29), B2 => n169, C1 => A_neg_shifted(29),
                           C2 => n163, ZN => n229);
   U243 : AOI222_X1 port map( A1 => A_shifted(31), A2 => n179, B1 => 
                           zeroSignal(31), B2 => n170, C1 => A_neg_shifted(31),
                           C2 => n163, ZN => n235);
   U244 : AOI22_X1 port map( A1 => A_neg(30), A2 => n152, B1 => A_signal(30), 
                           B2 => n143, ZN => n234);

end SYN_BEHAVIORAL_2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity encoder_31 is

   port( pieceofB : in std_logic_vector (2 downto 0);  sel : out 
         std_logic_vector (2 downto 0));

end encoder_31;

architecture SYN_behavioral of encoder_31 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n9, n10, n11 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => n10, A2 => n7, ZN => n4);
   U4 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => n7);
   U5 : NAND2_X1 port map( A1 => n7, A2 => n10, ZN => n9);
   U6 : INV_X1 port map( A => pieceofB(1), ZN => n5);
   U7 : INV_X1 port map( A => pieceofB(0), ZN => n6);
   U8 : INV_X1 port map( A => pieceofB(2), ZN => n11);
   U9 : NAND2_X1 port map( A1 => pieceofB(1), A2 => pieceofB(0), ZN => n10);
   U10 : AND3_X1 port map( A1 => pieceofB(2), A2 => n10, A3 => n9, ZN => sel(2)
                           );
   U11 : AOI21_X1 port map( B1 => n9, B2 => n10, A => pieceofB(2), ZN => sel(0)
                           );
   U12 : OAI22_X1 port map( A1 => n11, A2 => n4, B1 => pieceofB(2), B2 => n10, 
                           ZN => sel(1));

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity encoder_30 is

   port( pieceofB : in std_logic_vector (2 downto 0);  sel : out 
         std_logic_vector (2 downto 0));

end encoder_30;

architecture SYN_behavioral of encoder_30 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n6, n7 : std_logic;

begin
   
   U3 : INV_X1 port map( A => pieceofB(2), ZN => n7);
   U4 : NAND2_X1 port map( A1 => pieceofB(1), A2 => pieceofB(0), ZN => n6);
   U5 : AOI21_X1 port map( B1 => n5, B2 => n6, A => pieceofB(2), ZN => sel(0));
   U6 : AND3_X1 port map( A1 => pieceofB(2), A2 => n6, A3 => n5, ZN => sel(2));
   U7 : OAI22_X1 port map( A1 => n7, A2 => n5, B1 => pieceofB(2), B2 => n6, ZN 
                           => sel(1));
   U8 : OAI21_X1 port map( B1 => pieceofB(1), B2 => pieceofB(0), A => n6, ZN =>
                           n5);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity encoder_29 is

   port( pieceofB : in std_logic_vector (2 downto 0);  sel : out 
         std_logic_vector (2 downto 0));

end encoder_29;

architecture SYN_behavioral of encoder_29 is

   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n6, n7 : std_logic;

begin
   
   U3 : OAI22_X1 port map( A1 => n7, A2 => n5, B1 => pieceofB(2), B2 => n6, ZN 
                           => sel(1));
   U4 : INV_X1 port map( A => pieceofB(2), ZN => n7);
   U5 : OAI21_X1 port map( B1 => pieceofB(1), B2 => pieceofB(0), A => n6, ZN =>
                           n5);
   U6 : NAND2_X1 port map( A1 => pieceofB(1), A2 => pieceofB(0), ZN => n6);
   U7 : AOI21_X1 port map( B1 => n5, B2 => n6, A => pieceofB(2), ZN => sel(0));
   U8 : AND3_X1 port map( A1 => pieceofB(2), A2 => n6, A3 => n5, ZN => sel(2));

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity encoder_28 is

   port( pieceofB : in std_logic_vector (2 downto 0);  sel : out 
         std_logic_vector (2 downto 0));

end encoder_28;

architecture SYN_behavioral of encoder_28 is

   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n6, n7 : std_logic;

begin
   
   U3 : OAI22_X1 port map( A1 => n7, A2 => n5, B1 => pieceofB(2), B2 => n6, ZN 
                           => sel(1));
   U4 : INV_X1 port map( A => pieceofB(2), ZN => n7);
   U5 : OAI21_X1 port map( B1 => pieceofB(1), B2 => pieceofB(0), A => n6, ZN =>
                           n5);
   U6 : NAND2_X1 port map( A1 => pieceofB(1), A2 => pieceofB(0), ZN => n6);
   U7 : AOI21_X1 port map( B1 => n5, B2 => n6, A => pieceofB(2), ZN => sel(0));
   U8 : AND3_X1 port map( A1 => pieceofB(2), A2 => n6, A3 => n5, ZN => sel(2));

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity encoder_27 is

   port( pieceofB : in std_logic_vector (2 downto 0);  sel : out 
         std_logic_vector (2 downto 0));

end encoder_27;

architecture SYN_behavioral of encoder_27 is

   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n6, n7 : std_logic;

begin
   
   U3 : OAI22_X1 port map( A1 => n7, A2 => n5, B1 => pieceofB(2), B2 => n6, ZN 
                           => sel(1));
   U4 : INV_X1 port map( A => pieceofB(2), ZN => n7);
   U5 : OAI21_X1 port map( B1 => pieceofB(1), B2 => pieceofB(0), A => n6, ZN =>
                           n5);
   U6 : NAND2_X1 port map( A1 => pieceofB(1), A2 => pieceofB(0), ZN => n6);
   U7 : AOI21_X1 port map( B1 => n5, B2 => n6, A => pieceofB(2), ZN => sel(0));
   U8 : AND3_X1 port map( A1 => pieceofB(2), A2 => n6, A3 => n5, ZN => sel(2));

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity encoder_26 is

   port( pieceofB : in std_logic_vector (2 downto 0);  sel : out 
         std_logic_vector (2 downto 0));

end encoder_26;

architecture SYN_behavioral of encoder_26 is

   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n6, n7 : std_logic;

begin
   
   U3 : OAI22_X1 port map( A1 => n7, A2 => n5, B1 => pieceofB(2), B2 => n6, ZN 
                           => sel(1));
   U4 : INV_X1 port map( A => pieceofB(2), ZN => n7);
   U5 : OAI21_X1 port map( B1 => pieceofB(1), B2 => pieceofB(0), A => n6, ZN =>
                           n5);
   U6 : NAND2_X1 port map( A1 => pieceofB(1), A2 => pieceofB(0), ZN => n6);
   U7 : AOI21_X1 port map( B1 => n5, B2 => n6, A => pieceofB(2), ZN => sel(0));
   U8 : AND3_X1 port map( A1 => pieceofB(2), A2 => n6, A3 => n5, ZN => sel(2));

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity encoder_25 is

   port( pieceofB : in std_logic_vector (2 downto 0);  sel : out 
         std_logic_vector (2 downto 0));

end encoder_25;

architecture SYN_behavioral of encoder_25 is

   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n6, n7 : std_logic;

begin
   
   U3 : OAI22_X1 port map( A1 => n7, A2 => n5, B1 => pieceofB(2), B2 => n6, ZN 
                           => sel(1));
   U4 : INV_X1 port map( A => pieceofB(2), ZN => n7);
   U5 : OAI21_X1 port map( B1 => pieceofB(1), B2 => pieceofB(0), A => n6, ZN =>
                           n5);
   U6 : NAND2_X1 port map( A1 => pieceofB(1), A2 => pieceofB(0), ZN => n6);
   U7 : AOI21_X1 port map( B1 => n5, B2 => n6, A => pieceofB(2), ZN => sel(0));
   U8 : AND3_X1 port map( A1 => pieceofB(2), A2 => n6, A3 => n5, ZN => sel(2));

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity encoder_24 is

   port( pieceofB : in std_logic_vector (2 downto 0);  sel : out 
         std_logic_vector (2 downto 0));

end encoder_24;

architecture SYN_behavioral of encoder_24 is

   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n6, n7 : std_logic;

begin
   
   U3 : OAI22_X1 port map( A1 => n7, A2 => n5, B1 => pieceofB(2), B2 => n6, ZN 
                           => sel(1));
   U4 : INV_X1 port map( A => pieceofB(2), ZN => n7);
   U5 : OAI21_X1 port map( B1 => pieceofB(1), B2 => pieceofB(0), A => n6, ZN =>
                           n5);
   U6 : NAND2_X1 port map( A1 => pieceofB(1), A2 => pieceofB(0), ZN => n6);
   U7 : AOI21_X1 port map( B1 => n5, B2 => n6, A => pieceofB(2), ZN => sel(0));
   U8 : AND3_X1 port map( A1 => pieceofB(2), A2 => n6, A3 => n5, ZN => sel(2));

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity encoder_23 is

   port( pieceofB : in std_logic_vector (2 downto 0);  sel : out 
         std_logic_vector (2 downto 0));

end encoder_23;

architecture SYN_behavioral of encoder_23 is

   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n6, n7 : std_logic;

begin
   
   U3 : OAI22_X1 port map( A1 => n7, A2 => n5, B1 => pieceofB(2), B2 => n6, ZN 
                           => sel(1));
   U4 : INV_X1 port map( A => pieceofB(2), ZN => n7);
   U5 : OAI21_X1 port map( B1 => pieceofB(1), B2 => pieceofB(0), A => n6, ZN =>
                           n5);
   U6 : NAND2_X1 port map( A1 => pieceofB(1), A2 => pieceofB(0), ZN => n6);
   U7 : AOI21_X1 port map( B1 => n5, B2 => n6, A => pieceofB(2), ZN => sel(0));
   U8 : AND3_X1 port map( A1 => pieceofB(2), A2 => n6, A3 => n5, ZN => sel(2));

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity encoder_22 is

   port( pieceofB : in std_logic_vector (2 downto 0);  sel : out 
         std_logic_vector (2 downto 0));

end encoder_22;

architecture SYN_behavioral of encoder_22 is

   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n6, n7 : std_logic;

begin
   
   U3 : OAI22_X1 port map( A1 => n7, A2 => n5, B1 => pieceofB(2), B2 => n6, ZN 
                           => sel(1));
   U4 : INV_X1 port map( A => pieceofB(2), ZN => n7);
   U5 : OAI21_X1 port map( B1 => pieceofB(1), B2 => pieceofB(0), A => n6, ZN =>
                           n5);
   U6 : NAND2_X1 port map( A1 => pieceofB(1), A2 => pieceofB(0), ZN => n6);
   U7 : AOI21_X1 port map( B1 => n5, B2 => n6, A => pieceofB(2), ZN => sel(0));
   U8 : AND3_X1 port map( A1 => pieceofB(2), A2 => n6, A3 => n5, ZN => sel(2));

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity encoder_21 is

   port( pieceofB : in std_logic_vector (2 downto 0);  sel : out 
         std_logic_vector (2 downto 0));

end encoder_21;

architecture SYN_behavioral of encoder_21 is

   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n6, n7 : std_logic;

begin
   
   U3 : OAI22_X1 port map( A1 => n7, A2 => n5, B1 => pieceofB(2), B2 => n6, ZN 
                           => sel(1));
   U4 : INV_X1 port map( A => pieceofB(2), ZN => n7);
   U5 : OAI21_X1 port map( B1 => pieceofB(1), B2 => pieceofB(0), A => n6, ZN =>
                           n5);
   U6 : NAND2_X1 port map( A1 => pieceofB(1), A2 => pieceofB(0), ZN => n6);
   U7 : AOI21_X1 port map( B1 => n5, B2 => n6, A => pieceofB(2), ZN => sel(0));
   U8 : AND3_X1 port map( A1 => pieceofB(2), A2 => n6, A3 => n5, ZN => sel(2));

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity encoder_20 is

   port( pieceofB : in std_logic_vector (2 downto 0);  sel : out 
         std_logic_vector (2 downto 0));

end encoder_20;

architecture SYN_behavioral of encoder_20 is

   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n6, n7 : std_logic;

begin
   
   U3 : OAI22_X1 port map( A1 => n7, A2 => n5, B1 => pieceofB(2), B2 => n6, ZN 
                           => sel(1));
   U4 : INV_X1 port map( A => pieceofB(2), ZN => n7);
   U5 : OAI21_X1 port map( B1 => pieceofB(1), B2 => pieceofB(0), A => n6, ZN =>
                           n5);
   U6 : NAND2_X1 port map( A1 => pieceofB(1), A2 => pieceofB(0), ZN => n6);
   U7 : AOI21_X1 port map( B1 => n5, B2 => n6, A => pieceofB(2), ZN => sel(0));
   U8 : AND3_X1 port map( A1 => pieceofB(2), A2 => n6, A3 => n5, ZN => sel(2));

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity encoder_19 is

   port( pieceofB : in std_logic_vector (2 downto 0);  sel : out 
         std_logic_vector (2 downto 0));

end encoder_19;

architecture SYN_behavioral of encoder_19 is

   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n6, n7 : std_logic;

begin
   
   U3 : OAI22_X1 port map( A1 => n7, A2 => n5, B1 => pieceofB(2), B2 => n6, ZN 
                           => sel(1));
   U4 : INV_X1 port map( A => pieceofB(2), ZN => n7);
   U5 : OAI21_X1 port map( B1 => pieceofB(1), B2 => pieceofB(0), A => n6, ZN =>
                           n5);
   U6 : NAND2_X1 port map( A1 => pieceofB(1), A2 => pieceofB(0), ZN => n6);
   U7 : AOI21_X1 port map( B1 => n5, B2 => n6, A => pieceofB(2), ZN => sel(0));
   U8 : AND3_X1 port map( A1 => pieceofB(2), A2 => n6, A3 => n5, ZN => sel(2));

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity encoder_18 is

   port( pieceofB : in std_logic_vector (2 downto 0);  sel : out 
         std_logic_vector (2 downto 0));

end encoder_18;

architecture SYN_behavioral of encoder_18 is

   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n6, n7 : std_logic;

begin
   
   U3 : OAI22_X1 port map( A1 => n7, A2 => n5, B1 => pieceofB(2), B2 => n6, ZN 
                           => sel(1));
   U4 : INV_X1 port map( A => pieceofB(2), ZN => n7);
   U5 : OAI21_X1 port map( B1 => pieceofB(1), B2 => pieceofB(0), A => n6, ZN =>
                           n5);
   U6 : NAND2_X1 port map( A1 => pieceofB(1), A2 => pieceofB(0), ZN => n6);
   U7 : AOI21_X1 port map( B1 => n5, B2 => n6, A => pieceofB(2), ZN => sel(0));
   U8 : AND3_X1 port map( A1 => pieceofB(2), A2 => n6, A3 => n5, ZN => sel(2));

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity encoder_17 is

   port( pieceofB : in std_logic_vector (2 downto 0);  sel : out 
         std_logic_vector (2 downto 0));

end encoder_17;

architecture SYN_behavioral of encoder_17 is

   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n6, n7 : std_logic;

begin
   
   U3 : OAI22_X1 port map( A1 => n7, A2 => n5, B1 => pieceofB(2), B2 => n6, ZN 
                           => sel(1));
   U4 : INV_X1 port map( A => pieceofB(2), ZN => n7);
   U5 : OAI21_X1 port map( B1 => pieceofB(1), B2 => pieceofB(0), A => n6, ZN =>
                           n5);
   U6 : NAND2_X1 port map( A1 => pieceofB(1), A2 => pieceofB(0), ZN => n6);
   U7 : AOI21_X1 port map( B1 => n5, B2 => n6, A => pieceofB(2), ZN => sel(0));
   U8 : AND3_X1 port map( A1 => pieceofB(2), A2 => n6, A3 => n5, ZN => sel(2));

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity leftshifter_NbitShifter64_125 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_125;

architecture SYN_behavioral of leftshifter_NbitShifter64_125 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity leftshifter_NbitShifter64_124 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_124;

architecture SYN_behavioral of leftshifter_NbitShifter64_124 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity leftshifter_NbitShifter64_123 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_123;

architecture SYN_behavioral of leftshifter_NbitShifter64_123 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity leftshifter_NbitShifter64_122 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_122;

architecture SYN_behavioral of leftshifter_NbitShifter64_122 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity leftshifter_NbitShifter64_121 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_121;

architecture SYN_behavioral of leftshifter_NbitShifter64_121 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity leftshifter_NbitShifter64_120 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_120;

architecture SYN_behavioral of leftshifter_NbitShifter64_120 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity leftshifter_NbitShifter64_119 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_119;

architecture SYN_behavioral of leftshifter_NbitShifter64_119 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity leftshifter_NbitShifter64_118 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_118;

architecture SYN_behavioral of leftshifter_NbitShifter64_118 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity leftshifter_NbitShifter64_117 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_117;

architecture SYN_behavioral of leftshifter_NbitShifter64_117 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity leftshifter_NbitShifter64_116 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_116;

architecture SYN_behavioral of leftshifter_NbitShifter64_116 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity leftshifter_NbitShifter64_115 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_115;

architecture SYN_behavioral of leftshifter_NbitShifter64_115 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity leftshifter_NbitShifter64_114 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_114;

architecture SYN_behavioral of leftshifter_NbitShifter64_114 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity leftshifter_NbitShifter64_113 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_113;

architecture SYN_behavioral of leftshifter_NbitShifter64_113 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity leftshifter_NbitShifter64_112 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_112;

architecture SYN_behavioral of leftshifter_NbitShifter64_112 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity leftshifter_NbitShifter64_111 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_111;

architecture SYN_behavioral of leftshifter_NbitShifter64_111 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity leftshifter_NbitShifter64_110 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_110;

architecture SYN_behavioral of leftshifter_NbitShifter64_110 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity leftshifter_NbitShifter64_109 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_109;

architecture SYN_behavioral of leftshifter_NbitShifter64_109 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity leftshifter_NbitShifter64_108 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_108;

architecture SYN_behavioral of leftshifter_NbitShifter64_108 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity leftshifter_NbitShifter64_107 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_107;

architecture SYN_behavioral of leftshifter_NbitShifter64_107 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity leftshifter_NbitShifter64_106 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_106;

architecture SYN_behavioral of leftshifter_NbitShifter64_106 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity leftshifter_NbitShifter64_105 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_105;

architecture SYN_behavioral of leftshifter_NbitShifter64_105 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity leftshifter_NbitShifter64_104 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_104;

architecture SYN_behavioral of leftshifter_NbitShifter64_104 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity leftshifter_NbitShifter64_103 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_103;

architecture SYN_behavioral of leftshifter_NbitShifter64_103 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity leftshifter_NbitShifter64_102 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_102;

architecture SYN_behavioral of leftshifter_NbitShifter64_102 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity leftshifter_NbitShifter64_101 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_101;

architecture SYN_behavioral of leftshifter_NbitShifter64_101 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity leftshifter_NbitShifter64_100 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_100;

architecture SYN_behavioral of leftshifter_NbitShifter64_100 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity leftshifter_NbitShifter64_99 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_99;

architecture SYN_behavioral of leftshifter_NbitShifter64_99 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity leftshifter_NbitShifter64_98 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_98;

architecture SYN_behavioral of leftshifter_NbitShifter64_98 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity leftshifter_NbitShifter64_97 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_97;

architecture SYN_behavioral of leftshifter_NbitShifter64_97 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity leftshifter_NbitShifter64_96 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_96;

architecture SYN_behavioral of leftshifter_NbitShifter64_96 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity leftshifter_NbitShifter64_95 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_95;

architecture SYN_behavioral of leftshifter_NbitShifter64_95 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity leftshifter_NbitShifter64_94 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_94;

architecture SYN_behavioral of leftshifter_NbitShifter64_94 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity leftshifter_NbitShifter64_93 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_93;

architecture SYN_behavioral of leftshifter_NbitShifter64_93 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity leftshifter_NbitShifter64_92 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_92;

architecture SYN_behavioral of leftshifter_NbitShifter64_92 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity leftshifter_NbitShifter64_91 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_91;

architecture SYN_behavioral of leftshifter_NbitShifter64_91 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity leftshifter_NbitShifter64_90 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_90;

architecture SYN_behavioral of leftshifter_NbitShifter64_90 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity leftshifter_NbitShifter64_89 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_89;

architecture SYN_behavioral of leftshifter_NbitShifter64_89 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity leftshifter_NbitShifter64_88 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_88;

architecture SYN_behavioral of leftshifter_NbitShifter64_88 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity leftshifter_NbitShifter64_87 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_87;

architecture SYN_behavioral of leftshifter_NbitShifter64_87 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity leftshifter_NbitShifter64_86 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_86;

architecture SYN_behavioral of leftshifter_NbitShifter64_86 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity leftshifter_NbitShifter64_85 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_85;

architecture SYN_behavioral of leftshifter_NbitShifter64_85 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity leftshifter_NbitShifter64_84 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_84;

architecture SYN_behavioral of leftshifter_NbitShifter64_84 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity leftshifter_NbitShifter64_83 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_83;

architecture SYN_behavioral of leftshifter_NbitShifter64_83 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity leftshifter_NbitShifter64_82 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_82;

architecture SYN_behavioral of leftshifter_NbitShifter64_82 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity leftshifter_NbitShifter64_81 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_81;

architecture SYN_behavioral of leftshifter_NbitShifter64_81 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity leftshifter_NbitShifter64_80 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_80;

architecture SYN_behavioral of leftshifter_NbitShifter64_80 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity leftshifter_NbitShifter64_79 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_79;

architecture SYN_behavioral of leftshifter_NbitShifter64_79 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity leftshifter_NbitShifter64_78 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_78;

architecture SYN_behavioral of leftshifter_NbitShifter64_78 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity leftshifter_NbitShifter64_77 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_77;

architecture SYN_behavioral of leftshifter_NbitShifter64_77 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity leftshifter_NbitShifter64_76 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_76;

architecture SYN_behavioral of leftshifter_NbitShifter64_76 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity leftshifter_NbitShifter64_75 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_75;

architecture SYN_behavioral of leftshifter_NbitShifter64_75 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity leftshifter_NbitShifter64_74 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_74;

architecture SYN_behavioral of leftshifter_NbitShifter64_74 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity leftshifter_NbitShifter64_73 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_73;

architecture SYN_behavioral of leftshifter_NbitShifter64_73 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity leftshifter_NbitShifter64_72 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_72;

architecture SYN_behavioral of leftshifter_NbitShifter64_72 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity leftshifter_NbitShifter64_71 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_71;

architecture SYN_behavioral of leftshifter_NbitShifter64_71 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity leftshifter_NbitShifter64_70 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_70;

architecture SYN_behavioral of leftshifter_NbitShifter64_70 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity leftshifter_NbitShifter64_69 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_69;

architecture SYN_behavioral of leftshifter_NbitShifter64_69 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity leftshifter_NbitShifter64_68 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_68;

architecture SYN_behavioral of leftshifter_NbitShifter64_68 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity leftshifter_NbitShifter64_67 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_67;

architecture SYN_behavioral of leftshifter_NbitShifter64_67 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity leftshifter_NbitShifter64_66 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_66;

architecture SYN_behavioral of leftshifter_NbitShifter64_66 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity leftshifter_NbitShifter64_65 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_65;

architecture SYN_behavioral of leftshifter_NbitShifter64_65 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity leftshifter_NbitShifter64_64 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_64;

architecture SYN_behavioral of leftshifter_NbitShifter64_64 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity RCA_NbitRca64_30 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_NbitRca64_30;

architecture SYN_STRUCTURAL of RCA_NbitRca64_30 is

   component FA_1857
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1858
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1859
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1860
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1861
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1862
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1863
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1864
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1865
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1866
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1867
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1868
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1869
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1870
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1871
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1872
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1873
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1874
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1875
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1876
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1877
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1878
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1879
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1880
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1881
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1882
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1883
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1884
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1885
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1886
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1887
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1888
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1889
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1890
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1891
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1892
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1893
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1894
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1895
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1896
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1897
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1898
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1899
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1900
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1901
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1902
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1903
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1904
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1905
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1906
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1907
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1908
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1909
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1910
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1911
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1912
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1913
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1914
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1915
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1916
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1917
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1918
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1919
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1920
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_63_port, CTMP_62_port, CTMP_61_port, CTMP_60_port, CTMP_59_port,
      CTMP_58_port, CTMP_57_port, CTMP_56_port, CTMP_55_port, CTMP_54_port, 
      CTMP_53_port, CTMP_52_port, CTMP_51_port, CTMP_50_port, CTMP_49_port, 
      CTMP_48_port, CTMP_47_port, CTMP_46_port, CTMP_45_port, CTMP_44_port, 
      CTMP_43_port, CTMP_42_port, CTMP_41_port, CTMP_40_port, CTMP_39_port, 
      CTMP_38_port, CTMP_37_port, CTMP_36_port, CTMP_35_port, CTMP_34_port, 
      CTMP_33_port, CTMP_32_port, CTMP_31_port, CTMP_30_port, CTMP_29_port, 
      CTMP_28_port, CTMP_27_port, CTMP_26_port, CTMP_25_port, CTMP_24_port, 
      CTMP_23_port, CTMP_22_port, CTMP_21_port, CTMP_20_port, CTMP_19_port, 
      CTMP_18_port, CTMP_17_port, CTMP_16_port, CTMP_15_port, CTMP_14_port, 
      CTMP_13_port, CTMP_12_port, CTMP_11_port, CTMP_10_port, CTMP_9_port, 
      CTMP_8_port, CTMP_7_port, CTMP_6_port, CTMP_5_port, CTMP_4_port, 
      CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_1920 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_1919 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1)
                           , Co => CTMP_2_port);
   FAI_3 : FA_1918 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2)
                           , Co => CTMP_3_port);
   FAI_4 : FA_1917 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3)
                           , Co => CTMP_4_port);
   FAI_5 : FA_1916 port map( A => A(4), B => B(4), Ci => CTMP_4_port, S => S(4)
                           , Co => CTMP_5_port);
   FAI_6 : FA_1915 port map( A => A(5), B => B(5), Ci => CTMP_5_port, S => S(5)
                           , Co => CTMP_6_port);
   FAI_7 : FA_1914 port map( A => A(6), B => B(6), Ci => CTMP_6_port, S => S(6)
                           , Co => CTMP_7_port);
   FAI_8 : FA_1913 port map( A => A(7), B => B(7), Ci => CTMP_7_port, S => S(7)
                           , Co => CTMP_8_port);
   FAI_9 : FA_1912 port map( A => A(8), B => B(8), Ci => CTMP_8_port, S => S(8)
                           , Co => CTMP_9_port);
   FAI_10 : FA_1911 port map( A => A(9), B => B(9), Ci => CTMP_9_port, S => 
                           S(9), Co => CTMP_10_port);
   FAI_11 : FA_1910 port map( A => A(10), B => B(10), Ci => CTMP_10_port, S => 
                           S(10), Co => CTMP_11_port);
   FAI_12 : FA_1909 port map( A => A(11), B => B(11), Ci => CTMP_11_port, S => 
                           S(11), Co => CTMP_12_port);
   FAI_13 : FA_1908 port map( A => A(12), B => B(12), Ci => CTMP_12_port, S => 
                           S(12), Co => CTMP_13_port);
   FAI_14 : FA_1907 port map( A => A(13), B => B(13), Ci => CTMP_13_port, S => 
                           S(13), Co => CTMP_14_port);
   FAI_15 : FA_1906 port map( A => A(14), B => B(14), Ci => CTMP_14_port, S => 
                           S(14), Co => CTMP_15_port);
   FAI_16 : FA_1905 port map( A => A(15), B => B(15), Ci => CTMP_15_port, S => 
                           S(15), Co => CTMP_16_port);
   FAI_17 : FA_1904 port map( A => A(16), B => B(16), Ci => CTMP_16_port, S => 
                           S(16), Co => CTMP_17_port);
   FAI_18 : FA_1903 port map( A => A(17), B => B(17), Ci => CTMP_17_port, S => 
                           S(17), Co => CTMP_18_port);
   FAI_19 : FA_1902 port map( A => A(18), B => B(18), Ci => CTMP_18_port, S => 
                           S(18), Co => CTMP_19_port);
   FAI_20 : FA_1901 port map( A => A(19), B => B(19), Ci => CTMP_19_port, S => 
                           S(19), Co => CTMP_20_port);
   FAI_21 : FA_1900 port map( A => A(20), B => B(20), Ci => CTMP_20_port, S => 
                           S(20), Co => CTMP_21_port);
   FAI_22 : FA_1899 port map( A => A(21), B => B(21), Ci => CTMP_21_port, S => 
                           S(21), Co => CTMP_22_port);
   FAI_23 : FA_1898 port map( A => A(22), B => B(22), Ci => CTMP_22_port, S => 
                           S(22), Co => CTMP_23_port);
   FAI_24 : FA_1897 port map( A => A(23), B => B(23), Ci => CTMP_23_port, S => 
                           S(23), Co => CTMP_24_port);
   FAI_25 : FA_1896 port map( A => A(24), B => B(24), Ci => CTMP_24_port, S => 
                           S(24), Co => CTMP_25_port);
   FAI_26 : FA_1895 port map( A => A(25), B => B(25), Ci => CTMP_25_port, S => 
                           S(25), Co => CTMP_26_port);
   FAI_27 : FA_1894 port map( A => A(26), B => B(26), Ci => CTMP_26_port, S => 
                           S(26), Co => CTMP_27_port);
   FAI_28 : FA_1893 port map( A => A(27), B => B(27), Ci => CTMP_27_port, S => 
                           S(27), Co => CTMP_28_port);
   FAI_29 : FA_1892 port map( A => A(28), B => B(28), Ci => CTMP_28_port, S => 
                           S(28), Co => CTMP_29_port);
   FAI_30 : FA_1891 port map( A => A(29), B => B(29), Ci => CTMP_29_port, S => 
                           S(29), Co => CTMP_30_port);
   FAI_31 : FA_1890 port map( A => A(30), B => B(30), Ci => CTMP_30_port, S => 
                           S(30), Co => CTMP_31_port);
   FAI_32 : FA_1889 port map( A => A(31), B => B(31), Ci => CTMP_31_port, S => 
                           S(31), Co => CTMP_32_port);
   FAI_33 : FA_1888 port map( A => A(32), B => B(32), Ci => CTMP_32_port, S => 
                           S(32), Co => CTMP_33_port);
   FAI_34 : FA_1887 port map( A => A(33), B => B(33), Ci => CTMP_33_port, S => 
                           S(33), Co => CTMP_34_port);
   FAI_35 : FA_1886 port map( A => A(34), B => B(34), Ci => CTMP_34_port, S => 
                           S(34), Co => CTMP_35_port);
   FAI_36 : FA_1885 port map( A => A(35), B => B(35), Ci => CTMP_35_port, S => 
                           S(35), Co => CTMP_36_port);
   FAI_37 : FA_1884 port map( A => A(36), B => B(36), Ci => CTMP_36_port, S => 
                           S(36), Co => CTMP_37_port);
   FAI_38 : FA_1883 port map( A => A(37), B => B(37), Ci => CTMP_37_port, S => 
                           S(37), Co => CTMP_38_port);
   FAI_39 : FA_1882 port map( A => A(38), B => B(38), Ci => CTMP_38_port, S => 
                           S(38), Co => CTMP_39_port);
   FAI_40 : FA_1881 port map( A => A(39), B => B(39), Ci => CTMP_39_port, S => 
                           S(39), Co => CTMP_40_port);
   FAI_41 : FA_1880 port map( A => A(40), B => B(40), Ci => CTMP_40_port, S => 
                           S(40), Co => CTMP_41_port);
   FAI_42 : FA_1879 port map( A => A(41), B => B(41), Ci => CTMP_41_port, S => 
                           S(41), Co => CTMP_42_port);
   FAI_43 : FA_1878 port map( A => A(42), B => B(42), Ci => CTMP_42_port, S => 
                           S(42), Co => CTMP_43_port);
   FAI_44 : FA_1877 port map( A => A(43), B => B(43), Ci => CTMP_43_port, S => 
                           S(43), Co => CTMP_44_port);
   FAI_45 : FA_1876 port map( A => A(44), B => B(44), Ci => CTMP_44_port, S => 
                           S(44), Co => CTMP_45_port);
   FAI_46 : FA_1875 port map( A => A(45), B => B(45), Ci => CTMP_45_port, S => 
                           S(45), Co => CTMP_46_port);
   FAI_47 : FA_1874 port map( A => A(46), B => B(46), Ci => CTMP_46_port, S => 
                           S(46), Co => CTMP_47_port);
   FAI_48 : FA_1873 port map( A => A(47), B => B(47), Ci => CTMP_47_port, S => 
                           S(47), Co => CTMP_48_port);
   FAI_49 : FA_1872 port map( A => A(48), B => B(48), Ci => CTMP_48_port, S => 
                           S(48), Co => CTMP_49_port);
   FAI_50 : FA_1871 port map( A => A(49), B => B(49), Ci => CTMP_49_port, S => 
                           S(49), Co => CTMP_50_port);
   FAI_51 : FA_1870 port map( A => A(50), B => B(50), Ci => CTMP_50_port, S => 
                           S(50), Co => CTMP_51_port);
   FAI_52 : FA_1869 port map( A => A(51), B => B(51), Ci => CTMP_51_port, S => 
                           S(51), Co => CTMP_52_port);
   FAI_53 : FA_1868 port map( A => A(52), B => B(52), Ci => CTMP_52_port, S => 
                           S(52), Co => CTMP_53_port);
   FAI_54 : FA_1867 port map( A => A(53), B => B(53), Ci => CTMP_53_port, S => 
                           S(53), Co => CTMP_54_port);
   FAI_55 : FA_1866 port map( A => A(54), B => B(54), Ci => CTMP_54_port, S => 
                           S(54), Co => CTMP_55_port);
   FAI_56 : FA_1865 port map( A => A(55), B => B(55), Ci => CTMP_55_port, S => 
                           S(55), Co => CTMP_56_port);
   FAI_57 : FA_1864 port map( A => A(56), B => B(56), Ci => CTMP_56_port, S => 
                           S(56), Co => CTMP_57_port);
   FAI_58 : FA_1863 port map( A => A(57), B => B(57), Ci => CTMP_57_port, S => 
                           S(57), Co => CTMP_58_port);
   FAI_59 : FA_1862 port map( A => A(58), B => B(58), Ci => CTMP_58_port, S => 
                           S(58), Co => CTMP_59_port);
   FAI_60 : FA_1861 port map( A => A(59), B => B(59), Ci => CTMP_59_port, S => 
                           S(59), Co => CTMP_60_port);
   FAI_61 : FA_1860 port map( A => A(60), B => B(60), Ci => CTMP_60_port, S => 
                           S(60), Co => CTMP_61_port);
   FAI_62 : FA_1859 port map( A => A(61), B => B(61), Ci => CTMP_61_port, S => 
                           S(61), Co => CTMP_62_port);
   FAI_63 : FA_1858 port map( A => A(62), B => B(62), Ci => CTMP_62_port, S => 
                           S(62), Co => CTMP_63_port);
   FAI_64 : FA_1857 port map( A => A(63), B => B(63), Ci => CTMP_63_port, S => 
                           S(63), Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity RCA_NbitRca64_29 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_NbitRca64_29;

architecture SYN_STRUCTURAL of RCA_NbitRca64_29 is

   component FA_1793
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1794
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1795
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1796
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1797
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1798
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1799
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1800
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1801
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1802
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1803
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1804
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1805
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1806
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1807
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1808
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1809
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1810
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1811
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1812
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1813
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1814
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1815
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1816
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1817
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1818
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1819
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1820
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1821
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1822
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1823
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1824
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1825
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1826
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1827
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1828
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1829
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1830
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1831
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1832
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1833
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1834
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1835
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1836
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1837
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1838
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1839
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1840
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1841
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1842
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1843
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1844
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1845
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1846
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1847
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1848
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1849
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1850
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1851
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1852
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1853
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1854
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1855
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1856
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_63_port, CTMP_62_port, CTMP_61_port, CTMP_60_port, CTMP_59_port,
      CTMP_58_port, CTMP_57_port, CTMP_56_port, CTMP_55_port, CTMP_54_port, 
      CTMP_53_port, CTMP_52_port, CTMP_51_port, CTMP_50_port, CTMP_49_port, 
      CTMP_48_port, CTMP_47_port, CTMP_46_port, CTMP_45_port, CTMP_44_port, 
      CTMP_43_port, CTMP_42_port, CTMP_41_port, CTMP_40_port, CTMP_39_port, 
      CTMP_38_port, CTMP_37_port, CTMP_36_port, CTMP_35_port, CTMP_34_port, 
      CTMP_33_port, CTMP_32_port, CTMP_31_port, CTMP_30_port, CTMP_29_port, 
      CTMP_28_port, CTMP_27_port, CTMP_26_port, CTMP_25_port, CTMP_24_port, 
      CTMP_23_port, CTMP_22_port, CTMP_21_port, CTMP_20_port, CTMP_19_port, 
      CTMP_18_port, CTMP_17_port, CTMP_16_port, CTMP_15_port, CTMP_14_port, 
      CTMP_13_port, CTMP_12_port, CTMP_11_port, CTMP_10_port, CTMP_9_port, 
      CTMP_8_port, CTMP_7_port, CTMP_6_port, CTMP_5_port, CTMP_4_port, 
      CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_1856 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_1855 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1)
                           , Co => CTMP_2_port);
   FAI_3 : FA_1854 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2)
                           , Co => CTMP_3_port);
   FAI_4 : FA_1853 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3)
                           , Co => CTMP_4_port);
   FAI_5 : FA_1852 port map( A => A(4), B => B(4), Ci => CTMP_4_port, S => S(4)
                           , Co => CTMP_5_port);
   FAI_6 : FA_1851 port map( A => A(5), B => B(5), Ci => CTMP_5_port, S => S(5)
                           , Co => CTMP_6_port);
   FAI_7 : FA_1850 port map( A => A(6), B => B(6), Ci => CTMP_6_port, S => S(6)
                           , Co => CTMP_7_port);
   FAI_8 : FA_1849 port map( A => A(7), B => B(7), Ci => CTMP_7_port, S => S(7)
                           , Co => CTMP_8_port);
   FAI_9 : FA_1848 port map( A => A(8), B => B(8), Ci => CTMP_8_port, S => S(8)
                           , Co => CTMP_9_port);
   FAI_10 : FA_1847 port map( A => A(9), B => B(9), Ci => CTMP_9_port, S => 
                           S(9), Co => CTMP_10_port);
   FAI_11 : FA_1846 port map( A => A(10), B => B(10), Ci => CTMP_10_port, S => 
                           S(10), Co => CTMP_11_port);
   FAI_12 : FA_1845 port map( A => A(11), B => B(11), Ci => CTMP_11_port, S => 
                           S(11), Co => CTMP_12_port);
   FAI_13 : FA_1844 port map( A => A(12), B => B(12), Ci => CTMP_12_port, S => 
                           S(12), Co => CTMP_13_port);
   FAI_14 : FA_1843 port map( A => A(13), B => B(13), Ci => CTMP_13_port, S => 
                           S(13), Co => CTMP_14_port);
   FAI_15 : FA_1842 port map( A => A(14), B => B(14), Ci => CTMP_14_port, S => 
                           S(14), Co => CTMP_15_port);
   FAI_16 : FA_1841 port map( A => A(15), B => B(15), Ci => CTMP_15_port, S => 
                           S(15), Co => CTMP_16_port);
   FAI_17 : FA_1840 port map( A => A(16), B => B(16), Ci => CTMP_16_port, S => 
                           S(16), Co => CTMP_17_port);
   FAI_18 : FA_1839 port map( A => A(17), B => B(17), Ci => CTMP_17_port, S => 
                           S(17), Co => CTMP_18_port);
   FAI_19 : FA_1838 port map( A => A(18), B => B(18), Ci => CTMP_18_port, S => 
                           S(18), Co => CTMP_19_port);
   FAI_20 : FA_1837 port map( A => A(19), B => B(19), Ci => CTMP_19_port, S => 
                           S(19), Co => CTMP_20_port);
   FAI_21 : FA_1836 port map( A => A(20), B => B(20), Ci => CTMP_20_port, S => 
                           S(20), Co => CTMP_21_port);
   FAI_22 : FA_1835 port map( A => A(21), B => B(21), Ci => CTMP_21_port, S => 
                           S(21), Co => CTMP_22_port);
   FAI_23 : FA_1834 port map( A => A(22), B => B(22), Ci => CTMP_22_port, S => 
                           S(22), Co => CTMP_23_port);
   FAI_24 : FA_1833 port map( A => A(23), B => B(23), Ci => CTMP_23_port, S => 
                           S(23), Co => CTMP_24_port);
   FAI_25 : FA_1832 port map( A => A(24), B => B(24), Ci => CTMP_24_port, S => 
                           S(24), Co => CTMP_25_port);
   FAI_26 : FA_1831 port map( A => A(25), B => B(25), Ci => CTMP_25_port, S => 
                           S(25), Co => CTMP_26_port);
   FAI_27 : FA_1830 port map( A => A(26), B => B(26), Ci => CTMP_26_port, S => 
                           S(26), Co => CTMP_27_port);
   FAI_28 : FA_1829 port map( A => A(27), B => B(27), Ci => CTMP_27_port, S => 
                           S(27), Co => CTMP_28_port);
   FAI_29 : FA_1828 port map( A => A(28), B => B(28), Ci => CTMP_28_port, S => 
                           S(28), Co => CTMP_29_port);
   FAI_30 : FA_1827 port map( A => A(29), B => B(29), Ci => CTMP_29_port, S => 
                           S(29), Co => CTMP_30_port);
   FAI_31 : FA_1826 port map( A => A(30), B => B(30), Ci => CTMP_30_port, S => 
                           S(30), Co => CTMP_31_port);
   FAI_32 : FA_1825 port map( A => A(31), B => B(31), Ci => CTMP_31_port, S => 
                           S(31), Co => CTMP_32_port);
   FAI_33 : FA_1824 port map( A => A(32), B => B(32), Ci => CTMP_32_port, S => 
                           S(32), Co => CTMP_33_port);
   FAI_34 : FA_1823 port map( A => A(33), B => B(33), Ci => CTMP_33_port, S => 
                           S(33), Co => CTMP_34_port);
   FAI_35 : FA_1822 port map( A => A(34), B => B(34), Ci => CTMP_34_port, S => 
                           S(34), Co => CTMP_35_port);
   FAI_36 : FA_1821 port map( A => A(35), B => B(35), Ci => CTMP_35_port, S => 
                           S(35), Co => CTMP_36_port);
   FAI_37 : FA_1820 port map( A => A(36), B => B(36), Ci => CTMP_36_port, S => 
                           S(36), Co => CTMP_37_port);
   FAI_38 : FA_1819 port map( A => A(37), B => B(37), Ci => CTMP_37_port, S => 
                           S(37), Co => CTMP_38_port);
   FAI_39 : FA_1818 port map( A => A(38), B => B(38), Ci => CTMP_38_port, S => 
                           S(38), Co => CTMP_39_port);
   FAI_40 : FA_1817 port map( A => A(39), B => B(39), Ci => CTMP_39_port, S => 
                           S(39), Co => CTMP_40_port);
   FAI_41 : FA_1816 port map( A => A(40), B => B(40), Ci => CTMP_40_port, S => 
                           S(40), Co => CTMP_41_port);
   FAI_42 : FA_1815 port map( A => A(41), B => B(41), Ci => CTMP_41_port, S => 
                           S(41), Co => CTMP_42_port);
   FAI_43 : FA_1814 port map( A => A(42), B => B(42), Ci => CTMP_42_port, S => 
                           S(42), Co => CTMP_43_port);
   FAI_44 : FA_1813 port map( A => A(43), B => B(43), Ci => CTMP_43_port, S => 
                           S(43), Co => CTMP_44_port);
   FAI_45 : FA_1812 port map( A => A(44), B => B(44), Ci => CTMP_44_port, S => 
                           S(44), Co => CTMP_45_port);
   FAI_46 : FA_1811 port map( A => A(45), B => B(45), Ci => CTMP_45_port, S => 
                           S(45), Co => CTMP_46_port);
   FAI_47 : FA_1810 port map( A => A(46), B => B(46), Ci => CTMP_46_port, S => 
                           S(46), Co => CTMP_47_port);
   FAI_48 : FA_1809 port map( A => A(47), B => B(47), Ci => CTMP_47_port, S => 
                           S(47), Co => CTMP_48_port);
   FAI_49 : FA_1808 port map( A => A(48), B => B(48), Ci => CTMP_48_port, S => 
                           S(48), Co => CTMP_49_port);
   FAI_50 : FA_1807 port map( A => A(49), B => B(49), Ci => CTMP_49_port, S => 
                           S(49), Co => CTMP_50_port);
   FAI_51 : FA_1806 port map( A => A(50), B => B(50), Ci => CTMP_50_port, S => 
                           S(50), Co => CTMP_51_port);
   FAI_52 : FA_1805 port map( A => A(51), B => B(51), Ci => CTMP_51_port, S => 
                           S(51), Co => CTMP_52_port);
   FAI_53 : FA_1804 port map( A => A(52), B => B(52), Ci => CTMP_52_port, S => 
                           S(52), Co => CTMP_53_port);
   FAI_54 : FA_1803 port map( A => A(53), B => B(53), Ci => CTMP_53_port, S => 
                           S(53), Co => CTMP_54_port);
   FAI_55 : FA_1802 port map( A => A(54), B => B(54), Ci => CTMP_54_port, S => 
                           S(54), Co => CTMP_55_port);
   FAI_56 : FA_1801 port map( A => A(55), B => B(55), Ci => CTMP_55_port, S => 
                           S(55), Co => CTMP_56_port);
   FAI_57 : FA_1800 port map( A => A(56), B => B(56), Ci => CTMP_56_port, S => 
                           S(56), Co => CTMP_57_port);
   FAI_58 : FA_1799 port map( A => A(57), B => B(57), Ci => CTMP_57_port, S => 
                           S(57), Co => CTMP_58_port);
   FAI_59 : FA_1798 port map( A => A(58), B => B(58), Ci => CTMP_58_port, S => 
                           S(58), Co => CTMP_59_port);
   FAI_60 : FA_1797 port map( A => A(59), B => B(59), Ci => CTMP_59_port, S => 
                           S(59), Co => CTMP_60_port);
   FAI_61 : FA_1796 port map( A => A(60), B => B(60), Ci => CTMP_60_port, S => 
                           S(60), Co => CTMP_61_port);
   FAI_62 : FA_1795 port map( A => A(61), B => B(61), Ci => CTMP_61_port, S => 
                           S(61), Co => CTMP_62_port);
   FAI_63 : FA_1794 port map( A => A(62), B => B(62), Ci => CTMP_62_port, S => 
                           S(62), Co => CTMP_63_port);
   FAI_64 : FA_1793 port map( A => A(63), B => B(63), Ci => CTMP_63_port, S => 
                           S(63), Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity RCA_NbitRca64_28 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_NbitRca64_28;

architecture SYN_STRUCTURAL of RCA_NbitRca64_28 is

   component FA_1729
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1730
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1731
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1732
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1733
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1734
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1735
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1736
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1737
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1738
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1739
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1740
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1741
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1742
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1743
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1744
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1745
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1746
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1747
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1748
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1749
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1750
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1751
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1752
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1753
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1754
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1755
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1756
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1757
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1758
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1759
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1760
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1761
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1762
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1763
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1764
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1765
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1766
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1767
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1768
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1769
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1770
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1771
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1772
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1773
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1774
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1775
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1776
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1777
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1778
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1779
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1780
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1781
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1782
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1783
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1784
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1785
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1786
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1787
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1788
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1789
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1790
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1791
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1792
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_63_port, CTMP_62_port, CTMP_61_port, CTMP_60_port, CTMP_59_port,
      CTMP_58_port, CTMP_57_port, CTMP_56_port, CTMP_55_port, CTMP_54_port, 
      CTMP_53_port, CTMP_52_port, CTMP_51_port, CTMP_50_port, CTMP_49_port, 
      CTMP_48_port, CTMP_47_port, CTMP_46_port, CTMP_45_port, CTMP_44_port, 
      CTMP_43_port, CTMP_42_port, CTMP_41_port, CTMP_40_port, CTMP_39_port, 
      CTMP_38_port, CTMP_37_port, CTMP_36_port, CTMP_35_port, CTMP_34_port, 
      CTMP_33_port, CTMP_32_port, CTMP_31_port, CTMP_30_port, CTMP_29_port, 
      CTMP_28_port, CTMP_27_port, CTMP_26_port, CTMP_25_port, CTMP_24_port, 
      CTMP_23_port, CTMP_22_port, CTMP_21_port, CTMP_20_port, CTMP_19_port, 
      CTMP_18_port, CTMP_17_port, CTMP_16_port, CTMP_15_port, CTMP_14_port, 
      CTMP_13_port, CTMP_12_port, CTMP_11_port, CTMP_10_port, CTMP_9_port, 
      CTMP_8_port, CTMP_7_port, CTMP_6_port, CTMP_5_port, CTMP_4_port, 
      CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_1792 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_1791 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1)
                           , Co => CTMP_2_port);
   FAI_3 : FA_1790 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2)
                           , Co => CTMP_3_port);
   FAI_4 : FA_1789 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3)
                           , Co => CTMP_4_port);
   FAI_5 : FA_1788 port map( A => A(4), B => B(4), Ci => CTMP_4_port, S => S(4)
                           , Co => CTMP_5_port);
   FAI_6 : FA_1787 port map( A => A(5), B => B(5), Ci => CTMP_5_port, S => S(5)
                           , Co => CTMP_6_port);
   FAI_7 : FA_1786 port map( A => A(6), B => B(6), Ci => CTMP_6_port, S => S(6)
                           , Co => CTMP_7_port);
   FAI_8 : FA_1785 port map( A => A(7), B => B(7), Ci => CTMP_7_port, S => S(7)
                           , Co => CTMP_8_port);
   FAI_9 : FA_1784 port map( A => A(8), B => B(8), Ci => CTMP_8_port, S => S(8)
                           , Co => CTMP_9_port);
   FAI_10 : FA_1783 port map( A => A(9), B => B(9), Ci => CTMP_9_port, S => 
                           S(9), Co => CTMP_10_port);
   FAI_11 : FA_1782 port map( A => A(10), B => B(10), Ci => CTMP_10_port, S => 
                           S(10), Co => CTMP_11_port);
   FAI_12 : FA_1781 port map( A => A(11), B => B(11), Ci => CTMP_11_port, S => 
                           S(11), Co => CTMP_12_port);
   FAI_13 : FA_1780 port map( A => A(12), B => B(12), Ci => CTMP_12_port, S => 
                           S(12), Co => CTMP_13_port);
   FAI_14 : FA_1779 port map( A => A(13), B => B(13), Ci => CTMP_13_port, S => 
                           S(13), Co => CTMP_14_port);
   FAI_15 : FA_1778 port map( A => A(14), B => B(14), Ci => CTMP_14_port, S => 
                           S(14), Co => CTMP_15_port);
   FAI_16 : FA_1777 port map( A => A(15), B => B(15), Ci => CTMP_15_port, S => 
                           S(15), Co => CTMP_16_port);
   FAI_17 : FA_1776 port map( A => A(16), B => B(16), Ci => CTMP_16_port, S => 
                           S(16), Co => CTMP_17_port);
   FAI_18 : FA_1775 port map( A => A(17), B => B(17), Ci => CTMP_17_port, S => 
                           S(17), Co => CTMP_18_port);
   FAI_19 : FA_1774 port map( A => A(18), B => B(18), Ci => CTMP_18_port, S => 
                           S(18), Co => CTMP_19_port);
   FAI_20 : FA_1773 port map( A => A(19), B => B(19), Ci => CTMP_19_port, S => 
                           S(19), Co => CTMP_20_port);
   FAI_21 : FA_1772 port map( A => A(20), B => B(20), Ci => CTMP_20_port, S => 
                           S(20), Co => CTMP_21_port);
   FAI_22 : FA_1771 port map( A => A(21), B => B(21), Ci => CTMP_21_port, S => 
                           S(21), Co => CTMP_22_port);
   FAI_23 : FA_1770 port map( A => A(22), B => B(22), Ci => CTMP_22_port, S => 
                           S(22), Co => CTMP_23_port);
   FAI_24 : FA_1769 port map( A => A(23), B => B(23), Ci => CTMP_23_port, S => 
                           S(23), Co => CTMP_24_port);
   FAI_25 : FA_1768 port map( A => A(24), B => B(24), Ci => CTMP_24_port, S => 
                           S(24), Co => CTMP_25_port);
   FAI_26 : FA_1767 port map( A => A(25), B => B(25), Ci => CTMP_25_port, S => 
                           S(25), Co => CTMP_26_port);
   FAI_27 : FA_1766 port map( A => A(26), B => B(26), Ci => CTMP_26_port, S => 
                           S(26), Co => CTMP_27_port);
   FAI_28 : FA_1765 port map( A => A(27), B => B(27), Ci => CTMP_27_port, S => 
                           S(27), Co => CTMP_28_port);
   FAI_29 : FA_1764 port map( A => A(28), B => B(28), Ci => CTMP_28_port, S => 
                           S(28), Co => CTMP_29_port);
   FAI_30 : FA_1763 port map( A => A(29), B => B(29), Ci => CTMP_29_port, S => 
                           S(29), Co => CTMP_30_port);
   FAI_31 : FA_1762 port map( A => A(30), B => B(30), Ci => CTMP_30_port, S => 
                           S(30), Co => CTMP_31_port);
   FAI_32 : FA_1761 port map( A => A(31), B => B(31), Ci => CTMP_31_port, S => 
                           S(31), Co => CTMP_32_port);
   FAI_33 : FA_1760 port map( A => A(32), B => B(32), Ci => CTMP_32_port, S => 
                           S(32), Co => CTMP_33_port);
   FAI_34 : FA_1759 port map( A => A(33), B => B(33), Ci => CTMP_33_port, S => 
                           S(33), Co => CTMP_34_port);
   FAI_35 : FA_1758 port map( A => A(34), B => B(34), Ci => CTMP_34_port, S => 
                           S(34), Co => CTMP_35_port);
   FAI_36 : FA_1757 port map( A => A(35), B => B(35), Ci => CTMP_35_port, S => 
                           S(35), Co => CTMP_36_port);
   FAI_37 : FA_1756 port map( A => A(36), B => B(36), Ci => CTMP_36_port, S => 
                           S(36), Co => CTMP_37_port);
   FAI_38 : FA_1755 port map( A => A(37), B => B(37), Ci => CTMP_37_port, S => 
                           S(37), Co => CTMP_38_port);
   FAI_39 : FA_1754 port map( A => A(38), B => B(38), Ci => CTMP_38_port, S => 
                           S(38), Co => CTMP_39_port);
   FAI_40 : FA_1753 port map( A => A(39), B => B(39), Ci => CTMP_39_port, S => 
                           S(39), Co => CTMP_40_port);
   FAI_41 : FA_1752 port map( A => A(40), B => B(40), Ci => CTMP_40_port, S => 
                           S(40), Co => CTMP_41_port);
   FAI_42 : FA_1751 port map( A => A(41), B => B(41), Ci => CTMP_41_port, S => 
                           S(41), Co => CTMP_42_port);
   FAI_43 : FA_1750 port map( A => A(42), B => B(42), Ci => CTMP_42_port, S => 
                           S(42), Co => CTMP_43_port);
   FAI_44 : FA_1749 port map( A => A(43), B => B(43), Ci => CTMP_43_port, S => 
                           S(43), Co => CTMP_44_port);
   FAI_45 : FA_1748 port map( A => A(44), B => B(44), Ci => CTMP_44_port, S => 
                           S(44), Co => CTMP_45_port);
   FAI_46 : FA_1747 port map( A => A(45), B => B(45), Ci => CTMP_45_port, S => 
                           S(45), Co => CTMP_46_port);
   FAI_47 : FA_1746 port map( A => A(46), B => B(46), Ci => CTMP_46_port, S => 
                           S(46), Co => CTMP_47_port);
   FAI_48 : FA_1745 port map( A => A(47), B => B(47), Ci => CTMP_47_port, S => 
                           S(47), Co => CTMP_48_port);
   FAI_49 : FA_1744 port map( A => A(48), B => B(48), Ci => CTMP_48_port, S => 
                           S(48), Co => CTMP_49_port);
   FAI_50 : FA_1743 port map( A => A(49), B => B(49), Ci => CTMP_49_port, S => 
                           S(49), Co => CTMP_50_port);
   FAI_51 : FA_1742 port map( A => A(50), B => B(50), Ci => CTMP_50_port, S => 
                           S(50), Co => CTMP_51_port);
   FAI_52 : FA_1741 port map( A => A(51), B => B(51), Ci => CTMP_51_port, S => 
                           S(51), Co => CTMP_52_port);
   FAI_53 : FA_1740 port map( A => A(52), B => B(52), Ci => CTMP_52_port, S => 
                           S(52), Co => CTMP_53_port);
   FAI_54 : FA_1739 port map( A => A(53), B => B(53), Ci => CTMP_53_port, S => 
                           S(53), Co => CTMP_54_port);
   FAI_55 : FA_1738 port map( A => A(54), B => B(54), Ci => CTMP_54_port, S => 
                           S(54), Co => CTMP_55_port);
   FAI_56 : FA_1737 port map( A => A(55), B => B(55), Ci => CTMP_55_port, S => 
                           S(55), Co => CTMP_56_port);
   FAI_57 : FA_1736 port map( A => A(56), B => B(56), Ci => CTMP_56_port, S => 
                           S(56), Co => CTMP_57_port);
   FAI_58 : FA_1735 port map( A => A(57), B => B(57), Ci => CTMP_57_port, S => 
                           S(57), Co => CTMP_58_port);
   FAI_59 : FA_1734 port map( A => A(58), B => B(58), Ci => CTMP_58_port, S => 
                           S(58), Co => CTMP_59_port);
   FAI_60 : FA_1733 port map( A => A(59), B => B(59), Ci => CTMP_59_port, S => 
                           S(59), Co => CTMP_60_port);
   FAI_61 : FA_1732 port map( A => A(60), B => B(60), Ci => CTMP_60_port, S => 
                           S(60), Co => CTMP_61_port);
   FAI_62 : FA_1731 port map( A => A(61), B => B(61), Ci => CTMP_61_port, S => 
                           S(61), Co => CTMP_62_port);
   FAI_63 : FA_1730 port map( A => A(62), B => B(62), Ci => CTMP_62_port, S => 
                           S(62), Co => CTMP_63_port);
   FAI_64 : FA_1729 port map( A => A(63), B => B(63), Ci => CTMP_63_port, S => 
                           S(63), Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity RCA_NbitRca64_27 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_NbitRca64_27;

architecture SYN_STRUCTURAL of RCA_NbitRca64_27 is

   component FA_1665
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1666
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1667
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1668
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1669
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1670
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1671
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1672
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1673
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1674
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1675
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1676
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1677
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1678
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1679
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1680
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1681
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1682
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1683
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1684
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1685
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1686
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1687
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1688
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1689
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1690
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1691
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1692
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1693
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1694
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1695
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1696
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1697
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1698
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1699
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1700
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1701
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1702
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1703
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1704
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1705
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1706
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1707
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1708
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1709
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1710
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1711
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1712
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1713
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1714
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1715
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1716
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1717
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1718
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1719
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1720
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1721
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1722
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1723
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1724
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1725
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1726
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1727
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1728
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_63_port, CTMP_62_port, CTMP_61_port, CTMP_60_port, CTMP_59_port,
      CTMP_58_port, CTMP_57_port, CTMP_56_port, CTMP_55_port, CTMP_54_port, 
      CTMP_53_port, CTMP_52_port, CTMP_51_port, CTMP_50_port, CTMP_49_port, 
      CTMP_48_port, CTMP_47_port, CTMP_46_port, CTMP_45_port, CTMP_44_port, 
      CTMP_43_port, CTMP_42_port, CTMP_41_port, CTMP_40_port, CTMP_39_port, 
      CTMP_38_port, CTMP_37_port, CTMP_36_port, CTMP_35_port, CTMP_34_port, 
      CTMP_33_port, CTMP_32_port, CTMP_31_port, CTMP_30_port, CTMP_29_port, 
      CTMP_28_port, CTMP_27_port, CTMP_26_port, CTMP_25_port, CTMP_24_port, 
      CTMP_23_port, CTMP_22_port, CTMP_21_port, CTMP_20_port, CTMP_19_port, 
      CTMP_18_port, CTMP_17_port, CTMP_16_port, CTMP_15_port, CTMP_14_port, 
      CTMP_13_port, CTMP_12_port, CTMP_11_port, CTMP_10_port, CTMP_9_port, 
      CTMP_8_port, CTMP_7_port, CTMP_6_port, CTMP_5_port, CTMP_4_port, 
      CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_1728 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_1727 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1)
                           , Co => CTMP_2_port);
   FAI_3 : FA_1726 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2)
                           , Co => CTMP_3_port);
   FAI_4 : FA_1725 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3)
                           , Co => CTMP_4_port);
   FAI_5 : FA_1724 port map( A => A(4), B => B(4), Ci => CTMP_4_port, S => S(4)
                           , Co => CTMP_5_port);
   FAI_6 : FA_1723 port map( A => A(5), B => B(5), Ci => CTMP_5_port, S => S(5)
                           , Co => CTMP_6_port);
   FAI_7 : FA_1722 port map( A => A(6), B => B(6), Ci => CTMP_6_port, S => S(6)
                           , Co => CTMP_7_port);
   FAI_8 : FA_1721 port map( A => A(7), B => B(7), Ci => CTMP_7_port, S => S(7)
                           , Co => CTMP_8_port);
   FAI_9 : FA_1720 port map( A => A(8), B => B(8), Ci => CTMP_8_port, S => S(8)
                           , Co => CTMP_9_port);
   FAI_10 : FA_1719 port map( A => A(9), B => B(9), Ci => CTMP_9_port, S => 
                           S(9), Co => CTMP_10_port);
   FAI_11 : FA_1718 port map( A => A(10), B => B(10), Ci => CTMP_10_port, S => 
                           S(10), Co => CTMP_11_port);
   FAI_12 : FA_1717 port map( A => A(11), B => B(11), Ci => CTMP_11_port, S => 
                           S(11), Co => CTMP_12_port);
   FAI_13 : FA_1716 port map( A => A(12), B => B(12), Ci => CTMP_12_port, S => 
                           S(12), Co => CTMP_13_port);
   FAI_14 : FA_1715 port map( A => A(13), B => B(13), Ci => CTMP_13_port, S => 
                           S(13), Co => CTMP_14_port);
   FAI_15 : FA_1714 port map( A => A(14), B => B(14), Ci => CTMP_14_port, S => 
                           S(14), Co => CTMP_15_port);
   FAI_16 : FA_1713 port map( A => A(15), B => B(15), Ci => CTMP_15_port, S => 
                           S(15), Co => CTMP_16_port);
   FAI_17 : FA_1712 port map( A => A(16), B => B(16), Ci => CTMP_16_port, S => 
                           S(16), Co => CTMP_17_port);
   FAI_18 : FA_1711 port map( A => A(17), B => B(17), Ci => CTMP_17_port, S => 
                           S(17), Co => CTMP_18_port);
   FAI_19 : FA_1710 port map( A => A(18), B => B(18), Ci => CTMP_18_port, S => 
                           S(18), Co => CTMP_19_port);
   FAI_20 : FA_1709 port map( A => A(19), B => B(19), Ci => CTMP_19_port, S => 
                           S(19), Co => CTMP_20_port);
   FAI_21 : FA_1708 port map( A => A(20), B => B(20), Ci => CTMP_20_port, S => 
                           S(20), Co => CTMP_21_port);
   FAI_22 : FA_1707 port map( A => A(21), B => B(21), Ci => CTMP_21_port, S => 
                           S(21), Co => CTMP_22_port);
   FAI_23 : FA_1706 port map( A => A(22), B => B(22), Ci => CTMP_22_port, S => 
                           S(22), Co => CTMP_23_port);
   FAI_24 : FA_1705 port map( A => A(23), B => B(23), Ci => CTMP_23_port, S => 
                           S(23), Co => CTMP_24_port);
   FAI_25 : FA_1704 port map( A => A(24), B => B(24), Ci => CTMP_24_port, S => 
                           S(24), Co => CTMP_25_port);
   FAI_26 : FA_1703 port map( A => A(25), B => B(25), Ci => CTMP_25_port, S => 
                           S(25), Co => CTMP_26_port);
   FAI_27 : FA_1702 port map( A => A(26), B => B(26), Ci => CTMP_26_port, S => 
                           S(26), Co => CTMP_27_port);
   FAI_28 : FA_1701 port map( A => A(27), B => B(27), Ci => CTMP_27_port, S => 
                           S(27), Co => CTMP_28_port);
   FAI_29 : FA_1700 port map( A => A(28), B => B(28), Ci => CTMP_28_port, S => 
                           S(28), Co => CTMP_29_port);
   FAI_30 : FA_1699 port map( A => A(29), B => B(29), Ci => CTMP_29_port, S => 
                           S(29), Co => CTMP_30_port);
   FAI_31 : FA_1698 port map( A => A(30), B => B(30), Ci => CTMP_30_port, S => 
                           S(30), Co => CTMP_31_port);
   FAI_32 : FA_1697 port map( A => A(31), B => B(31), Ci => CTMP_31_port, S => 
                           S(31), Co => CTMP_32_port);
   FAI_33 : FA_1696 port map( A => A(32), B => B(32), Ci => CTMP_32_port, S => 
                           S(32), Co => CTMP_33_port);
   FAI_34 : FA_1695 port map( A => A(33), B => B(33), Ci => CTMP_33_port, S => 
                           S(33), Co => CTMP_34_port);
   FAI_35 : FA_1694 port map( A => A(34), B => B(34), Ci => CTMP_34_port, S => 
                           S(34), Co => CTMP_35_port);
   FAI_36 : FA_1693 port map( A => A(35), B => B(35), Ci => CTMP_35_port, S => 
                           S(35), Co => CTMP_36_port);
   FAI_37 : FA_1692 port map( A => A(36), B => B(36), Ci => CTMP_36_port, S => 
                           S(36), Co => CTMP_37_port);
   FAI_38 : FA_1691 port map( A => A(37), B => B(37), Ci => CTMP_37_port, S => 
                           S(37), Co => CTMP_38_port);
   FAI_39 : FA_1690 port map( A => A(38), B => B(38), Ci => CTMP_38_port, S => 
                           S(38), Co => CTMP_39_port);
   FAI_40 : FA_1689 port map( A => A(39), B => B(39), Ci => CTMP_39_port, S => 
                           S(39), Co => CTMP_40_port);
   FAI_41 : FA_1688 port map( A => A(40), B => B(40), Ci => CTMP_40_port, S => 
                           S(40), Co => CTMP_41_port);
   FAI_42 : FA_1687 port map( A => A(41), B => B(41), Ci => CTMP_41_port, S => 
                           S(41), Co => CTMP_42_port);
   FAI_43 : FA_1686 port map( A => A(42), B => B(42), Ci => CTMP_42_port, S => 
                           S(42), Co => CTMP_43_port);
   FAI_44 : FA_1685 port map( A => A(43), B => B(43), Ci => CTMP_43_port, S => 
                           S(43), Co => CTMP_44_port);
   FAI_45 : FA_1684 port map( A => A(44), B => B(44), Ci => CTMP_44_port, S => 
                           S(44), Co => CTMP_45_port);
   FAI_46 : FA_1683 port map( A => A(45), B => B(45), Ci => CTMP_45_port, S => 
                           S(45), Co => CTMP_46_port);
   FAI_47 : FA_1682 port map( A => A(46), B => B(46), Ci => CTMP_46_port, S => 
                           S(46), Co => CTMP_47_port);
   FAI_48 : FA_1681 port map( A => A(47), B => B(47), Ci => CTMP_47_port, S => 
                           S(47), Co => CTMP_48_port);
   FAI_49 : FA_1680 port map( A => A(48), B => B(48), Ci => CTMP_48_port, S => 
                           S(48), Co => CTMP_49_port);
   FAI_50 : FA_1679 port map( A => A(49), B => B(49), Ci => CTMP_49_port, S => 
                           S(49), Co => CTMP_50_port);
   FAI_51 : FA_1678 port map( A => A(50), B => B(50), Ci => CTMP_50_port, S => 
                           S(50), Co => CTMP_51_port);
   FAI_52 : FA_1677 port map( A => A(51), B => B(51), Ci => CTMP_51_port, S => 
                           S(51), Co => CTMP_52_port);
   FAI_53 : FA_1676 port map( A => A(52), B => B(52), Ci => CTMP_52_port, S => 
                           S(52), Co => CTMP_53_port);
   FAI_54 : FA_1675 port map( A => A(53), B => B(53), Ci => CTMP_53_port, S => 
                           S(53), Co => CTMP_54_port);
   FAI_55 : FA_1674 port map( A => A(54), B => B(54), Ci => CTMP_54_port, S => 
                           S(54), Co => CTMP_55_port);
   FAI_56 : FA_1673 port map( A => A(55), B => B(55), Ci => CTMP_55_port, S => 
                           S(55), Co => CTMP_56_port);
   FAI_57 : FA_1672 port map( A => A(56), B => B(56), Ci => CTMP_56_port, S => 
                           S(56), Co => CTMP_57_port);
   FAI_58 : FA_1671 port map( A => A(57), B => B(57), Ci => CTMP_57_port, S => 
                           S(57), Co => CTMP_58_port);
   FAI_59 : FA_1670 port map( A => A(58), B => B(58), Ci => CTMP_58_port, S => 
                           S(58), Co => CTMP_59_port);
   FAI_60 : FA_1669 port map( A => A(59), B => B(59), Ci => CTMP_59_port, S => 
                           S(59), Co => CTMP_60_port);
   FAI_61 : FA_1668 port map( A => A(60), B => B(60), Ci => CTMP_60_port, S => 
                           S(60), Co => CTMP_61_port);
   FAI_62 : FA_1667 port map( A => A(61), B => B(61), Ci => CTMP_61_port, S => 
                           S(61), Co => CTMP_62_port);
   FAI_63 : FA_1666 port map( A => A(62), B => B(62), Ci => CTMP_62_port, S => 
                           S(62), Co => CTMP_63_port);
   FAI_64 : FA_1665 port map( A => A(63), B => B(63), Ci => CTMP_63_port, S => 
                           S(63), Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity RCA_NbitRca64_26 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_NbitRca64_26;

architecture SYN_STRUCTURAL of RCA_NbitRca64_26 is

   component FA_1601
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1602
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1603
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1604
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1605
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1606
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1607
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1608
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1609
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1610
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1611
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1612
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1613
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1614
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1615
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1616
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1617
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1618
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1619
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1620
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1621
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1622
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1623
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1624
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1625
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1626
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1627
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1628
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1629
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1630
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1631
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1632
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1633
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1634
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1635
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1636
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1637
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1638
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1639
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1640
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1641
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1642
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1643
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1644
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1645
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1646
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1647
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1648
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1649
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1650
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1651
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1652
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1653
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1654
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1655
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1656
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1657
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1658
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1659
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1660
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1661
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1662
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1663
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1664
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_63_port, CTMP_62_port, CTMP_61_port, CTMP_60_port, CTMP_59_port,
      CTMP_58_port, CTMP_57_port, CTMP_56_port, CTMP_55_port, CTMP_54_port, 
      CTMP_53_port, CTMP_52_port, CTMP_51_port, CTMP_50_port, CTMP_49_port, 
      CTMP_48_port, CTMP_47_port, CTMP_46_port, CTMP_45_port, CTMP_44_port, 
      CTMP_43_port, CTMP_42_port, CTMP_41_port, CTMP_40_port, CTMP_39_port, 
      CTMP_38_port, CTMP_37_port, CTMP_36_port, CTMP_35_port, CTMP_34_port, 
      CTMP_33_port, CTMP_32_port, CTMP_31_port, CTMP_30_port, CTMP_29_port, 
      CTMP_28_port, CTMP_27_port, CTMP_26_port, CTMP_25_port, CTMP_24_port, 
      CTMP_23_port, CTMP_22_port, CTMP_21_port, CTMP_20_port, CTMP_19_port, 
      CTMP_18_port, CTMP_17_port, CTMP_16_port, CTMP_15_port, CTMP_14_port, 
      CTMP_13_port, CTMP_12_port, CTMP_11_port, CTMP_10_port, CTMP_9_port, 
      CTMP_8_port, CTMP_7_port, CTMP_6_port, CTMP_5_port, CTMP_4_port, 
      CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_1664 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_1663 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1)
                           , Co => CTMP_2_port);
   FAI_3 : FA_1662 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2)
                           , Co => CTMP_3_port);
   FAI_4 : FA_1661 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3)
                           , Co => CTMP_4_port);
   FAI_5 : FA_1660 port map( A => A(4), B => B(4), Ci => CTMP_4_port, S => S(4)
                           , Co => CTMP_5_port);
   FAI_6 : FA_1659 port map( A => A(5), B => B(5), Ci => CTMP_5_port, S => S(5)
                           , Co => CTMP_6_port);
   FAI_7 : FA_1658 port map( A => A(6), B => B(6), Ci => CTMP_6_port, S => S(6)
                           , Co => CTMP_7_port);
   FAI_8 : FA_1657 port map( A => A(7), B => B(7), Ci => CTMP_7_port, S => S(7)
                           , Co => CTMP_8_port);
   FAI_9 : FA_1656 port map( A => A(8), B => B(8), Ci => CTMP_8_port, S => S(8)
                           , Co => CTMP_9_port);
   FAI_10 : FA_1655 port map( A => A(9), B => B(9), Ci => CTMP_9_port, S => 
                           S(9), Co => CTMP_10_port);
   FAI_11 : FA_1654 port map( A => A(10), B => B(10), Ci => CTMP_10_port, S => 
                           S(10), Co => CTMP_11_port);
   FAI_12 : FA_1653 port map( A => A(11), B => B(11), Ci => CTMP_11_port, S => 
                           S(11), Co => CTMP_12_port);
   FAI_13 : FA_1652 port map( A => A(12), B => B(12), Ci => CTMP_12_port, S => 
                           S(12), Co => CTMP_13_port);
   FAI_14 : FA_1651 port map( A => A(13), B => B(13), Ci => CTMP_13_port, S => 
                           S(13), Co => CTMP_14_port);
   FAI_15 : FA_1650 port map( A => A(14), B => B(14), Ci => CTMP_14_port, S => 
                           S(14), Co => CTMP_15_port);
   FAI_16 : FA_1649 port map( A => A(15), B => B(15), Ci => CTMP_15_port, S => 
                           S(15), Co => CTMP_16_port);
   FAI_17 : FA_1648 port map( A => A(16), B => B(16), Ci => CTMP_16_port, S => 
                           S(16), Co => CTMP_17_port);
   FAI_18 : FA_1647 port map( A => A(17), B => B(17), Ci => CTMP_17_port, S => 
                           S(17), Co => CTMP_18_port);
   FAI_19 : FA_1646 port map( A => A(18), B => B(18), Ci => CTMP_18_port, S => 
                           S(18), Co => CTMP_19_port);
   FAI_20 : FA_1645 port map( A => A(19), B => B(19), Ci => CTMP_19_port, S => 
                           S(19), Co => CTMP_20_port);
   FAI_21 : FA_1644 port map( A => A(20), B => B(20), Ci => CTMP_20_port, S => 
                           S(20), Co => CTMP_21_port);
   FAI_22 : FA_1643 port map( A => A(21), B => B(21), Ci => CTMP_21_port, S => 
                           S(21), Co => CTMP_22_port);
   FAI_23 : FA_1642 port map( A => A(22), B => B(22), Ci => CTMP_22_port, S => 
                           S(22), Co => CTMP_23_port);
   FAI_24 : FA_1641 port map( A => A(23), B => B(23), Ci => CTMP_23_port, S => 
                           S(23), Co => CTMP_24_port);
   FAI_25 : FA_1640 port map( A => A(24), B => B(24), Ci => CTMP_24_port, S => 
                           S(24), Co => CTMP_25_port);
   FAI_26 : FA_1639 port map( A => A(25), B => B(25), Ci => CTMP_25_port, S => 
                           S(25), Co => CTMP_26_port);
   FAI_27 : FA_1638 port map( A => A(26), B => B(26), Ci => CTMP_26_port, S => 
                           S(26), Co => CTMP_27_port);
   FAI_28 : FA_1637 port map( A => A(27), B => B(27), Ci => CTMP_27_port, S => 
                           S(27), Co => CTMP_28_port);
   FAI_29 : FA_1636 port map( A => A(28), B => B(28), Ci => CTMP_28_port, S => 
                           S(28), Co => CTMP_29_port);
   FAI_30 : FA_1635 port map( A => A(29), B => B(29), Ci => CTMP_29_port, S => 
                           S(29), Co => CTMP_30_port);
   FAI_31 : FA_1634 port map( A => A(30), B => B(30), Ci => CTMP_30_port, S => 
                           S(30), Co => CTMP_31_port);
   FAI_32 : FA_1633 port map( A => A(31), B => B(31), Ci => CTMP_31_port, S => 
                           S(31), Co => CTMP_32_port);
   FAI_33 : FA_1632 port map( A => A(32), B => B(32), Ci => CTMP_32_port, S => 
                           S(32), Co => CTMP_33_port);
   FAI_34 : FA_1631 port map( A => A(33), B => B(33), Ci => CTMP_33_port, S => 
                           S(33), Co => CTMP_34_port);
   FAI_35 : FA_1630 port map( A => A(34), B => B(34), Ci => CTMP_34_port, S => 
                           S(34), Co => CTMP_35_port);
   FAI_36 : FA_1629 port map( A => A(35), B => B(35), Ci => CTMP_35_port, S => 
                           S(35), Co => CTMP_36_port);
   FAI_37 : FA_1628 port map( A => A(36), B => B(36), Ci => CTMP_36_port, S => 
                           S(36), Co => CTMP_37_port);
   FAI_38 : FA_1627 port map( A => A(37), B => B(37), Ci => CTMP_37_port, S => 
                           S(37), Co => CTMP_38_port);
   FAI_39 : FA_1626 port map( A => A(38), B => B(38), Ci => CTMP_38_port, S => 
                           S(38), Co => CTMP_39_port);
   FAI_40 : FA_1625 port map( A => A(39), B => B(39), Ci => CTMP_39_port, S => 
                           S(39), Co => CTMP_40_port);
   FAI_41 : FA_1624 port map( A => A(40), B => B(40), Ci => CTMP_40_port, S => 
                           S(40), Co => CTMP_41_port);
   FAI_42 : FA_1623 port map( A => A(41), B => B(41), Ci => CTMP_41_port, S => 
                           S(41), Co => CTMP_42_port);
   FAI_43 : FA_1622 port map( A => A(42), B => B(42), Ci => CTMP_42_port, S => 
                           S(42), Co => CTMP_43_port);
   FAI_44 : FA_1621 port map( A => A(43), B => B(43), Ci => CTMP_43_port, S => 
                           S(43), Co => CTMP_44_port);
   FAI_45 : FA_1620 port map( A => A(44), B => B(44), Ci => CTMP_44_port, S => 
                           S(44), Co => CTMP_45_port);
   FAI_46 : FA_1619 port map( A => A(45), B => B(45), Ci => CTMP_45_port, S => 
                           S(45), Co => CTMP_46_port);
   FAI_47 : FA_1618 port map( A => A(46), B => B(46), Ci => CTMP_46_port, S => 
                           S(46), Co => CTMP_47_port);
   FAI_48 : FA_1617 port map( A => A(47), B => B(47), Ci => CTMP_47_port, S => 
                           S(47), Co => CTMP_48_port);
   FAI_49 : FA_1616 port map( A => A(48), B => B(48), Ci => CTMP_48_port, S => 
                           S(48), Co => CTMP_49_port);
   FAI_50 : FA_1615 port map( A => A(49), B => B(49), Ci => CTMP_49_port, S => 
                           S(49), Co => CTMP_50_port);
   FAI_51 : FA_1614 port map( A => A(50), B => B(50), Ci => CTMP_50_port, S => 
                           S(50), Co => CTMP_51_port);
   FAI_52 : FA_1613 port map( A => A(51), B => B(51), Ci => CTMP_51_port, S => 
                           S(51), Co => CTMP_52_port);
   FAI_53 : FA_1612 port map( A => A(52), B => B(52), Ci => CTMP_52_port, S => 
                           S(52), Co => CTMP_53_port);
   FAI_54 : FA_1611 port map( A => A(53), B => B(53), Ci => CTMP_53_port, S => 
                           S(53), Co => CTMP_54_port);
   FAI_55 : FA_1610 port map( A => A(54), B => B(54), Ci => CTMP_54_port, S => 
                           S(54), Co => CTMP_55_port);
   FAI_56 : FA_1609 port map( A => A(55), B => B(55), Ci => CTMP_55_port, S => 
                           S(55), Co => CTMP_56_port);
   FAI_57 : FA_1608 port map( A => A(56), B => B(56), Ci => CTMP_56_port, S => 
                           S(56), Co => CTMP_57_port);
   FAI_58 : FA_1607 port map( A => A(57), B => B(57), Ci => CTMP_57_port, S => 
                           S(57), Co => CTMP_58_port);
   FAI_59 : FA_1606 port map( A => A(58), B => B(58), Ci => CTMP_58_port, S => 
                           S(58), Co => CTMP_59_port);
   FAI_60 : FA_1605 port map( A => A(59), B => B(59), Ci => CTMP_59_port, S => 
                           S(59), Co => CTMP_60_port);
   FAI_61 : FA_1604 port map( A => A(60), B => B(60), Ci => CTMP_60_port, S => 
                           S(60), Co => CTMP_61_port);
   FAI_62 : FA_1603 port map( A => A(61), B => B(61), Ci => CTMP_61_port, S => 
                           S(61), Co => CTMP_62_port);
   FAI_63 : FA_1602 port map( A => A(62), B => B(62), Ci => CTMP_62_port, S => 
                           S(62), Co => CTMP_63_port);
   FAI_64 : FA_1601 port map( A => A(63), B => B(63), Ci => CTMP_63_port, S => 
                           S(63), Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity RCA_NbitRca64_25 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_NbitRca64_25;

architecture SYN_STRUCTURAL of RCA_NbitRca64_25 is

   component FA_1537
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1538
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1539
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1540
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1541
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1542
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1543
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1544
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1545
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1546
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1547
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1548
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1549
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1550
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1551
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1552
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1553
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1554
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1555
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1556
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1557
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1558
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1559
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1560
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1561
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1562
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1563
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1564
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1565
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1566
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1567
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1568
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1569
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1570
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1571
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1572
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1573
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1574
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1575
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1576
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1577
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1578
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1579
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1580
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1581
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1582
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1583
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1584
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1585
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1586
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1587
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1588
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1589
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1590
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1591
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1592
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1593
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1594
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1595
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1596
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1597
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1598
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1599
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1600
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_63_port, CTMP_62_port, CTMP_61_port, CTMP_60_port, CTMP_59_port,
      CTMP_58_port, CTMP_57_port, CTMP_56_port, CTMP_55_port, CTMP_54_port, 
      CTMP_53_port, CTMP_52_port, CTMP_51_port, CTMP_50_port, CTMP_49_port, 
      CTMP_48_port, CTMP_47_port, CTMP_46_port, CTMP_45_port, CTMP_44_port, 
      CTMP_43_port, CTMP_42_port, CTMP_41_port, CTMP_40_port, CTMP_39_port, 
      CTMP_38_port, CTMP_37_port, CTMP_36_port, CTMP_35_port, CTMP_34_port, 
      CTMP_33_port, CTMP_32_port, CTMP_31_port, CTMP_30_port, CTMP_29_port, 
      CTMP_28_port, CTMP_27_port, CTMP_26_port, CTMP_25_port, CTMP_24_port, 
      CTMP_23_port, CTMP_22_port, CTMP_21_port, CTMP_20_port, CTMP_19_port, 
      CTMP_18_port, CTMP_17_port, CTMP_16_port, CTMP_15_port, CTMP_14_port, 
      CTMP_13_port, CTMP_12_port, CTMP_11_port, CTMP_10_port, CTMP_9_port, 
      CTMP_8_port, CTMP_7_port, CTMP_6_port, CTMP_5_port, CTMP_4_port, 
      CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_1600 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_1599 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1)
                           , Co => CTMP_2_port);
   FAI_3 : FA_1598 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2)
                           , Co => CTMP_3_port);
   FAI_4 : FA_1597 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3)
                           , Co => CTMP_4_port);
   FAI_5 : FA_1596 port map( A => A(4), B => B(4), Ci => CTMP_4_port, S => S(4)
                           , Co => CTMP_5_port);
   FAI_6 : FA_1595 port map( A => A(5), B => B(5), Ci => CTMP_5_port, S => S(5)
                           , Co => CTMP_6_port);
   FAI_7 : FA_1594 port map( A => A(6), B => B(6), Ci => CTMP_6_port, S => S(6)
                           , Co => CTMP_7_port);
   FAI_8 : FA_1593 port map( A => A(7), B => B(7), Ci => CTMP_7_port, S => S(7)
                           , Co => CTMP_8_port);
   FAI_9 : FA_1592 port map( A => A(8), B => B(8), Ci => CTMP_8_port, S => S(8)
                           , Co => CTMP_9_port);
   FAI_10 : FA_1591 port map( A => A(9), B => B(9), Ci => CTMP_9_port, S => 
                           S(9), Co => CTMP_10_port);
   FAI_11 : FA_1590 port map( A => A(10), B => B(10), Ci => CTMP_10_port, S => 
                           S(10), Co => CTMP_11_port);
   FAI_12 : FA_1589 port map( A => A(11), B => B(11), Ci => CTMP_11_port, S => 
                           S(11), Co => CTMP_12_port);
   FAI_13 : FA_1588 port map( A => A(12), B => B(12), Ci => CTMP_12_port, S => 
                           S(12), Co => CTMP_13_port);
   FAI_14 : FA_1587 port map( A => A(13), B => B(13), Ci => CTMP_13_port, S => 
                           S(13), Co => CTMP_14_port);
   FAI_15 : FA_1586 port map( A => A(14), B => B(14), Ci => CTMP_14_port, S => 
                           S(14), Co => CTMP_15_port);
   FAI_16 : FA_1585 port map( A => A(15), B => B(15), Ci => CTMP_15_port, S => 
                           S(15), Co => CTMP_16_port);
   FAI_17 : FA_1584 port map( A => A(16), B => B(16), Ci => CTMP_16_port, S => 
                           S(16), Co => CTMP_17_port);
   FAI_18 : FA_1583 port map( A => A(17), B => B(17), Ci => CTMP_17_port, S => 
                           S(17), Co => CTMP_18_port);
   FAI_19 : FA_1582 port map( A => A(18), B => B(18), Ci => CTMP_18_port, S => 
                           S(18), Co => CTMP_19_port);
   FAI_20 : FA_1581 port map( A => A(19), B => B(19), Ci => CTMP_19_port, S => 
                           S(19), Co => CTMP_20_port);
   FAI_21 : FA_1580 port map( A => A(20), B => B(20), Ci => CTMP_20_port, S => 
                           S(20), Co => CTMP_21_port);
   FAI_22 : FA_1579 port map( A => A(21), B => B(21), Ci => CTMP_21_port, S => 
                           S(21), Co => CTMP_22_port);
   FAI_23 : FA_1578 port map( A => A(22), B => B(22), Ci => CTMP_22_port, S => 
                           S(22), Co => CTMP_23_port);
   FAI_24 : FA_1577 port map( A => A(23), B => B(23), Ci => CTMP_23_port, S => 
                           S(23), Co => CTMP_24_port);
   FAI_25 : FA_1576 port map( A => A(24), B => B(24), Ci => CTMP_24_port, S => 
                           S(24), Co => CTMP_25_port);
   FAI_26 : FA_1575 port map( A => A(25), B => B(25), Ci => CTMP_25_port, S => 
                           S(25), Co => CTMP_26_port);
   FAI_27 : FA_1574 port map( A => A(26), B => B(26), Ci => CTMP_26_port, S => 
                           S(26), Co => CTMP_27_port);
   FAI_28 : FA_1573 port map( A => A(27), B => B(27), Ci => CTMP_27_port, S => 
                           S(27), Co => CTMP_28_port);
   FAI_29 : FA_1572 port map( A => A(28), B => B(28), Ci => CTMP_28_port, S => 
                           S(28), Co => CTMP_29_port);
   FAI_30 : FA_1571 port map( A => A(29), B => B(29), Ci => CTMP_29_port, S => 
                           S(29), Co => CTMP_30_port);
   FAI_31 : FA_1570 port map( A => A(30), B => B(30), Ci => CTMP_30_port, S => 
                           S(30), Co => CTMP_31_port);
   FAI_32 : FA_1569 port map( A => A(31), B => B(31), Ci => CTMP_31_port, S => 
                           S(31), Co => CTMP_32_port);
   FAI_33 : FA_1568 port map( A => A(32), B => B(32), Ci => CTMP_32_port, S => 
                           S(32), Co => CTMP_33_port);
   FAI_34 : FA_1567 port map( A => A(33), B => B(33), Ci => CTMP_33_port, S => 
                           S(33), Co => CTMP_34_port);
   FAI_35 : FA_1566 port map( A => A(34), B => B(34), Ci => CTMP_34_port, S => 
                           S(34), Co => CTMP_35_port);
   FAI_36 : FA_1565 port map( A => A(35), B => B(35), Ci => CTMP_35_port, S => 
                           S(35), Co => CTMP_36_port);
   FAI_37 : FA_1564 port map( A => A(36), B => B(36), Ci => CTMP_36_port, S => 
                           S(36), Co => CTMP_37_port);
   FAI_38 : FA_1563 port map( A => A(37), B => B(37), Ci => CTMP_37_port, S => 
                           S(37), Co => CTMP_38_port);
   FAI_39 : FA_1562 port map( A => A(38), B => B(38), Ci => CTMP_38_port, S => 
                           S(38), Co => CTMP_39_port);
   FAI_40 : FA_1561 port map( A => A(39), B => B(39), Ci => CTMP_39_port, S => 
                           S(39), Co => CTMP_40_port);
   FAI_41 : FA_1560 port map( A => A(40), B => B(40), Ci => CTMP_40_port, S => 
                           S(40), Co => CTMP_41_port);
   FAI_42 : FA_1559 port map( A => A(41), B => B(41), Ci => CTMP_41_port, S => 
                           S(41), Co => CTMP_42_port);
   FAI_43 : FA_1558 port map( A => A(42), B => B(42), Ci => CTMP_42_port, S => 
                           S(42), Co => CTMP_43_port);
   FAI_44 : FA_1557 port map( A => A(43), B => B(43), Ci => CTMP_43_port, S => 
                           S(43), Co => CTMP_44_port);
   FAI_45 : FA_1556 port map( A => A(44), B => B(44), Ci => CTMP_44_port, S => 
                           S(44), Co => CTMP_45_port);
   FAI_46 : FA_1555 port map( A => A(45), B => B(45), Ci => CTMP_45_port, S => 
                           S(45), Co => CTMP_46_port);
   FAI_47 : FA_1554 port map( A => A(46), B => B(46), Ci => CTMP_46_port, S => 
                           S(46), Co => CTMP_47_port);
   FAI_48 : FA_1553 port map( A => A(47), B => B(47), Ci => CTMP_47_port, S => 
                           S(47), Co => CTMP_48_port);
   FAI_49 : FA_1552 port map( A => A(48), B => B(48), Ci => CTMP_48_port, S => 
                           S(48), Co => CTMP_49_port);
   FAI_50 : FA_1551 port map( A => A(49), B => B(49), Ci => CTMP_49_port, S => 
                           S(49), Co => CTMP_50_port);
   FAI_51 : FA_1550 port map( A => A(50), B => B(50), Ci => CTMP_50_port, S => 
                           S(50), Co => CTMP_51_port);
   FAI_52 : FA_1549 port map( A => A(51), B => B(51), Ci => CTMP_51_port, S => 
                           S(51), Co => CTMP_52_port);
   FAI_53 : FA_1548 port map( A => A(52), B => B(52), Ci => CTMP_52_port, S => 
                           S(52), Co => CTMP_53_port);
   FAI_54 : FA_1547 port map( A => A(53), B => B(53), Ci => CTMP_53_port, S => 
                           S(53), Co => CTMP_54_port);
   FAI_55 : FA_1546 port map( A => A(54), B => B(54), Ci => CTMP_54_port, S => 
                           S(54), Co => CTMP_55_port);
   FAI_56 : FA_1545 port map( A => A(55), B => B(55), Ci => CTMP_55_port, S => 
                           S(55), Co => CTMP_56_port);
   FAI_57 : FA_1544 port map( A => A(56), B => B(56), Ci => CTMP_56_port, S => 
                           S(56), Co => CTMP_57_port);
   FAI_58 : FA_1543 port map( A => A(57), B => B(57), Ci => CTMP_57_port, S => 
                           S(57), Co => CTMP_58_port);
   FAI_59 : FA_1542 port map( A => A(58), B => B(58), Ci => CTMP_58_port, S => 
                           S(58), Co => CTMP_59_port);
   FAI_60 : FA_1541 port map( A => A(59), B => B(59), Ci => CTMP_59_port, S => 
                           S(59), Co => CTMP_60_port);
   FAI_61 : FA_1540 port map( A => A(60), B => B(60), Ci => CTMP_60_port, S => 
                           S(60), Co => CTMP_61_port);
   FAI_62 : FA_1539 port map( A => A(61), B => B(61), Ci => CTMP_61_port, S => 
                           S(61), Co => CTMP_62_port);
   FAI_63 : FA_1538 port map( A => A(62), B => B(62), Ci => CTMP_62_port, S => 
                           S(62), Co => CTMP_63_port);
   FAI_64 : FA_1537 port map( A => A(63), B => B(63), Ci => CTMP_63_port, S => 
                           S(63), Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity RCA_NbitRca64_24 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_NbitRca64_24;

architecture SYN_STRUCTURAL of RCA_NbitRca64_24 is

   component FA_1473
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1474
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1475
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1476
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1477
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1478
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1479
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1480
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1481
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1482
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1483
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1484
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1485
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1486
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1487
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1488
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1489
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1490
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1491
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1492
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1493
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1494
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1495
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1496
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1497
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1498
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1499
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1500
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1501
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1502
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1503
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1504
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1505
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1506
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1507
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1508
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1509
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1510
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1511
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1512
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1513
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1514
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1515
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1516
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1517
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1518
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1519
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1520
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1521
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1522
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1523
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1524
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1525
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1526
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1527
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1528
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1529
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1530
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1531
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1532
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1533
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1534
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1535
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1536
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_63_port, CTMP_62_port, CTMP_61_port, CTMP_60_port, CTMP_59_port,
      CTMP_58_port, CTMP_57_port, CTMP_56_port, CTMP_55_port, CTMP_54_port, 
      CTMP_53_port, CTMP_52_port, CTMP_51_port, CTMP_50_port, CTMP_49_port, 
      CTMP_48_port, CTMP_47_port, CTMP_46_port, CTMP_45_port, CTMP_44_port, 
      CTMP_43_port, CTMP_42_port, CTMP_41_port, CTMP_40_port, CTMP_39_port, 
      CTMP_38_port, CTMP_37_port, CTMP_36_port, CTMP_35_port, CTMP_34_port, 
      CTMP_33_port, CTMP_32_port, CTMP_31_port, CTMP_30_port, CTMP_29_port, 
      CTMP_28_port, CTMP_27_port, CTMP_26_port, CTMP_25_port, CTMP_24_port, 
      CTMP_23_port, CTMP_22_port, CTMP_21_port, CTMP_20_port, CTMP_19_port, 
      CTMP_18_port, CTMP_17_port, CTMP_16_port, CTMP_15_port, CTMP_14_port, 
      CTMP_13_port, CTMP_12_port, CTMP_11_port, CTMP_10_port, CTMP_9_port, 
      CTMP_8_port, CTMP_7_port, CTMP_6_port, CTMP_5_port, CTMP_4_port, 
      CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_1536 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_1535 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1)
                           , Co => CTMP_2_port);
   FAI_3 : FA_1534 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2)
                           , Co => CTMP_3_port);
   FAI_4 : FA_1533 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3)
                           , Co => CTMP_4_port);
   FAI_5 : FA_1532 port map( A => A(4), B => B(4), Ci => CTMP_4_port, S => S(4)
                           , Co => CTMP_5_port);
   FAI_6 : FA_1531 port map( A => A(5), B => B(5), Ci => CTMP_5_port, S => S(5)
                           , Co => CTMP_6_port);
   FAI_7 : FA_1530 port map( A => A(6), B => B(6), Ci => CTMP_6_port, S => S(6)
                           , Co => CTMP_7_port);
   FAI_8 : FA_1529 port map( A => A(7), B => B(7), Ci => CTMP_7_port, S => S(7)
                           , Co => CTMP_8_port);
   FAI_9 : FA_1528 port map( A => A(8), B => B(8), Ci => CTMP_8_port, S => S(8)
                           , Co => CTMP_9_port);
   FAI_10 : FA_1527 port map( A => A(9), B => B(9), Ci => CTMP_9_port, S => 
                           S(9), Co => CTMP_10_port);
   FAI_11 : FA_1526 port map( A => A(10), B => B(10), Ci => CTMP_10_port, S => 
                           S(10), Co => CTMP_11_port);
   FAI_12 : FA_1525 port map( A => A(11), B => B(11), Ci => CTMP_11_port, S => 
                           S(11), Co => CTMP_12_port);
   FAI_13 : FA_1524 port map( A => A(12), B => B(12), Ci => CTMP_12_port, S => 
                           S(12), Co => CTMP_13_port);
   FAI_14 : FA_1523 port map( A => A(13), B => B(13), Ci => CTMP_13_port, S => 
                           S(13), Co => CTMP_14_port);
   FAI_15 : FA_1522 port map( A => A(14), B => B(14), Ci => CTMP_14_port, S => 
                           S(14), Co => CTMP_15_port);
   FAI_16 : FA_1521 port map( A => A(15), B => B(15), Ci => CTMP_15_port, S => 
                           S(15), Co => CTMP_16_port);
   FAI_17 : FA_1520 port map( A => A(16), B => B(16), Ci => CTMP_16_port, S => 
                           S(16), Co => CTMP_17_port);
   FAI_18 : FA_1519 port map( A => A(17), B => B(17), Ci => CTMP_17_port, S => 
                           S(17), Co => CTMP_18_port);
   FAI_19 : FA_1518 port map( A => A(18), B => B(18), Ci => CTMP_18_port, S => 
                           S(18), Co => CTMP_19_port);
   FAI_20 : FA_1517 port map( A => A(19), B => B(19), Ci => CTMP_19_port, S => 
                           S(19), Co => CTMP_20_port);
   FAI_21 : FA_1516 port map( A => A(20), B => B(20), Ci => CTMP_20_port, S => 
                           S(20), Co => CTMP_21_port);
   FAI_22 : FA_1515 port map( A => A(21), B => B(21), Ci => CTMP_21_port, S => 
                           S(21), Co => CTMP_22_port);
   FAI_23 : FA_1514 port map( A => A(22), B => B(22), Ci => CTMP_22_port, S => 
                           S(22), Co => CTMP_23_port);
   FAI_24 : FA_1513 port map( A => A(23), B => B(23), Ci => CTMP_23_port, S => 
                           S(23), Co => CTMP_24_port);
   FAI_25 : FA_1512 port map( A => A(24), B => B(24), Ci => CTMP_24_port, S => 
                           S(24), Co => CTMP_25_port);
   FAI_26 : FA_1511 port map( A => A(25), B => B(25), Ci => CTMP_25_port, S => 
                           S(25), Co => CTMP_26_port);
   FAI_27 : FA_1510 port map( A => A(26), B => B(26), Ci => CTMP_26_port, S => 
                           S(26), Co => CTMP_27_port);
   FAI_28 : FA_1509 port map( A => A(27), B => B(27), Ci => CTMP_27_port, S => 
                           S(27), Co => CTMP_28_port);
   FAI_29 : FA_1508 port map( A => A(28), B => B(28), Ci => CTMP_28_port, S => 
                           S(28), Co => CTMP_29_port);
   FAI_30 : FA_1507 port map( A => A(29), B => B(29), Ci => CTMP_29_port, S => 
                           S(29), Co => CTMP_30_port);
   FAI_31 : FA_1506 port map( A => A(30), B => B(30), Ci => CTMP_30_port, S => 
                           S(30), Co => CTMP_31_port);
   FAI_32 : FA_1505 port map( A => A(31), B => B(31), Ci => CTMP_31_port, S => 
                           S(31), Co => CTMP_32_port);
   FAI_33 : FA_1504 port map( A => A(32), B => B(32), Ci => CTMP_32_port, S => 
                           S(32), Co => CTMP_33_port);
   FAI_34 : FA_1503 port map( A => A(33), B => B(33), Ci => CTMP_33_port, S => 
                           S(33), Co => CTMP_34_port);
   FAI_35 : FA_1502 port map( A => A(34), B => B(34), Ci => CTMP_34_port, S => 
                           S(34), Co => CTMP_35_port);
   FAI_36 : FA_1501 port map( A => A(35), B => B(35), Ci => CTMP_35_port, S => 
                           S(35), Co => CTMP_36_port);
   FAI_37 : FA_1500 port map( A => A(36), B => B(36), Ci => CTMP_36_port, S => 
                           S(36), Co => CTMP_37_port);
   FAI_38 : FA_1499 port map( A => A(37), B => B(37), Ci => CTMP_37_port, S => 
                           S(37), Co => CTMP_38_port);
   FAI_39 : FA_1498 port map( A => A(38), B => B(38), Ci => CTMP_38_port, S => 
                           S(38), Co => CTMP_39_port);
   FAI_40 : FA_1497 port map( A => A(39), B => B(39), Ci => CTMP_39_port, S => 
                           S(39), Co => CTMP_40_port);
   FAI_41 : FA_1496 port map( A => A(40), B => B(40), Ci => CTMP_40_port, S => 
                           S(40), Co => CTMP_41_port);
   FAI_42 : FA_1495 port map( A => A(41), B => B(41), Ci => CTMP_41_port, S => 
                           S(41), Co => CTMP_42_port);
   FAI_43 : FA_1494 port map( A => A(42), B => B(42), Ci => CTMP_42_port, S => 
                           S(42), Co => CTMP_43_port);
   FAI_44 : FA_1493 port map( A => A(43), B => B(43), Ci => CTMP_43_port, S => 
                           S(43), Co => CTMP_44_port);
   FAI_45 : FA_1492 port map( A => A(44), B => B(44), Ci => CTMP_44_port, S => 
                           S(44), Co => CTMP_45_port);
   FAI_46 : FA_1491 port map( A => A(45), B => B(45), Ci => CTMP_45_port, S => 
                           S(45), Co => CTMP_46_port);
   FAI_47 : FA_1490 port map( A => A(46), B => B(46), Ci => CTMP_46_port, S => 
                           S(46), Co => CTMP_47_port);
   FAI_48 : FA_1489 port map( A => A(47), B => B(47), Ci => CTMP_47_port, S => 
                           S(47), Co => CTMP_48_port);
   FAI_49 : FA_1488 port map( A => A(48), B => B(48), Ci => CTMP_48_port, S => 
                           S(48), Co => CTMP_49_port);
   FAI_50 : FA_1487 port map( A => A(49), B => B(49), Ci => CTMP_49_port, S => 
                           S(49), Co => CTMP_50_port);
   FAI_51 : FA_1486 port map( A => A(50), B => B(50), Ci => CTMP_50_port, S => 
                           S(50), Co => CTMP_51_port);
   FAI_52 : FA_1485 port map( A => A(51), B => B(51), Ci => CTMP_51_port, S => 
                           S(51), Co => CTMP_52_port);
   FAI_53 : FA_1484 port map( A => A(52), B => B(52), Ci => CTMP_52_port, S => 
                           S(52), Co => CTMP_53_port);
   FAI_54 : FA_1483 port map( A => A(53), B => B(53), Ci => CTMP_53_port, S => 
                           S(53), Co => CTMP_54_port);
   FAI_55 : FA_1482 port map( A => A(54), B => B(54), Ci => CTMP_54_port, S => 
                           S(54), Co => CTMP_55_port);
   FAI_56 : FA_1481 port map( A => A(55), B => B(55), Ci => CTMP_55_port, S => 
                           S(55), Co => CTMP_56_port);
   FAI_57 : FA_1480 port map( A => A(56), B => B(56), Ci => CTMP_56_port, S => 
                           S(56), Co => CTMP_57_port);
   FAI_58 : FA_1479 port map( A => A(57), B => B(57), Ci => CTMP_57_port, S => 
                           S(57), Co => CTMP_58_port);
   FAI_59 : FA_1478 port map( A => A(58), B => B(58), Ci => CTMP_58_port, S => 
                           S(58), Co => CTMP_59_port);
   FAI_60 : FA_1477 port map( A => A(59), B => B(59), Ci => CTMP_59_port, S => 
                           S(59), Co => CTMP_60_port);
   FAI_61 : FA_1476 port map( A => A(60), B => B(60), Ci => CTMP_60_port, S => 
                           S(60), Co => CTMP_61_port);
   FAI_62 : FA_1475 port map( A => A(61), B => B(61), Ci => CTMP_61_port, S => 
                           S(61), Co => CTMP_62_port);
   FAI_63 : FA_1474 port map( A => A(62), B => B(62), Ci => CTMP_62_port, S => 
                           S(62), Co => CTMP_63_port);
   FAI_64 : FA_1473 port map( A => A(63), B => B(63), Ci => CTMP_63_port, S => 
                           S(63), Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity RCA_NbitRca64_23 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_NbitRca64_23;

architecture SYN_STRUCTURAL of RCA_NbitRca64_23 is

   component FA_1409
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1410
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1411
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1412
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1413
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1414
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1415
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1416
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1417
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1418
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1419
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1420
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1421
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1422
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1423
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1424
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1425
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1426
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1427
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1428
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1429
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1430
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1431
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1432
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1433
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1434
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1435
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1436
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1437
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1438
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1439
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1440
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1441
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1442
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1443
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1444
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1445
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1446
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1447
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1448
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1449
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1450
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1451
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1452
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1453
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1454
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1455
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1456
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1457
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1458
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1459
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1460
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1461
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1462
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1463
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1464
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1465
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1466
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1467
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1468
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1469
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1470
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1471
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1472
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_63_port, CTMP_62_port, CTMP_61_port, CTMP_60_port, CTMP_59_port,
      CTMP_58_port, CTMP_57_port, CTMP_56_port, CTMP_55_port, CTMP_54_port, 
      CTMP_53_port, CTMP_52_port, CTMP_51_port, CTMP_50_port, CTMP_49_port, 
      CTMP_48_port, CTMP_47_port, CTMP_46_port, CTMP_45_port, CTMP_44_port, 
      CTMP_43_port, CTMP_42_port, CTMP_41_port, CTMP_40_port, CTMP_39_port, 
      CTMP_38_port, CTMP_37_port, CTMP_36_port, CTMP_35_port, CTMP_34_port, 
      CTMP_33_port, CTMP_32_port, CTMP_31_port, CTMP_30_port, CTMP_29_port, 
      CTMP_28_port, CTMP_27_port, CTMP_26_port, CTMP_25_port, CTMP_24_port, 
      CTMP_23_port, CTMP_22_port, CTMP_21_port, CTMP_20_port, CTMP_19_port, 
      CTMP_18_port, CTMP_17_port, CTMP_16_port, CTMP_15_port, CTMP_14_port, 
      CTMP_13_port, CTMP_12_port, CTMP_11_port, CTMP_10_port, CTMP_9_port, 
      CTMP_8_port, CTMP_7_port, CTMP_6_port, CTMP_5_port, CTMP_4_port, 
      CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_1472 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_1471 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1)
                           , Co => CTMP_2_port);
   FAI_3 : FA_1470 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2)
                           , Co => CTMP_3_port);
   FAI_4 : FA_1469 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3)
                           , Co => CTMP_4_port);
   FAI_5 : FA_1468 port map( A => A(4), B => B(4), Ci => CTMP_4_port, S => S(4)
                           , Co => CTMP_5_port);
   FAI_6 : FA_1467 port map( A => A(5), B => B(5), Ci => CTMP_5_port, S => S(5)
                           , Co => CTMP_6_port);
   FAI_7 : FA_1466 port map( A => A(6), B => B(6), Ci => CTMP_6_port, S => S(6)
                           , Co => CTMP_7_port);
   FAI_8 : FA_1465 port map( A => A(7), B => B(7), Ci => CTMP_7_port, S => S(7)
                           , Co => CTMP_8_port);
   FAI_9 : FA_1464 port map( A => A(8), B => B(8), Ci => CTMP_8_port, S => S(8)
                           , Co => CTMP_9_port);
   FAI_10 : FA_1463 port map( A => A(9), B => B(9), Ci => CTMP_9_port, S => 
                           S(9), Co => CTMP_10_port);
   FAI_11 : FA_1462 port map( A => A(10), B => B(10), Ci => CTMP_10_port, S => 
                           S(10), Co => CTMP_11_port);
   FAI_12 : FA_1461 port map( A => A(11), B => B(11), Ci => CTMP_11_port, S => 
                           S(11), Co => CTMP_12_port);
   FAI_13 : FA_1460 port map( A => A(12), B => B(12), Ci => CTMP_12_port, S => 
                           S(12), Co => CTMP_13_port);
   FAI_14 : FA_1459 port map( A => A(13), B => B(13), Ci => CTMP_13_port, S => 
                           S(13), Co => CTMP_14_port);
   FAI_15 : FA_1458 port map( A => A(14), B => B(14), Ci => CTMP_14_port, S => 
                           S(14), Co => CTMP_15_port);
   FAI_16 : FA_1457 port map( A => A(15), B => B(15), Ci => CTMP_15_port, S => 
                           S(15), Co => CTMP_16_port);
   FAI_17 : FA_1456 port map( A => A(16), B => B(16), Ci => CTMP_16_port, S => 
                           S(16), Co => CTMP_17_port);
   FAI_18 : FA_1455 port map( A => A(17), B => B(17), Ci => CTMP_17_port, S => 
                           S(17), Co => CTMP_18_port);
   FAI_19 : FA_1454 port map( A => A(18), B => B(18), Ci => CTMP_18_port, S => 
                           S(18), Co => CTMP_19_port);
   FAI_20 : FA_1453 port map( A => A(19), B => B(19), Ci => CTMP_19_port, S => 
                           S(19), Co => CTMP_20_port);
   FAI_21 : FA_1452 port map( A => A(20), B => B(20), Ci => CTMP_20_port, S => 
                           S(20), Co => CTMP_21_port);
   FAI_22 : FA_1451 port map( A => A(21), B => B(21), Ci => CTMP_21_port, S => 
                           S(21), Co => CTMP_22_port);
   FAI_23 : FA_1450 port map( A => A(22), B => B(22), Ci => CTMP_22_port, S => 
                           S(22), Co => CTMP_23_port);
   FAI_24 : FA_1449 port map( A => A(23), B => B(23), Ci => CTMP_23_port, S => 
                           S(23), Co => CTMP_24_port);
   FAI_25 : FA_1448 port map( A => A(24), B => B(24), Ci => CTMP_24_port, S => 
                           S(24), Co => CTMP_25_port);
   FAI_26 : FA_1447 port map( A => A(25), B => B(25), Ci => CTMP_25_port, S => 
                           S(25), Co => CTMP_26_port);
   FAI_27 : FA_1446 port map( A => A(26), B => B(26), Ci => CTMP_26_port, S => 
                           S(26), Co => CTMP_27_port);
   FAI_28 : FA_1445 port map( A => A(27), B => B(27), Ci => CTMP_27_port, S => 
                           S(27), Co => CTMP_28_port);
   FAI_29 : FA_1444 port map( A => A(28), B => B(28), Ci => CTMP_28_port, S => 
                           S(28), Co => CTMP_29_port);
   FAI_30 : FA_1443 port map( A => A(29), B => B(29), Ci => CTMP_29_port, S => 
                           S(29), Co => CTMP_30_port);
   FAI_31 : FA_1442 port map( A => A(30), B => B(30), Ci => CTMP_30_port, S => 
                           S(30), Co => CTMP_31_port);
   FAI_32 : FA_1441 port map( A => A(31), B => B(31), Ci => CTMP_31_port, S => 
                           S(31), Co => CTMP_32_port);
   FAI_33 : FA_1440 port map( A => A(32), B => B(32), Ci => CTMP_32_port, S => 
                           S(32), Co => CTMP_33_port);
   FAI_34 : FA_1439 port map( A => A(33), B => B(33), Ci => CTMP_33_port, S => 
                           S(33), Co => CTMP_34_port);
   FAI_35 : FA_1438 port map( A => A(34), B => B(34), Ci => CTMP_34_port, S => 
                           S(34), Co => CTMP_35_port);
   FAI_36 : FA_1437 port map( A => A(35), B => B(35), Ci => CTMP_35_port, S => 
                           S(35), Co => CTMP_36_port);
   FAI_37 : FA_1436 port map( A => A(36), B => B(36), Ci => CTMP_36_port, S => 
                           S(36), Co => CTMP_37_port);
   FAI_38 : FA_1435 port map( A => A(37), B => B(37), Ci => CTMP_37_port, S => 
                           S(37), Co => CTMP_38_port);
   FAI_39 : FA_1434 port map( A => A(38), B => B(38), Ci => CTMP_38_port, S => 
                           S(38), Co => CTMP_39_port);
   FAI_40 : FA_1433 port map( A => A(39), B => B(39), Ci => CTMP_39_port, S => 
                           S(39), Co => CTMP_40_port);
   FAI_41 : FA_1432 port map( A => A(40), B => B(40), Ci => CTMP_40_port, S => 
                           S(40), Co => CTMP_41_port);
   FAI_42 : FA_1431 port map( A => A(41), B => B(41), Ci => CTMP_41_port, S => 
                           S(41), Co => CTMP_42_port);
   FAI_43 : FA_1430 port map( A => A(42), B => B(42), Ci => CTMP_42_port, S => 
                           S(42), Co => CTMP_43_port);
   FAI_44 : FA_1429 port map( A => A(43), B => B(43), Ci => CTMP_43_port, S => 
                           S(43), Co => CTMP_44_port);
   FAI_45 : FA_1428 port map( A => A(44), B => B(44), Ci => CTMP_44_port, S => 
                           S(44), Co => CTMP_45_port);
   FAI_46 : FA_1427 port map( A => A(45), B => B(45), Ci => CTMP_45_port, S => 
                           S(45), Co => CTMP_46_port);
   FAI_47 : FA_1426 port map( A => A(46), B => B(46), Ci => CTMP_46_port, S => 
                           S(46), Co => CTMP_47_port);
   FAI_48 : FA_1425 port map( A => A(47), B => B(47), Ci => CTMP_47_port, S => 
                           S(47), Co => CTMP_48_port);
   FAI_49 : FA_1424 port map( A => A(48), B => B(48), Ci => CTMP_48_port, S => 
                           S(48), Co => CTMP_49_port);
   FAI_50 : FA_1423 port map( A => A(49), B => B(49), Ci => CTMP_49_port, S => 
                           S(49), Co => CTMP_50_port);
   FAI_51 : FA_1422 port map( A => A(50), B => B(50), Ci => CTMP_50_port, S => 
                           S(50), Co => CTMP_51_port);
   FAI_52 : FA_1421 port map( A => A(51), B => B(51), Ci => CTMP_51_port, S => 
                           S(51), Co => CTMP_52_port);
   FAI_53 : FA_1420 port map( A => A(52), B => B(52), Ci => CTMP_52_port, S => 
                           S(52), Co => CTMP_53_port);
   FAI_54 : FA_1419 port map( A => A(53), B => B(53), Ci => CTMP_53_port, S => 
                           S(53), Co => CTMP_54_port);
   FAI_55 : FA_1418 port map( A => A(54), B => B(54), Ci => CTMP_54_port, S => 
                           S(54), Co => CTMP_55_port);
   FAI_56 : FA_1417 port map( A => A(55), B => B(55), Ci => CTMP_55_port, S => 
                           S(55), Co => CTMP_56_port);
   FAI_57 : FA_1416 port map( A => A(56), B => B(56), Ci => CTMP_56_port, S => 
                           S(56), Co => CTMP_57_port);
   FAI_58 : FA_1415 port map( A => A(57), B => B(57), Ci => CTMP_57_port, S => 
                           S(57), Co => CTMP_58_port);
   FAI_59 : FA_1414 port map( A => A(58), B => B(58), Ci => CTMP_58_port, S => 
                           S(58), Co => CTMP_59_port);
   FAI_60 : FA_1413 port map( A => A(59), B => B(59), Ci => CTMP_59_port, S => 
                           S(59), Co => CTMP_60_port);
   FAI_61 : FA_1412 port map( A => A(60), B => B(60), Ci => CTMP_60_port, S => 
                           S(60), Co => CTMP_61_port);
   FAI_62 : FA_1411 port map( A => A(61), B => B(61), Ci => CTMP_61_port, S => 
                           S(61), Co => CTMP_62_port);
   FAI_63 : FA_1410 port map( A => A(62), B => B(62), Ci => CTMP_62_port, S => 
                           S(62), Co => CTMP_63_port);
   FAI_64 : FA_1409 port map( A => A(63), B => B(63), Ci => CTMP_63_port, S => 
                           S(63), Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity RCA_NbitRca64_22 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_NbitRca64_22;

architecture SYN_STRUCTURAL of RCA_NbitRca64_22 is

   component FA_1345
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1346
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1347
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1348
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1349
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1350
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1351
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1352
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1353
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1354
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1355
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1356
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1357
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1358
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1359
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1360
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1361
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1362
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1363
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1364
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1365
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1366
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1367
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1368
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1369
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1370
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1371
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1372
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1373
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1374
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1375
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1376
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1377
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1378
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1379
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1380
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1381
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1382
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1383
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1384
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1385
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1386
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1387
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1388
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1389
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1390
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1391
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1392
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1393
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1394
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1395
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1396
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1397
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1398
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1399
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1400
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1401
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1402
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1403
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1404
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1405
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1406
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1407
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1408
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_63_port, CTMP_62_port, CTMP_61_port, CTMP_60_port, CTMP_59_port,
      CTMP_58_port, CTMP_57_port, CTMP_56_port, CTMP_55_port, CTMP_54_port, 
      CTMP_53_port, CTMP_52_port, CTMP_51_port, CTMP_50_port, CTMP_49_port, 
      CTMP_48_port, CTMP_47_port, CTMP_46_port, CTMP_45_port, CTMP_44_port, 
      CTMP_43_port, CTMP_42_port, CTMP_41_port, CTMP_40_port, CTMP_39_port, 
      CTMP_38_port, CTMP_37_port, CTMP_36_port, CTMP_35_port, CTMP_34_port, 
      CTMP_33_port, CTMP_32_port, CTMP_31_port, CTMP_30_port, CTMP_29_port, 
      CTMP_28_port, CTMP_27_port, CTMP_26_port, CTMP_25_port, CTMP_24_port, 
      CTMP_23_port, CTMP_22_port, CTMP_21_port, CTMP_20_port, CTMP_19_port, 
      CTMP_18_port, CTMP_17_port, CTMP_16_port, CTMP_15_port, CTMP_14_port, 
      CTMP_13_port, CTMP_12_port, CTMP_11_port, CTMP_10_port, CTMP_9_port, 
      CTMP_8_port, CTMP_7_port, CTMP_6_port, CTMP_5_port, CTMP_4_port, 
      CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_1408 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_1407 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1)
                           , Co => CTMP_2_port);
   FAI_3 : FA_1406 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2)
                           , Co => CTMP_3_port);
   FAI_4 : FA_1405 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3)
                           , Co => CTMP_4_port);
   FAI_5 : FA_1404 port map( A => A(4), B => B(4), Ci => CTMP_4_port, S => S(4)
                           , Co => CTMP_5_port);
   FAI_6 : FA_1403 port map( A => A(5), B => B(5), Ci => CTMP_5_port, S => S(5)
                           , Co => CTMP_6_port);
   FAI_7 : FA_1402 port map( A => A(6), B => B(6), Ci => CTMP_6_port, S => S(6)
                           , Co => CTMP_7_port);
   FAI_8 : FA_1401 port map( A => A(7), B => B(7), Ci => CTMP_7_port, S => S(7)
                           , Co => CTMP_8_port);
   FAI_9 : FA_1400 port map( A => A(8), B => B(8), Ci => CTMP_8_port, S => S(8)
                           , Co => CTMP_9_port);
   FAI_10 : FA_1399 port map( A => A(9), B => B(9), Ci => CTMP_9_port, S => 
                           S(9), Co => CTMP_10_port);
   FAI_11 : FA_1398 port map( A => A(10), B => B(10), Ci => CTMP_10_port, S => 
                           S(10), Co => CTMP_11_port);
   FAI_12 : FA_1397 port map( A => A(11), B => B(11), Ci => CTMP_11_port, S => 
                           S(11), Co => CTMP_12_port);
   FAI_13 : FA_1396 port map( A => A(12), B => B(12), Ci => CTMP_12_port, S => 
                           S(12), Co => CTMP_13_port);
   FAI_14 : FA_1395 port map( A => A(13), B => B(13), Ci => CTMP_13_port, S => 
                           S(13), Co => CTMP_14_port);
   FAI_15 : FA_1394 port map( A => A(14), B => B(14), Ci => CTMP_14_port, S => 
                           S(14), Co => CTMP_15_port);
   FAI_16 : FA_1393 port map( A => A(15), B => B(15), Ci => CTMP_15_port, S => 
                           S(15), Co => CTMP_16_port);
   FAI_17 : FA_1392 port map( A => A(16), B => B(16), Ci => CTMP_16_port, S => 
                           S(16), Co => CTMP_17_port);
   FAI_18 : FA_1391 port map( A => A(17), B => B(17), Ci => CTMP_17_port, S => 
                           S(17), Co => CTMP_18_port);
   FAI_19 : FA_1390 port map( A => A(18), B => B(18), Ci => CTMP_18_port, S => 
                           S(18), Co => CTMP_19_port);
   FAI_20 : FA_1389 port map( A => A(19), B => B(19), Ci => CTMP_19_port, S => 
                           S(19), Co => CTMP_20_port);
   FAI_21 : FA_1388 port map( A => A(20), B => B(20), Ci => CTMP_20_port, S => 
                           S(20), Co => CTMP_21_port);
   FAI_22 : FA_1387 port map( A => A(21), B => B(21), Ci => CTMP_21_port, S => 
                           S(21), Co => CTMP_22_port);
   FAI_23 : FA_1386 port map( A => A(22), B => B(22), Ci => CTMP_22_port, S => 
                           S(22), Co => CTMP_23_port);
   FAI_24 : FA_1385 port map( A => A(23), B => B(23), Ci => CTMP_23_port, S => 
                           S(23), Co => CTMP_24_port);
   FAI_25 : FA_1384 port map( A => A(24), B => B(24), Ci => CTMP_24_port, S => 
                           S(24), Co => CTMP_25_port);
   FAI_26 : FA_1383 port map( A => A(25), B => B(25), Ci => CTMP_25_port, S => 
                           S(25), Co => CTMP_26_port);
   FAI_27 : FA_1382 port map( A => A(26), B => B(26), Ci => CTMP_26_port, S => 
                           S(26), Co => CTMP_27_port);
   FAI_28 : FA_1381 port map( A => A(27), B => B(27), Ci => CTMP_27_port, S => 
                           S(27), Co => CTMP_28_port);
   FAI_29 : FA_1380 port map( A => A(28), B => B(28), Ci => CTMP_28_port, S => 
                           S(28), Co => CTMP_29_port);
   FAI_30 : FA_1379 port map( A => A(29), B => B(29), Ci => CTMP_29_port, S => 
                           S(29), Co => CTMP_30_port);
   FAI_31 : FA_1378 port map( A => A(30), B => B(30), Ci => CTMP_30_port, S => 
                           S(30), Co => CTMP_31_port);
   FAI_32 : FA_1377 port map( A => A(31), B => B(31), Ci => CTMP_31_port, S => 
                           S(31), Co => CTMP_32_port);
   FAI_33 : FA_1376 port map( A => A(32), B => B(32), Ci => CTMP_32_port, S => 
                           S(32), Co => CTMP_33_port);
   FAI_34 : FA_1375 port map( A => A(33), B => B(33), Ci => CTMP_33_port, S => 
                           S(33), Co => CTMP_34_port);
   FAI_35 : FA_1374 port map( A => A(34), B => B(34), Ci => CTMP_34_port, S => 
                           S(34), Co => CTMP_35_port);
   FAI_36 : FA_1373 port map( A => A(35), B => B(35), Ci => CTMP_35_port, S => 
                           S(35), Co => CTMP_36_port);
   FAI_37 : FA_1372 port map( A => A(36), B => B(36), Ci => CTMP_36_port, S => 
                           S(36), Co => CTMP_37_port);
   FAI_38 : FA_1371 port map( A => A(37), B => B(37), Ci => CTMP_37_port, S => 
                           S(37), Co => CTMP_38_port);
   FAI_39 : FA_1370 port map( A => A(38), B => B(38), Ci => CTMP_38_port, S => 
                           S(38), Co => CTMP_39_port);
   FAI_40 : FA_1369 port map( A => A(39), B => B(39), Ci => CTMP_39_port, S => 
                           S(39), Co => CTMP_40_port);
   FAI_41 : FA_1368 port map( A => A(40), B => B(40), Ci => CTMP_40_port, S => 
                           S(40), Co => CTMP_41_port);
   FAI_42 : FA_1367 port map( A => A(41), B => B(41), Ci => CTMP_41_port, S => 
                           S(41), Co => CTMP_42_port);
   FAI_43 : FA_1366 port map( A => A(42), B => B(42), Ci => CTMP_42_port, S => 
                           S(42), Co => CTMP_43_port);
   FAI_44 : FA_1365 port map( A => A(43), B => B(43), Ci => CTMP_43_port, S => 
                           S(43), Co => CTMP_44_port);
   FAI_45 : FA_1364 port map( A => A(44), B => B(44), Ci => CTMP_44_port, S => 
                           S(44), Co => CTMP_45_port);
   FAI_46 : FA_1363 port map( A => A(45), B => B(45), Ci => CTMP_45_port, S => 
                           S(45), Co => CTMP_46_port);
   FAI_47 : FA_1362 port map( A => A(46), B => B(46), Ci => CTMP_46_port, S => 
                           S(46), Co => CTMP_47_port);
   FAI_48 : FA_1361 port map( A => A(47), B => B(47), Ci => CTMP_47_port, S => 
                           S(47), Co => CTMP_48_port);
   FAI_49 : FA_1360 port map( A => A(48), B => B(48), Ci => CTMP_48_port, S => 
                           S(48), Co => CTMP_49_port);
   FAI_50 : FA_1359 port map( A => A(49), B => B(49), Ci => CTMP_49_port, S => 
                           S(49), Co => CTMP_50_port);
   FAI_51 : FA_1358 port map( A => A(50), B => B(50), Ci => CTMP_50_port, S => 
                           S(50), Co => CTMP_51_port);
   FAI_52 : FA_1357 port map( A => A(51), B => B(51), Ci => CTMP_51_port, S => 
                           S(51), Co => CTMP_52_port);
   FAI_53 : FA_1356 port map( A => A(52), B => B(52), Ci => CTMP_52_port, S => 
                           S(52), Co => CTMP_53_port);
   FAI_54 : FA_1355 port map( A => A(53), B => B(53), Ci => CTMP_53_port, S => 
                           S(53), Co => CTMP_54_port);
   FAI_55 : FA_1354 port map( A => A(54), B => B(54), Ci => CTMP_54_port, S => 
                           S(54), Co => CTMP_55_port);
   FAI_56 : FA_1353 port map( A => A(55), B => B(55), Ci => CTMP_55_port, S => 
                           S(55), Co => CTMP_56_port);
   FAI_57 : FA_1352 port map( A => A(56), B => B(56), Ci => CTMP_56_port, S => 
                           S(56), Co => CTMP_57_port);
   FAI_58 : FA_1351 port map( A => A(57), B => B(57), Ci => CTMP_57_port, S => 
                           S(57), Co => CTMP_58_port);
   FAI_59 : FA_1350 port map( A => A(58), B => B(58), Ci => CTMP_58_port, S => 
                           S(58), Co => CTMP_59_port);
   FAI_60 : FA_1349 port map( A => A(59), B => B(59), Ci => CTMP_59_port, S => 
                           S(59), Co => CTMP_60_port);
   FAI_61 : FA_1348 port map( A => A(60), B => B(60), Ci => CTMP_60_port, S => 
                           S(60), Co => CTMP_61_port);
   FAI_62 : FA_1347 port map( A => A(61), B => B(61), Ci => CTMP_61_port, S => 
                           S(61), Co => CTMP_62_port);
   FAI_63 : FA_1346 port map( A => A(62), B => B(62), Ci => CTMP_62_port, S => 
                           S(62), Co => CTMP_63_port);
   FAI_64 : FA_1345 port map( A => A(63), B => B(63), Ci => CTMP_63_port, S => 
                           S(63), Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity RCA_NbitRca64_21 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_NbitRca64_21;

architecture SYN_STRUCTURAL of RCA_NbitRca64_21 is

   component FA_1281
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1282
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1283
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1284
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1285
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1286
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1287
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1288
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1289
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1290
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1291
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1292
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1293
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1294
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1295
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1296
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1297
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1298
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1299
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1300
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1301
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1302
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1303
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1304
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1305
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1306
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1307
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1308
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1309
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1310
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1311
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1312
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1313
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1314
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1315
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1316
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1317
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1318
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1319
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1320
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1321
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1322
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1323
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1324
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1325
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1326
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1327
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1328
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1329
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1330
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1331
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1332
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1333
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1334
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1335
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1336
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1337
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1338
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1339
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1340
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1341
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1342
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1343
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1344
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_63_port, CTMP_62_port, CTMP_61_port, CTMP_60_port, CTMP_59_port,
      CTMP_58_port, CTMP_57_port, CTMP_56_port, CTMP_55_port, CTMP_54_port, 
      CTMP_53_port, CTMP_52_port, CTMP_51_port, CTMP_50_port, CTMP_49_port, 
      CTMP_48_port, CTMP_47_port, CTMP_46_port, CTMP_45_port, CTMP_44_port, 
      CTMP_43_port, CTMP_42_port, CTMP_41_port, CTMP_40_port, CTMP_39_port, 
      CTMP_38_port, CTMP_37_port, CTMP_36_port, CTMP_35_port, CTMP_34_port, 
      CTMP_33_port, CTMP_32_port, CTMP_31_port, CTMP_30_port, CTMP_29_port, 
      CTMP_28_port, CTMP_27_port, CTMP_26_port, CTMP_25_port, CTMP_24_port, 
      CTMP_23_port, CTMP_22_port, CTMP_21_port, CTMP_20_port, CTMP_19_port, 
      CTMP_18_port, CTMP_17_port, CTMP_16_port, CTMP_15_port, CTMP_14_port, 
      CTMP_13_port, CTMP_12_port, CTMP_11_port, CTMP_10_port, CTMP_9_port, 
      CTMP_8_port, CTMP_7_port, CTMP_6_port, CTMP_5_port, CTMP_4_port, 
      CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_1344 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_1343 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1)
                           , Co => CTMP_2_port);
   FAI_3 : FA_1342 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2)
                           , Co => CTMP_3_port);
   FAI_4 : FA_1341 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3)
                           , Co => CTMP_4_port);
   FAI_5 : FA_1340 port map( A => A(4), B => B(4), Ci => CTMP_4_port, S => S(4)
                           , Co => CTMP_5_port);
   FAI_6 : FA_1339 port map( A => A(5), B => B(5), Ci => CTMP_5_port, S => S(5)
                           , Co => CTMP_6_port);
   FAI_7 : FA_1338 port map( A => A(6), B => B(6), Ci => CTMP_6_port, S => S(6)
                           , Co => CTMP_7_port);
   FAI_8 : FA_1337 port map( A => A(7), B => B(7), Ci => CTMP_7_port, S => S(7)
                           , Co => CTMP_8_port);
   FAI_9 : FA_1336 port map( A => A(8), B => B(8), Ci => CTMP_8_port, S => S(8)
                           , Co => CTMP_9_port);
   FAI_10 : FA_1335 port map( A => A(9), B => B(9), Ci => CTMP_9_port, S => 
                           S(9), Co => CTMP_10_port);
   FAI_11 : FA_1334 port map( A => A(10), B => B(10), Ci => CTMP_10_port, S => 
                           S(10), Co => CTMP_11_port);
   FAI_12 : FA_1333 port map( A => A(11), B => B(11), Ci => CTMP_11_port, S => 
                           S(11), Co => CTMP_12_port);
   FAI_13 : FA_1332 port map( A => A(12), B => B(12), Ci => CTMP_12_port, S => 
                           S(12), Co => CTMP_13_port);
   FAI_14 : FA_1331 port map( A => A(13), B => B(13), Ci => CTMP_13_port, S => 
                           S(13), Co => CTMP_14_port);
   FAI_15 : FA_1330 port map( A => A(14), B => B(14), Ci => CTMP_14_port, S => 
                           S(14), Co => CTMP_15_port);
   FAI_16 : FA_1329 port map( A => A(15), B => B(15), Ci => CTMP_15_port, S => 
                           S(15), Co => CTMP_16_port);
   FAI_17 : FA_1328 port map( A => A(16), B => B(16), Ci => CTMP_16_port, S => 
                           S(16), Co => CTMP_17_port);
   FAI_18 : FA_1327 port map( A => A(17), B => B(17), Ci => CTMP_17_port, S => 
                           S(17), Co => CTMP_18_port);
   FAI_19 : FA_1326 port map( A => A(18), B => B(18), Ci => CTMP_18_port, S => 
                           S(18), Co => CTMP_19_port);
   FAI_20 : FA_1325 port map( A => A(19), B => B(19), Ci => CTMP_19_port, S => 
                           S(19), Co => CTMP_20_port);
   FAI_21 : FA_1324 port map( A => A(20), B => B(20), Ci => CTMP_20_port, S => 
                           S(20), Co => CTMP_21_port);
   FAI_22 : FA_1323 port map( A => A(21), B => B(21), Ci => CTMP_21_port, S => 
                           S(21), Co => CTMP_22_port);
   FAI_23 : FA_1322 port map( A => A(22), B => B(22), Ci => CTMP_22_port, S => 
                           S(22), Co => CTMP_23_port);
   FAI_24 : FA_1321 port map( A => A(23), B => B(23), Ci => CTMP_23_port, S => 
                           S(23), Co => CTMP_24_port);
   FAI_25 : FA_1320 port map( A => A(24), B => B(24), Ci => CTMP_24_port, S => 
                           S(24), Co => CTMP_25_port);
   FAI_26 : FA_1319 port map( A => A(25), B => B(25), Ci => CTMP_25_port, S => 
                           S(25), Co => CTMP_26_port);
   FAI_27 : FA_1318 port map( A => A(26), B => B(26), Ci => CTMP_26_port, S => 
                           S(26), Co => CTMP_27_port);
   FAI_28 : FA_1317 port map( A => A(27), B => B(27), Ci => CTMP_27_port, S => 
                           S(27), Co => CTMP_28_port);
   FAI_29 : FA_1316 port map( A => A(28), B => B(28), Ci => CTMP_28_port, S => 
                           S(28), Co => CTMP_29_port);
   FAI_30 : FA_1315 port map( A => A(29), B => B(29), Ci => CTMP_29_port, S => 
                           S(29), Co => CTMP_30_port);
   FAI_31 : FA_1314 port map( A => A(30), B => B(30), Ci => CTMP_30_port, S => 
                           S(30), Co => CTMP_31_port);
   FAI_32 : FA_1313 port map( A => A(31), B => B(31), Ci => CTMP_31_port, S => 
                           S(31), Co => CTMP_32_port);
   FAI_33 : FA_1312 port map( A => A(32), B => B(32), Ci => CTMP_32_port, S => 
                           S(32), Co => CTMP_33_port);
   FAI_34 : FA_1311 port map( A => A(33), B => B(33), Ci => CTMP_33_port, S => 
                           S(33), Co => CTMP_34_port);
   FAI_35 : FA_1310 port map( A => A(34), B => B(34), Ci => CTMP_34_port, S => 
                           S(34), Co => CTMP_35_port);
   FAI_36 : FA_1309 port map( A => A(35), B => B(35), Ci => CTMP_35_port, S => 
                           S(35), Co => CTMP_36_port);
   FAI_37 : FA_1308 port map( A => A(36), B => B(36), Ci => CTMP_36_port, S => 
                           S(36), Co => CTMP_37_port);
   FAI_38 : FA_1307 port map( A => A(37), B => B(37), Ci => CTMP_37_port, S => 
                           S(37), Co => CTMP_38_port);
   FAI_39 : FA_1306 port map( A => A(38), B => B(38), Ci => CTMP_38_port, S => 
                           S(38), Co => CTMP_39_port);
   FAI_40 : FA_1305 port map( A => A(39), B => B(39), Ci => CTMP_39_port, S => 
                           S(39), Co => CTMP_40_port);
   FAI_41 : FA_1304 port map( A => A(40), B => B(40), Ci => CTMP_40_port, S => 
                           S(40), Co => CTMP_41_port);
   FAI_42 : FA_1303 port map( A => A(41), B => B(41), Ci => CTMP_41_port, S => 
                           S(41), Co => CTMP_42_port);
   FAI_43 : FA_1302 port map( A => A(42), B => B(42), Ci => CTMP_42_port, S => 
                           S(42), Co => CTMP_43_port);
   FAI_44 : FA_1301 port map( A => A(43), B => B(43), Ci => CTMP_43_port, S => 
                           S(43), Co => CTMP_44_port);
   FAI_45 : FA_1300 port map( A => A(44), B => B(44), Ci => CTMP_44_port, S => 
                           S(44), Co => CTMP_45_port);
   FAI_46 : FA_1299 port map( A => A(45), B => B(45), Ci => CTMP_45_port, S => 
                           S(45), Co => CTMP_46_port);
   FAI_47 : FA_1298 port map( A => A(46), B => B(46), Ci => CTMP_46_port, S => 
                           S(46), Co => CTMP_47_port);
   FAI_48 : FA_1297 port map( A => A(47), B => B(47), Ci => CTMP_47_port, S => 
                           S(47), Co => CTMP_48_port);
   FAI_49 : FA_1296 port map( A => A(48), B => B(48), Ci => CTMP_48_port, S => 
                           S(48), Co => CTMP_49_port);
   FAI_50 : FA_1295 port map( A => A(49), B => B(49), Ci => CTMP_49_port, S => 
                           S(49), Co => CTMP_50_port);
   FAI_51 : FA_1294 port map( A => A(50), B => B(50), Ci => CTMP_50_port, S => 
                           S(50), Co => CTMP_51_port);
   FAI_52 : FA_1293 port map( A => A(51), B => B(51), Ci => CTMP_51_port, S => 
                           S(51), Co => CTMP_52_port);
   FAI_53 : FA_1292 port map( A => A(52), B => B(52), Ci => CTMP_52_port, S => 
                           S(52), Co => CTMP_53_port);
   FAI_54 : FA_1291 port map( A => A(53), B => B(53), Ci => CTMP_53_port, S => 
                           S(53), Co => CTMP_54_port);
   FAI_55 : FA_1290 port map( A => A(54), B => B(54), Ci => CTMP_54_port, S => 
                           S(54), Co => CTMP_55_port);
   FAI_56 : FA_1289 port map( A => A(55), B => B(55), Ci => CTMP_55_port, S => 
                           S(55), Co => CTMP_56_port);
   FAI_57 : FA_1288 port map( A => A(56), B => B(56), Ci => CTMP_56_port, S => 
                           S(56), Co => CTMP_57_port);
   FAI_58 : FA_1287 port map( A => A(57), B => B(57), Ci => CTMP_57_port, S => 
                           S(57), Co => CTMP_58_port);
   FAI_59 : FA_1286 port map( A => A(58), B => B(58), Ci => CTMP_58_port, S => 
                           S(58), Co => CTMP_59_port);
   FAI_60 : FA_1285 port map( A => A(59), B => B(59), Ci => CTMP_59_port, S => 
                           S(59), Co => CTMP_60_port);
   FAI_61 : FA_1284 port map( A => A(60), B => B(60), Ci => CTMP_60_port, S => 
                           S(60), Co => CTMP_61_port);
   FAI_62 : FA_1283 port map( A => A(61), B => B(61), Ci => CTMP_61_port, S => 
                           S(61), Co => CTMP_62_port);
   FAI_63 : FA_1282 port map( A => A(62), B => B(62), Ci => CTMP_62_port, S => 
                           S(62), Co => CTMP_63_port);
   FAI_64 : FA_1281 port map( A => A(63), B => B(63), Ci => CTMP_63_port, S => 
                           S(63), Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity RCA_NbitRca64_20 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_NbitRca64_20;

architecture SYN_STRUCTURAL of RCA_NbitRca64_20 is

   component FA_1217
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1218
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1219
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1220
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1221
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1222
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1223
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1224
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1225
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1226
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1227
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1228
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1229
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1230
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1231
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1232
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1233
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1234
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1235
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1236
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1237
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1238
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1239
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1240
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1241
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1242
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1243
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1244
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1245
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1246
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1247
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1248
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1249
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1250
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1251
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1252
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1253
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1254
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1255
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1256
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1257
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1258
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1259
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1260
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1261
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1262
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1263
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1264
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1265
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1266
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1267
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1268
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1269
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1270
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1271
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1272
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1273
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1274
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1275
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1276
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1277
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1278
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1279
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1280
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_63_port, CTMP_62_port, CTMP_61_port, CTMP_60_port, CTMP_59_port,
      CTMP_58_port, CTMP_57_port, CTMP_56_port, CTMP_55_port, CTMP_54_port, 
      CTMP_53_port, CTMP_52_port, CTMP_51_port, CTMP_50_port, CTMP_49_port, 
      CTMP_48_port, CTMP_47_port, CTMP_46_port, CTMP_45_port, CTMP_44_port, 
      CTMP_43_port, CTMP_42_port, CTMP_41_port, CTMP_40_port, CTMP_39_port, 
      CTMP_38_port, CTMP_37_port, CTMP_36_port, CTMP_35_port, CTMP_34_port, 
      CTMP_33_port, CTMP_32_port, CTMP_31_port, CTMP_30_port, CTMP_29_port, 
      CTMP_28_port, CTMP_27_port, CTMP_26_port, CTMP_25_port, CTMP_24_port, 
      CTMP_23_port, CTMP_22_port, CTMP_21_port, CTMP_20_port, CTMP_19_port, 
      CTMP_18_port, CTMP_17_port, CTMP_16_port, CTMP_15_port, CTMP_14_port, 
      CTMP_13_port, CTMP_12_port, CTMP_11_port, CTMP_10_port, CTMP_9_port, 
      CTMP_8_port, CTMP_7_port, CTMP_6_port, CTMP_5_port, CTMP_4_port, 
      CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_1280 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_1279 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1)
                           , Co => CTMP_2_port);
   FAI_3 : FA_1278 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2)
                           , Co => CTMP_3_port);
   FAI_4 : FA_1277 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3)
                           , Co => CTMP_4_port);
   FAI_5 : FA_1276 port map( A => A(4), B => B(4), Ci => CTMP_4_port, S => S(4)
                           , Co => CTMP_5_port);
   FAI_6 : FA_1275 port map( A => A(5), B => B(5), Ci => CTMP_5_port, S => S(5)
                           , Co => CTMP_6_port);
   FAI_7 : FA_1274 port map( A => A(6), B => B(6), Ci => CTMP_6_port, S => S(6)
                           , Co => CTMP_7_port);
   FAI_8 : FA_1273 port map( A => A(7), B => B(7), Ci => CTMP_7_port, S => S(7)
                           , Co => CTMP_8_port);
   FAI_9 : FA_1272 port map( A => A(8), B => B(8), Ci => CTMP_8_port, S => S(8)
                           , Co => CTMP_9_port);
   FAI_10 : FA_1271 port map( A => A(9), B => B(9), Ci => CTMP_9_port, S => 
                           S(9), Co => CTMP_10_port);
   FAI_11 : FA_1270 port map( A => A(10), B => B(10), Ci => CTMP_10_port, S => 
                           S(10), Co => CTMP_11_port);
   FAI_12 : FA_1269 port map( A => A(11), B => B(11), Ci => CTMP_11_port, S => 
                           S(11), Co => CTMP_12_port);
   FAI_13 : FA_1268 port map( A => A(12), B => B(12), Ci => CTMP_12_port, S => 
                           S(12), Co => CTMP_13_port);
   FAI_14 : FA_1267 port map( A => A(13), B => B(13), Ci => CTMP_13_port, S => 
                           S(13), Co => CTMP_14_port);
   FAI_15 : FA_1266 port map( A => A(14), B => B(14), Ci => CTMP_14_port, S => 
                           S(14), Co => CTMP_15_port);
   FAI_16 : FA_1265 port map( A => A(15), B => B(15), Ci => CTMP_15_port, S => 
                           S(15), Co => CTMP_16_port);
   FAI_17 : FA_1264 port map( A => A(16), B => B(16), Ci => CTMP_16_port, S => 
                           S(16), Co => CTMP_17_port);
   FAI_18 : FA_1263 port map( A => A(17), B => B(17), Ci => CTMP_17_port, S => 
                           S(17), Co => CTMP_18_port);
   FAI_19 : FA_1262 port map( A => A(18), B => B(18), Ci => CTMP_18_port, S => 
                           S(18), Co => CTMP_19_port);
   FAI_20 : FA_1261 port map( A => A(19), B => B(19), Ci => CTMP_19_port, S => 
                           S(19), Co => CTMP_20_port);
   FAI_21 : FA_1260 port map( A => A(20), B => B(20), Ci => CTMP_20_port, S => 
                           S(20), Co => CTMP_21_port);
   FAI_22 : FA_1259 port map( A => A(21), B => B(21), Ci => CTMP_21_port, S => 
                           S(21), Co => CTMP_22_port);
   FAI_23 : FA_1258 port map( A => A(22), B => B(22), Ci => CTMP_22_port, S => 
                           S(22), Co => CTMP_23_port);
   FAI_24 : FA_1257 port map( A => A(23), B => B(23), Ci => CTMP_23_port, S => 
                           S(23), Co => CTMP_24_port);
   FAI_25 : FA_1256 port map( A => A(24), B => B(24), Ci => CTMP_24_port, S => 
                           S(24), Co => CTMP_25_port);
   FAI_26 : FA_1255 port map( A => A(25), B => B(25), Ci => CTMP_25_port, S => 
                           S(25), Co => CTMP_26_port);
   FAI_27 : FA_1254 port map( A => A(26), B => B(26), Ci => CTMP_26_port, S => 
                           S(26), Co => CTMP_27_port);
   FAI_28 : FA_1253 port map( A => A(27), B => B(27), Ci => CTMP_27_port, S => 
                           S(27), Co => CTMP_28_port);
   FAI_29 : FA_1252 port map( A => A(28), B => B(28), Ci => CTMP_28_port, S => 
                           S(28), Co => CTMP_29_port);
   FAI_30 : FA_1251 port map( A => A(29), B => B(29), Ci => CTMP_29_port, S => 
                           S(29), Co => CTMP_30_port);
   FAI_31 : FA_1250 port map( A => A(30), B => B(30), Ci => CTMP_30_port, S => 
                           S(30), Co => CTMP_31_port);
   FAI_32 : FA_1249 port map( A => A(31), B => B(31), Ci => CTMP_31_port, S => 
                           S(31), Co => CTMP_32_port);
   FAI_33 : FA_1248 port map( A => A(32), B => B(32), Ci => CTMP_32_port, S => 
                           S(32), Co => CTMP_33_port);
   FAI_34 : FA_1247 port map( A => A(33), B => B(33), Ci => CTMP_33_port, S => 
                           S(33), Co => CTMP_34_port);
   FAI_35 : FA_1246 port map( A => A(34), B => B(34), Ci => CTMP_34_port, S => 
                           S(34), Co => CTMP_35_port);
   FAI_36 : FA_1245 port map( A => A(35), B => B(35), Ci => CTMP_35_port, S => 
                           S(35), Co => CTMP_36_port);
   FAI_37 : FA_1244 port map( A => A(36), B => B(36), Ci => CTMP_36_port, S => 
                           S(36), Co => CTMP_37_port);
   FAI_38 : FA_1243 port map( A => A(37), B => B(37), Ci => CTMP_37_port, S => 
                           S(37), Co => CTMP_38_port);
   FAI_39 : FA_1242 port map( A => A(38), B => B(38), Ci => CTMP_38_port, S => 
                           S(38), Co => CTMP_39_port);
   FAI_40 : FA_1241 port map( A => A(39), B => B(39), Ci => CTMP_39_port, S => 
                           S(39), Co => CTMP_40_port);
   FAI_41 : FA_1240 port map( A => A(40), B => B(40), Ci => CTMP_40_port, S => 
                           S(40), Co => CTMP_41_port);
   FAI_42 : FA_1239 port map( A => A(41), B => B(41), Ci => CTMP_41_port, S => 
                           S(41), Co => CTMP_42_port);
   FAI_43 : FA_1238 port map( A => A(42), B => B(42), Ci => CTMP_42_port, S => 
                           S(42), Co => CTMP_43_port);
   FAI_44 : FA_1237 port map( A => A(43), B => B(43), Ci => CTMP_43_port, S => 
                           S(43), Co => CTMP_44_port);
   FAI_45 : FA_1236 port map( A => A(44), B => B(44), Ci => CTMP_44_port, S => 
                           S(44), Co => CTMP_45_port);
   FAI_46 : FA_1235 port map( A => A(45), B => B(45), Ci => CTMP_45_port, S => 
                           S(45), Co => CTMP_46_port);
   FAI_47 : FA_1234 port map( A => A(46), B => B(46), Ci => CTMP_46_port, S => 
                           S(46), Co => CTMP_47_port);
   FAI_48 : FA_1233 port map( A => A(47), B => B(47), Ci => CTMP_47_port, S => 
                           S(47), Co => CTMP_48_port);
   FAI_49 : FA_1232 port map( A => A(48), B => B(48), Ci => CTMP_48_port, S => 
                           S(48), Co => CTMP_49_port);
   FAI_50 : FA_1231 port map( A => A(49), B => B(49), Ci => CTMP_49_port, S => 
                           S(49), Co => CTMP_50_port);
   FAI_51 : FA_1230 port map( A => A(50), B => B(50), Ci => CTMP_50_port, S => 
                           S(50), Co => CTMP_51_port);
   FAI_52 : FA_1229 port map( A => A(51), B => B(51), Ci => CTMP_51_port, S => 
                           S(51), Co => CTMP_52_port);
   FAI_53 : FA_1228 port map( A => A(52), B => B(52), Ci => CTMP_52_port, S => 
                           S(52), Co => CTMP_53_port);
   FAI_54 : FA_1227 port map( A => A(53), B => B(53), Ci => CTMP_53_port, S => 
                           S(53), Co => CTMP_54_port);
   FAI_55 : FA_1226 port map( A => A(54), B => B(54), Ci => CTMP_54_port, S => 
                           S(54), Co => CTMP_55_port);
   FAI_56 : FA_1225 port map( A => A(55), B => B(55), Ci => CTMP_55_port, S => 
                           S(55), Co => CTMP_56_port);
   FAI_57 : FA_1224 port map( A => A(56), B => B(56), Ci => CTMP_56_port, S => 
                           S(56), Co => CTMP_57_port);
   FAI_58 : FA_1223 port map( A => A(57), B => B(57), Ci => CTMP_57_port, S => 
                           S(57), Co => CTMP_58_port);
   FAI_59 : FA_1222 port map( A => A(58), B => B(58), Ci => CTMP_58_port, S => 
                           S(58), Co => CTMP_59_port);
   FAI_60 : FA_1221 port map( A => A(59), B => B(59), Ci => CTMP_59_port, S => 
                           S(59), Co => CTMP_60_port);
   FAI_61 : FA_1220 port map( A => A(60), B => B(60), Ci => CTMP_60_port, S => 
                           S(60), Co => CTMP_61_port);
   FAI_62 : FA_1219 port map( A => A(61), B => B(61), Ci => CTMP_61_port, S => 
                           S(61), Co => CTMP_62_port);
   FAI_63 : FA_1218 port map( A => A(62), B => B(62), Ci => CTMP_62_port, S => 
                           S(62), Co => CTMP_63_port);
   FAI_64 : FA_1217 port map( A => A(63), B => B(63), Ci => CTMP_63_port, S => 
                           S(63), Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity RCA_NbitRca64_19 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_NbitRca64_19;

architecture SYN_STRUCTURAL of RCA_NbitRca64_19 is

   component FA_1153
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1154
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1155
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1156
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1157
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1158
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1159
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1160
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1161
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1162
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1163
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1164
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1165
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1166
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1167
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1168
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1169
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1170
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1171
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1172
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1173
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1174
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1175
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1176
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1177
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1178
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1179
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1180
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1181
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1182
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1183
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1184
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1185
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1186
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1187
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1188
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1189
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1190
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1191
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1192
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1193
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1194
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1195
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1196
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1197
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1198
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1199
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1200
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1201
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1202
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1203
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1204
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1205
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1206
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1207
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1208
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1209
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1210
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1211
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1212
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1213
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1214
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1215
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1216
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_63_port, CTMP_62_port, CTMP_61_port, CTMP_60_port, CTMP_59_port,
      CTMP_58_port, CTMP_57_port, CTMP_56_port, CTMP_55_port, CTMP_54_port, 
      CTMP_53_port, CTMP_52_port, CTMP_51_port, CTMP_50_port, CTMP_49_port, 
      CTMP_48_port, CTMP_47_port, CTMP_46_port, CTMP_45_port, CTMP_44_port, 
      CTMP_43_port, CTMP_42_port, CTMP_41_port, CTMP_40_port, CTMP_39_port, 
      CTMP_38_port, CTMP_37_port, CTMP_36_port, CTMP_35_port, CTMP_34_port, 
      CTMP_33_port, CTMP_32_port, CTMP_31_port, CTMP_30_port, CTMP_29_port, 
      CTMP_28_port, CTMP_27_port, CTMP_26_port, CTMP_25_port, CTMP_24_port, 
      CTMP_23_port, CTMP_22_port, CTMP_21_port, CTMP_20_port, CTMP_19_port, 
      CTMP_18_port, CTMP_17_port, CTMP_16_port, CTMP_15_port, CTMP_14_port, 
      CTMP_13_port, CTMP_12_port, CTMP_11_port, CTMP_10_port, CTMP_9_port, 
      CTMP_8_port, CTMP_7_port, CTMP_6_port, CTMP_5_port, CTMP_4_port, 
      CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_1216 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_1215 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1)
                           , Co => CTMP_2_port);
   FAI_3 : FA_1214 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2)
                           , Co => CTMP_3_port);
   FAI_4 : FA_1213 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3)
                           , Co => CTMP_4_port);
   FAI_5 : FA_1212 port map( A => A(4), B => B(4), Ci => CTMP_4_port, S => S(4)
                           , Co => CTMP_5_port);
   FAI_6 : FA_1211 port map( A => A(5), B => B(5), Ci => CTMP_5_port, S => S(5)
                           , Co => CTMP_6_port);
   FAI_7 : FA_1210 port map( A => A(6), B => B(6), Ci => CTMP_6_port, S => S(6)
                           , Co => CTMP_7_port);
   FAI_8 : FA_1209 port map( A => A(7), B => B(7), Ci => CTMP_7_port, S => S(7)
                           , Co => CTMP_8_port);
   FAI_9 : FA_1208 port map( A => A(8), B => B(8), Ci => CTMP_8_port, S => S(8)
                           , Co => CTMP_9_port);
   FAI_10 : FA_1207 port map( A => A(9), B => B(9), Ci => CTMP_9_port, S => 
                           S(9), Co => CTMP_10_port);
   FAI_11 : FA_1206 port map( A => A(10), B => B(10), Ci => CTMP_10_port, S => 
                           S(10), Co => CTMP_11_port);
   FAI_12 : FA_1205 port map( A => A(11), B => B(11), Ci => CTMP_11_port, S => 
                           S(11), Co => CTMP_12_port);
   FAI_13 : FA_1204 port map( A => A(12), B => B(12), Ci => CTMP_12_port, S => 
                           S(12), Co => CTMP_13_port);
   FAI_14 : FA_1203 port map( A => A(13), B => B(13), Ci => CTMP_13_port, S => 
                           S(13), Co => CTMP_14_port);
   FAI_15 : FA_1202 port map( A => A(14), B => B(14), Ci => CTMP_14_port, S => 
                           S(14), Co => CTMP_15_port);
   FAI_16 : FA_1201 port map( A => A(15), B => B(15), Ci => CTMP_15_port, S => 
                           S(15), Co => CTMP_16_port);
   FAI_17 : FA_1200 port map( A => A(16), B => B(16), Ci => CTMP_16_port, S => 
                           S(16), Co => CTMP_17_port);
   FAI_18 : FA_1199 port map( A => A(17), B => B(17), Ci => CTMP_17_port, S => 
                           S(17), Co => CTMP_18_port);
   FAI_19 : FA_1198 port map( A => A(18), B => B(18), Ci => CTMP_18_port, S => 
                           S(18), Co => CTMP_19_port);
   FAI_20 : FA_1197 port map( A => A(19), B => B(19), Ci => CTMP_19_port, S => 
                           S(19), Co => CTMP_20_port);
   FAI_21 : FA_1196 port map( A => A(20), B => B(20), Ci => CTMP_20_port, S => 
                           S(20), Co => CTMP_21_port);
   FAI_22 : FA_1195 port map( A => A(21), B => B(21), Ci => CTMP_21_port, S => 
                           S(21), Co => CTMP_22_port);
   FAI_23 : FA_1194 port map( A => A(22), B => B(22), Ci => CTMP_22_port, S => 
                           S(22), Co => CTMP_23_port);
   FAI_24 : FA_1193 port map( A => A(23), B => B(23), Ci => CTMP_23_port, S => 
                           S(23), Co => CTMP_24_port);
   FAI_25 : FA_1192 port map( A => A(24), B => B(24), Ci => CTMP_24_port, S => 
                           S(24), Co => CTMP_25_port);
   FAI_26 : FA_1191 port map( A => A(25), B => B(25), Ci => CTMP_25_port, S => 
                           S(25), Co => CTMP_26_port);
   FAI_27 : FA_1190 port map( A => A(26), B => B(26), Ci => CTMP_26_port, S => 
                           S(26), Co => CTMP_27_port);
   FAI_28 : FA_1189 port map( A => A(27), B => B(27), Ci => CTMP_27_port, S => 
                           S(27), Co => CTMP_28_port);
   FAI_29 : FA_1188 port map( A => A(28), B => B(28), Ci => CTMP_28_port, S => 
                           S(28), Co => CTMP_29_port);
   FAI_30 : FA_1187 port map( A => A(29), B => B(29), Ci => CTMP_29_port, S => 
                           S(29), Co => CTMP_30_port);
   FAI_31 : FA_1186 port map( A => A(30), B => B(30), Ci => CTMP_30_port, S => 
                           S(30), Co => CTMP_31_port);
   FAI_32 : FA_1185 port map( A => A(31), B => B(31), Ci => CTMP_31_port, S => 
                           S(31), Co => CTMP_32_port);
   FAI_33 : FA_1184 port map( A => A(32), B => B(32), Ci => CTMP_32_port, S => 
                           S(32), Co => CTMP_33_port);
   FAI_34 : FA_1183 port map( A => A(33), B => B(33), Ci => CTMP_33_port, S => 
                           S(33), Co => CTMP_34_port);
   FAI_35 : FA_1182 port map( A => A(34), B => B(34), Ci => CTMP_34_port, S => 
                           S(34), Co => CTMP_35_port);
   FAI_36 : FA_1181 port map( A => A(35), B => B(35), Ci => CTMP_35_port, S => 
                           S(35), Co => CTMP_36_port);
   FAI_37 : FA_1180 port map( A => A(36), B => B(36), Ci => CTMP_36_port, S => 
                           S(36), Co => CTMP_37_port);
   FAI_38 : FA_1179 port map( A => A(37), B => B(37), Ci => CTMP_37_port, S => 
                           S(37), Co => CTMP_38_port);
   FAI_39 : FA_1178 port map( A => A(38), B => B(38), Ci => CTMP_38_port, S => 
                           S(38), Co => CTMP_39_port);
   FAI_40 : FA_1177 port map( A => A(39), B => B(39), Ci => CTMP_39_port, S => 
                           S(39), Co => CTMP_40_port);
   FAI_41 : FA_1176 port map( A => A(40), B => B(40), Ci => CTMP_40_port, S => 
                           S(40), Co => CTMP_41_port);
   FAI_42 : FA_1175 port map( A => A(41), B => B(41), Ci => CTMP_41_port, S => 
                           S(41), Co => CTMP_42_port);
   FAI_43 : FA_1174 port map( A => A(42), B => B(42), Ci => CTMP_42_port, S => 
                           S(42), Co => CTMP_43_port);
   FAI_44 : FA_1173 port map( A => A(43), B => B(43), Ci => CTMP_43_port, S => 
                           S(43), Co => CTMP_44_port);
   FAI_45 : FA_1172 port map( A => A(44), B => B(44), Ci => CTMP_44_port, S => 
                           S(44), Co => CTMP_45_port);
   FAI_46 : FA_1171 port map( A => A(45), B => B(45), Ci => CTMP_45_port, S => 
                           S(45), Co => CTMP_46_port);
   FAI_47 : FA_1170 port map( A => A(46), B => B(46), Ci => CTMP_46_port, S => 
                           S(46), Co => CTMP_47_port);
   FAI_48 : FA_1169 port map( A => A(47), B => B(47), Ci => CTMP_47_port, S => 
                           S(47), Co => CTMP_48_port);
   FAI_49 : FA_1168 port map( A => A(48), B => B(48), Ci => CTMP_48_port, S => 
                           S(48), Co => CTMP_49_port);
   FAI_50 : FA_1167 port map( A => A(49), B => B(49), Ci => CTMP_49_port, S => 
                           S(49), Co => CTMP_50_port);
   FAI_51 : FA_1166 port map( A => A(50), B => B(50), Ci => CTMP_50_port, S => 
                           S(50), Co => CTMP_51_port);
   FAI_52 : FA_1165 port map( A => A(51), B => B(51), Ci => CTMP_51_port, S => 
                           S(51), Co => CTMP_52_port);
   FAI_53 : FA_1164 port map( A => A(52), B => B(52), Ci => CTMP_52_port, S => 
                           S(52), Co => CTMP_53_port);
   FAI_54 : FA_1163 port map( A => A(53), B => B(53), Ci => CTMP_53_port, S => 
                           S(53), Co => CTMP_54_port);
   FAI_55 : FA_1162 port map( A => A(54), B => B(54), Ci => CTMP_54_port, S => 
                           S(54), Co => CTMP_55_port);
   FAI_56 : FA_1161 port map( A => A(55), B => B(55), Ci => CTMP_55_port, S => 
                           S(55), Co => CTMP_56_port);
   FAI_57 : FA_1160 port map( A => A(56), B => B(56), Ci => CTMP_56_port, S => 
                           S(56), Co => CTMP_57_port);
   FAI_58 : FA_1159 port map( A => A(57), B => B(57), Ci => CTMP_57_port, S => 
                           S(57), Co => CTMP_58_port);
   FAI_59 : FA_1158 port map( A => A(58), B => B(58), Ci => CTMP_58_port, S => 
                           S(58), Co => CTMP_59_port);
   FAI_60 : FA_1157 port map( A => A(59), B => B(59), Ci => CTMP_59_port, S => 
                           S(59), Co => CTMP_60_port);
   FAI_61 : FA_1156 port map( A => A(60), B => B(60), Ci => CTMP_60_port, S => 
                           S(60), Co => CTMP_61_port);
   FAI_62 : FA_1155 port map( A => A(61), B => B(61), Ci => CTMP_61_port, S => 
                           S(61), Co => CTMP_62_port);
   FAI_63 : FA_1154 port map( A => A(62), B => B(62), Ci => CTMP_62_port, S => 
                           S(62), Co => CTMP_63_port);
   FAI_64 : FA_1153 port map( A => A(63), B => B(63), Ci => CTMP_63_port, S => 
                           S(63), Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity RCA_NbitRca64_18 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_NbitRca64_18;

architecture SYN_STRUCTURAL of RCA_NbitRca64_18 is

   component FA_1089
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1090
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1091
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1092
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1093
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1094
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1095
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1096
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1097
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1098
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1099
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1100
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1101
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1102
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1103
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1104
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1105
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1106
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1107
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1108
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1109
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1110
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1111
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1112
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1113
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1114
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1115
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1116
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1117
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1118
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1119
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1120
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1121
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1122
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1123
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1124
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1125
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1126
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1127
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1128
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1129
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1130
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1131
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1132
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1133
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1134
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1135
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1136
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1137
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1138
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1139
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1140
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1141
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1142
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1143
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1144
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1145
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1146
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1147
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1148
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1149
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1150
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1151
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1152
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_63_port, CTMP_62_port, CTMP_61_port, CTMP_60_port, CTMP_59_port,
      CTMP_58_port, CTMP_57_port, CTMP_56_port, CTMP_55_port, CTMP_54_port, 
      CTMP_53_port, CTMP_52_port, CTMP_51_port, CTMP_50_port, CTMP_49_port, 
      CTMP_48_port, CTMP_47_port, CTMP_46_port, CTMP_45_port, CTMP_44_port, 
      CTMP_43_port, CTMP_42_port, CTMP_41_port, CTMP_40_port, CTMP_39_port, 
      CTMP_38_port, CTMP_37_port, CTMP_36_port, CTMP_35_port, CTMP_34_port, 
      CTMP_33_port, CTMP_32_port, CTMP_31_port, CTMP_30_port, CTMP_29_port, 
      CTMP_28_port, CTMP_27_port, CTMP_26_port, CTMP_25_port, CTMP_24_port, 
      CTMP_23_port, CTMP_22_port, CTMP_21_port, CTMP_20_port, CTMP_19_port, 
      CTMP_18_port, CTMP_17_port, CTMP_16_port, CTMP_15_port, CTMP_14_port, 
      CTMP_13_port, CTMP_12_port, CTMP_11_port, CTMP_10_port, CTMP_9_port, 
      CTMP_8_port, CTMP_7_port, CTMP_6_port, CTMP_5_port, CTMP_4_port, 
      CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_1152 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_1151 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1)
                           , Co => CTMP_2_port);
   FAI_3 : FA_1150 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2)
                           , Co => CTMP_3_port);
   FAI_4 : FA_1149 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3)
                           , Co => CTMP_4_port);
   FAI_5 : FA_1148 port map( A => A(4), B => B(4), Ci => CTMP_4_port, S => S(4)
                           , Co => CTMP_5_port);
   FAI_6 : FA_1147 port map( A => A(5), B => B(5), Ci => CTMP_5_port, S => S(5)
                           , Co => CTMP_6_port);
   FAI_7 : FA_1146 port map( A => A(6), B => B(6), Ci => CTMP_6_port, S => S(6)
                           , Co => CTMP_7_port);
   FAI_8 : FA_1145 port map( A => A(7), B => B(7), Ci => CTMP_7_port, S => S(7)
                           , Co => CTMP_8_port);
   FAI_9 : FA_1144 port map( A => A(8), B => B(8), Ci => CTMP_8_port, S => S(8)
                           , Co => CTMP_9_port);
   FAI_10 : FA_1143 port map( A => A(9), B => B(9), Ci => CTMP_9_port, S => 
                           S(9), Co => CTMP_10_port);
   FAI_11 : FA_1142 port map( A => A(10), B => B(10), Ci => CTMP_10_port, S => 
                           S(10), Co => CTMP_11_port);
   FAI_12 : FA_1141 port map( A => A(11), B => B(11), Ci => CTMP_11_port, S => 
                           S(11), Co => CTMP_12_port);
   FAI_13 : FA_1140 port map( A => A(12), B => B(12), Ci => CTMP_12_port, S => 
                           S(12), Co => CTMP_13_port);
   FAI_14 : FA_1139 port map( A => A(13), B => B(13), Ci => CTMP_13_port, S => 
                           S(13), Co => CTMP_14_port);
   FAI_15 : FA_1138 port map( A => A(14), B => B(14), Ci => CTMP_14_port, S => 
                           S(14), Co => CTMP_15_port);
   FAI_16 : FA_1137 port map( A => A(15), B => B(15), Ci => CTMP_15_port, S => 
                           S(15), Co => CTMP_16_port);
   FAI_17 : FA_1136 port map( A => A(16), B => B(16), Ci => CTMP_16_port, S => 
                           S(16), Co => CTMP_17_port);
   FAI_18 : FA_1135 port map( A => A(17), B => B(17), Ci => CTMP_17_port, S => 
                           S(17), Co => CTMP_18_port);
   FAI_19 : FA_1134 port map( A => A(18), B => B(18), Ci => CTMP_18_port, S => 
                           S(18), Co => CTMP_19_port);
   FAI_20 : FA_1133 port map( A => A(19), B => B(19), Ci => CTMP_19_port, S => 
                           S(19), Co => CTMP_20_port);
   FAI_21 : FA_1132 port map( A => A(20), B => B(20), Ci => CTMP_20_port, S => 
                           S(20), Co => CTMP_21_port);
   FAI_22 : FA_1131 port map( A => A(21), B => B(21), Ci => CTMP_21_port, S => 
                           S(21), Co => CTMP_22_port);
   FAI_23 : FA_1130 port map( A => A(22), B => B(22), Ci => CTMP_22_port, S => 
                           S(22), Co => CTMP_23_port);
   FAI_24 : FA_1129 port map( A => A(23), B => B(23), Ci => CTMP_23_port, S => 
                           S(23), Co => CTMP_24_port);
   FAI_25 : FA_1128 port map( A => A(24), B => B(24), Ci => CTMP_24_port, S => 
                           S(24), Co => CTMP_25_port);
   FAI_26 : FA_1127 port map( A => A(25), B => B(25), Ci => CTMP_25_port, S => 
                           S(25), Co => CTMP_26_port);
   FAI_27 : FA_1126 port map( A => A(26), B => B(26), Ci => CTMP_26_port, S => 
                           S(26), Co => CTMP_27_port);
   FAI_28 : FA_1125 port map( A => A(27), B => B(27), Ci => CTMP_27_port, S => 
                           S(27), Co => CTMP_28_port);
   FAI_29 : FA_1124 port map( A => A(28), B => B(28), Ci => CTMP_28_port, S => 
                           S(28), Co => CTMP_29_port);
   FAI_30 : FA_1123 port map( A => A(29), B => B(29), Ci => CTMP_29_port, S => 
                           S(29), Co => CTMP_30_port);
   FAI_31 : FA_1122 port map( A => A(30), B => B(30), Ci => CTMP_30_port, S => 
                           S(30), Co => CTMP_31_port);
   FAI_32 : FA_1121 port map( A => A(31), B => B(31), Ci => CTMP_31_port, S => 
                           S(31), Co => CTMP_32_port);
   FAI_33 : FA_1120 port map( A => A(32), B => B(32), Ci => CTMP_32_port, S => 
                           S(32), Co => CTMP_33_port);
   FAI_34 : FA_1119 port map( A => A(33), B => B(33), Ci => CTMP_33_port, S => 
                           S(33), Co => CTMP_34_port);
   FAI_35 : FA_1118 port map( A => A(34), B => B(34), Ci => CTMP_34_port, S => 
                           S(34), Co => CTMP_35_port);
   FAI_36 : FA_1117 port map( A => A(35), B => B(35), Ci => CTMP_35_port, S => 
                           S(35), Co => CTMP_36_port);
   FAI_37 : FA_1116 port map( A => A(36), B => B(36), Ci => CTMP_36_port, S => 
                           S(36), Co => CTMP_37_port);
   FAI_38 : FA_1115 port map( A => A(37), B => B(37), Ci => CTMP_37_port, S => 
                           S(37), Co => CTMP_38_port);
   FAI_39 : FA_1114 port map( A => A(38), B => B(38), Ci => CTMP_38_port, S => 
                           S(38), Co => CTMP_39_port);
   FAI_40 : FA_1113 port map( A => A(39), B => B(39), Ci => CTMP_39_port, S => 
                           S(39), Co => CTMP_40_port);
   FAI_41 : FA_1112 port map( A => A(40), B => B(40), Ci => CTMP_40_port, S => 
                           S(40), Co => CTMP_41_port);
   FAI_42 : FA_1111 port map( A => A(41), B => B(41), Ci => CTMP_41_port, S => 
                           S(41), Co => CTMP_42_port);
   FAI_43 : FA_1110 port map( A => A(42), B => B(42), Ci => CTMP_42_port, S => 
                           S(42), Co => CTMP_43_port);
   FAI_44 : FA_1109 port map( A => A(43), B => B(43), Ci => CTMP_43_port, S => 
                           S(43), Co => CTMP_44_port);
   FAI_45 : FA_1108 port map( A => A(44), B => B(44), Ci => CTMP_44_port, S => 
                           S(44), Co => CTMP_45_port);
   FAI_46 : FA_1107 port map( A => A(45), B => B(45), Ci => CTMP_45_port, S => 
                           S(45), Co => CTMP_46_port);
   FAI_47 : FA_1106 port map( A => A(46), B => B(46), Ci => CTMP_46_port, S => 
                           S(46), Co => CTMP_47_port);
   FAI_48 : FA_1105 port map( A => A(47), B => B(47), Ci => CTMP_47_port, S => 
                           S(47), Co => CTMP_48_port);
   FAI_49 : FA_1104 port map( A => A(48), B => B(48), Ci => CTMP_48_port, S => 
                           S(48), Co => CTMP_49_port);
   FAI_50 : FA_1103 port map( A => A(49), B => B(49), Ci => CTMP_49_port, S => 
                           S(49), Co => CTMP_50_port);
   FAI_51 : FA_1102 port map( A => A(50), B => B(50), Ci => CTMP_50_port, S => 
                           S(50), Co => CTMP_51_port);
   FAI_52 : FA_1101 port map( A => A(51), B => B(51), Ci => CTMP_51_port, S => 
                           S(51), Co => CTMP_52_port);
   FAI_53 : FA_1100 port map( A => A(52), B => B(52), Ci => CTMP_52_port, S => 
                           S(52), Co => CTMP_53_port);
   FAI_54 : FA_1099 port map( A => A(53), B => B(53), Ci => CTMP_53_port, S => 
                           S(53), Co => CTMP_54_port);
   FAI_55 : FA_1098 port map( A => A(54), B => B(54), Ci => CTMP_54_port, S => 
                           S(54), Co => CTMP_55_port);
   FAI_56 : FA_1097 port map( A => A(55), B => B(55), Ci => CTMP_55_port, S => 
                           S(55), Co => CTMP_56_port);
   FAI_57 : FA_1096 port map( A => A(56), B => B(56), Ci => CTMP_56_port, S => 
                           S(56), Co => CTMP_57_port);
   FAI_58 : FA_1095 port map( A => A(57), B => B(57), Ci => CTMP_57_port, S => 
                           S(57), Co => CTMP_58_port);
   FAI_59 : FA_1094 port map( A => A(58), B => B(58), Ci => CTMP_58_port, S => 
                           S(58), Co => CTMP_59_port);
   FAI_60 : FA_1093 port map( A => A(59), B => B(59), Ci => CTMP_59_port, S => 
                           S(59), Co => CTMP_60_port);
   FAI_61 : FA_1092 port map( A => A(60), B => B(60), Ci => CTMP_60_port, S => 
                           S(60), Co => CTMP_61_port);
   FAI_62 : FA_1091 port map( A => A(61), B => B(61), Ci => CTMP_61_port, S => 
                           S(61), Co => CTMP_62_port);
   FAI_63 : FA_1090 port map( A => A(62), B => B(62), Ci => CTMP_62_port, S => 
                           S(62), Co => CTMP_63_port);
   FAI_64 : FA_1089 port map( A => A(63), B => B(63), Ci => CTMP_63_port, S => 
                           S(63), Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity RCA_NbitRca64_17 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_NbitRca64_17;

architecture SYN_STRUCTURAL of RCA_NbitRca64_17 is

   component FA_1025
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1026
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1027
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1028
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1029
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1030
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1031
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1032
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1033
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1034
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1035
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1036
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1037
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1038
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1039
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1040
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1041
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1042
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1043
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1044
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1045
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1046
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1047
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1048
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1049
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1050
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1051
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1052
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1053
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1054
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1055
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1056
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1057
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1058
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1059
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1060
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1061
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1062
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1063
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1064
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1065
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1066
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1067
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1068
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1069
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1070
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1071
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1072
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1073
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1074
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1075
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1076
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1077
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1078
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1079
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1080
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1081
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1082
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1083
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1084
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1085
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1086
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1087
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1088
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_63_port, CTMP_62_port, CTMP_61_port, CTMP_60_port, CTMP_59_port,
      CTMP_58_port, CTMP_57_port, CTMP_56_port, CTMP_55_port, CTMP_54_port, 
      CTMP_53_port, CTMP_52_port, CTMP_51_port, CTMP_50_port, CTMP_49_port, 
      CTMP_48_port, CTMP_47_port, CTMP_46_port, CTMP_45_port, CTMP_44_port, 
      CTMP_43_port, CTMP_42_port, CTMP_41_port, CTMP_40_port, CTMP_39_port, 
      CTMP_38_port, CTMP_37_port, CTMP_36_port, CTMP_35_port, CTMP_34_port, 
      CTMP_33_port, CTMP_32_port, CTMP_31_port, CTMP_30_port, CTMP_29_port, 
      CTMP_28_port, CTMP_27_port, CTMP_26_port, CTMP_25_port, CTMP_24_port, 
      CTMP_23_port, CTMP_22_port, CTMP_21_port, CTMP_20_port, CTMP_19_port, 
      CTMP_18_port, CTMP_17_port, CTMP_16_port, CTMP_15_port, CTMP_14_port, 
      CTMP_13_port, CTMP_12_port, CTMP_11_port, CTMP_10_port, CTMP_9_port, 
      CTMP_8_port, CTMP_7_port, CTMP_6_port, CTMP_5_port, CTMP_4_port, 
      CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_1088 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_1087 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1)
                           , Co => CTMP_2_port);
   FAI_3 : FA_1086 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2)
                           , Co => CTMP_3_port);
   FAI_4 : FA_1085 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3)
                           , Co => CTMP_4_port);
   FAI_5 : FA_1084 port map( A => A(4), B => B(4), Ci => CTMP_4_port, S => S(4)
                           , Co => CTMP_5_port);
   FAI_6 : FA_1083 port map( A => A(5), B => B(5), Ci => CTMP_5_port, S => S(5)
                           , Co => CTMP_6_port);
   FAI_7 : FA_1082 port map( A => A(6), B => B(6), Ci => CTMP_6_port, S => S(6)
                           , Co => CTMP_7_port);
   FAI_8 : FA_1081 port map( A => A(7), B => B(7), Ci => CTMP_7_port, S => S(7)
                           , Co => CTMP_8_port);
   FAI_9 : FA_1080 port map( A => A(8), B => B(8), Ci => CTMP_8_port, S => S(8)
                           , Co => CTMP_9_port);
   FAI_10 : FA_1079 port map( A => A(9), B => B(9), Ci => CTMP_9_port, S => 
                           S(9), Co => CTMP_10_port);
   FAI_11 : FA_1078 port map( A => A(10), B => B(10), Ci => CTMP_10_port, S => 
                           S(10), Co => CTMP_11_port);
   FAI_12 : FA_1077 port map( A => A(11), B => B(11), Ci => CTMP_11_port, S => 
                           S(11), Co => CTMP_12_port);
   FAI_13 : FA_1076 port map( A => A(12), B => B(12), Ci => CTMP_12_port, S => 
                           S(12), Co => CTMP_13_port);
   FAI_14 : FA_1075 port map( A => A(13), B => B(13), Ci => CTMP_13_port, S => 
                           S(13), Co => CTMP_14_port);
   FAI_15 : FA_1074 port map( A => A(14), B => B(14), Ci => CTMP_14_port, S => 
                           S(14), Co => CTMP_15_port);
   FAI_16 : FA_1073 port map( A => A(15), B => B(15), Ci => CTMP_15_port, S => 
                           S(15), Co => CTMP_16_port);
   FAI_17 : FA_1072 port map( A => A(16), B => B(16), Ci => CTMP_16_port, S => 
                           S(16), Co => CTMP_17_port);
   FAI_18 : FA_1071 port map( A => A(17), B => B(17), Ci => CTMP_17_port, S => 
                           S(17), Co => CTMP_18_port);
   FAI_19 : FA_1070 port map( A => A(18), B => B(18), Ci => CTMP_18_port, S => 
                           S(18), Co => CTMP_19_port);
   FAI_20 : FA_1069 port map( A => A(19), B => B(19), Ci => CTMP_19_port, S => 
                           S(19), Co => CTMP_20_port);
   FAI_21 : FA_1068 port map( A => A(20), B => B(20), Ci => CTMP_20_port, S => 
                           S(20), Co => CTMP_21_port);
   FAI_22 : FA_1067 port map( A => A(21), B => B(21), Ci => CTMP_21_port, S => 
                           S(21), Co => CTMP_22_port);
   FAI_23 : FA_1066 port map( A => A(22), B => B(22), Ci => CTMP_22_port, S => 
                           S(22), Co => CTMP_23_port);
   FAI_24 : FA_1065 port map( A => A(23), B => B(23), Ci => CTMP_23_port, S => 
                           S(23), Co => CTMP_24_port);
   FAI_25 : FA_1064 port map( A => A(24), B => B(24), Ci => CTMP_24_port, S => 
                           S(24), Co => CTMP_25_port);
   FAI_26 : FA_1063 port map( A => A(25), B => B(25), Ci => CTMP_25_port, S => 
                           S(25), Co => CTMP_26_port);
   FAI_27 : FA_1062 port map( A => A(26), B => B(26), Ci => CTMP_26_port, S => 
                           S(26), Co => CTMP_27_port);
   FAI_28 : FA_1061 port map( A => A(27), B => B(27), Ci => CTMP_27_port, S => 
                           S(27), Co => CTMP_28_port);
   FAI_29 : FA_1060 port map( A => A(28), B => B(28), Ci => CTMP_28_port, S => 
                           S(28), Co => CTMP_29_port);
   FAI_30 : FA_1059 port map( A => A(29), B => B(29), Ci => CTMP_29_port, S => 
                           S(29), Co => CTMP_30_port);
   FAI_31 : FA_1058 port map( A => A(30), B => B(30), Ci => CTMP_30_port, S => 
                           S(30), Co => CTMP_31_port);
   FAI_32 : FA_1057 port map( A => A(31), B => B(31), Ci => CTMP_31_port, S => 
                           S(31), Co => CTMP_32_port);
   FAI_33 : FA_1056 port map( A => A(32), B => B(32), Ci => CTMP_32_port, S => 
                           S(32), Co => CTMP_33_port);
   FAI_34 : FA_1055 port map( A => A(33), B => B(33), Ci => CTMP_33_port, S => 
                           S(33), Co => CTMP_34_port);
   FAI_35 : FA_1054 port map( A => A(34), B => B(34), Ci => CTMP_34_port, S => 
                           S(34), Co => CTMP_35_port);
   FAI_36 : FA_1053 port map( A => A(35), B => B(35), Ci => CTMP_35_port, S => 
                           S(35), Co => CTMP_36_port);
   FAI_37 : FA_1052 port map( A => A(36), B => B(36), Ci => CTMP_36_port, S => 
                           S(36), Co => CTMP_37_port);
   FAI_38 : FA_1051 port map( A => A(37), B => B(37), Ci => CTMP_37_port, S => 
                           S(37), Co => CTMP_38_port);
   FAI_39 : FA_1050 port map( A => A(38), B => B(38), Ci => CTMP_38_port, S => 
                           S(38), Co => CTMP_39_port);
   FAI_40 : FA_1049 port map( A => A(39), B => B(39), Ci => CTMP_39_port, S => 
                           S(39), Co => CTMP_40_port);
   FAI_41 : FA_1048 port map( A => A(40), B => B(40), Ci => CTMP_40_port, S => 
                           S(40), Co => CTMP_41_port);
   FAI_42 : FA_1047 port map( A => A(41), B => B(41), Ci => CTMP_41_port, S => 
                           S(41), Co => CTMP_42_port);
   FAI_43 : FA_1046 port map( A => A(42), B => B(42), Ci => CTMP_42_port, S => 
                           S(42), Co => CTMP_43_port);
   FAI_44 : FA_1045 port map( A => A(43), B => B(43), Ci => CTMP_43_port, S => 
                           S(43), Co => CTMP_44_port);
   FAI_45 : FA_1044 port map( A => A(44), B => B(44), Ci => CTMP_44_port, S => 
                           S(44), Co => CTMP_45_port);
   FAI_46 : FA_1043 port map( A => A(45), B => B(45), Ci => CTMP_45_port, S => 
                           S(45), Co => CTMP_46_port);
   FAI_47 : FA_1042 port map( A => A(46), B => B(46), Ci => CTMP_46_port, S => 
                           S(46), Co => CTMP_47_port);
   FAI_48 : FA_1041 port map( A => A(47), B => B(47), Ci => CTMP_47_port, S => 
                           S(47), Co => CTMP_48_port);
   FAI_49 : FA_1040 port map( A => A(48), B => B(48), Ci => CTMP_48_port, S => 
                           S(48), Co => CTMP_49_port);
   FAI_50 : FA_1039 port map( A => A(49), B => B(49), Ci => CTMP_49_port, S => 
                           S(49), Co => CTMP_50_port);
   FAI_51 : FA_1038 port map( A => A(50), B => B(50), Ci => CTMP_50_port, S => 
                           S(50), Co => CTMP_51_port);
   FAI_52 : FA_1037 port map( A => A(51), B => B(51), Ci => CTMP_51_port, S => 
                           S(51), Co => CTMP_52_port);
   FAI_53 : FA_1036 port map( A => A(52), B => B(52), Ci => CTMP_52_port, S => 
                           S(52), Co => CTMP_53_port);
   FAI_54 : FA_1035 port map( A => A(53), B => B(53), Ci => CTMP_53_port, S => 
                           S(53), Co => CTMP_54_port);
   FAI_55 : FA_1034 port map( A => A(54), B => B(54), Ci => CTMP_54_port, S => 
                           S(54), Co => CTMP_55_port);
   FAI_56 : FA_1033 port map( A => A(55), B => B(55), Ci => CTMP_55_port, S => 
                           S(55), Co => CTMP_56_port);
   FAI_57 : FA_1032 port map( A => A(56), B => B(56), Ci => CTMP_56_port, S => 
                           S(56), Co => CTMP_57_port);
   FAI_58 : FA_1031 port map( A => A(57), B => B(57), Ci => CTMP_57_port, S => 
                           S(57), Co => CTMP_58_port);
   FAI_59 : FA_1030 port map( A => A(58), B => B(58), Ci => CTMP_58_port, S => 
                           S(58), Co => CTMP_59_port);
   FAI_60 : FA_1029 port map( A => A(59), B => B(59), Ci => CTMP_59_port, S => 
                           S(59), Co => CTMP_60_port);
   FAI_61 : FA_1028 port map( A => A(60), B => B(60), Ci => CTMP_60_port, S => 
                           S(60), Co => CTMP_61_port);
   FAI_62 : FA_1027 port map( A => A(61), B => B(61), Ci => CTMP_61_port, S => 
                           S(61), Co => CTMP_62_port);
   FAI_63 : FA_1026 port map( A => A(62), B => B(62), Ci => CTMP_62_port, S => 
                           S(62), Co => CTMP_63_port);
   FAI_64 : FA_1025 port map( A => A(63), B => B(63), Ci => CTMP_63_port, S => 
                           S(63), Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity IV_127 is

   port( A : in std_logic;  Y : out std_logic);

end IV_127;

architecture SYN_BEHAVIORAL of IV_127 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity IV_126 is

   port( A : in std_logic;  Y : out std_logic);

end IV_126;

architecture SYN_BEHAVIORAL of IV_126 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity IV_125 is

   port( A : in std_logic;  Y : out std_logic);

end IV_125;

architecture SYN_BEHAVIORAL of IV_125 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity IV_124 is

   port( A : in std_logic;  Y : out std_logic);

end IV_124;

architecture SYN_BEHAVIORAL of IV_124 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity IV_123 is

   port( A : in std_logic;  Y : out std_logic);

end IV_123;

architecture SYN_BEHAVIORAL of IV_123 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity IV_122 is

   port( A : in std_logic;  Y : out std_logic);

end IV_122;

architecture SYN_BEHAVIORAL of IV_122 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity IV_121 is

   port( A : in std_logic;  Y : out std_logic);

end IV_121;

architecture SYN_BEHAVIORAL of IV_121 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity IV_120 is

   port( A : in std_logic;  Y : out std_logic);

end IV_120;

architecture SYN_BEHAVIORAL of IV_120 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity IV_119 is

   port( A : in std_logic;  Y : out std_logic);

end IV_119;

architecture SYN_BEHAVIORAL of IV_119 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity IV_118 is

   port( A : in std_logic;  Y : out std_logic);

end IV_118;

architecture SYN_BEHAVIORAL of IV_118 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity IV_117 is

   port( A : in std_logic;  Y : out std_logic);

end IV_117;

architecture SYN_BEHAVIORAL of IV_117 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity IV_116 is

   port( A : in std_logic;  Y : out std_logic);

end IV_116;

architecture SYN_BEHAVIORAL of IV_116 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity IV_115 is

   port( A : in std_logic;  Y : out std_logic);

end IV_115;

architecture SYN_BEHAVIORAL of IV_115 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity IV_114 is

   port( A : in std_logic;  Y : out std_logic);

end IV_114;

architecture SYN_BEHAVIORAL of IV_114 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity IV_113 is

   port( A : in std_logic;  Y : out std_logic);

end IV_113;

architecture SYN_BEHAVIORAL of IV_113 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity IV_112 is

   port( A : in std_logic;  Y : out std_logic);

end IV_112;

architecture SYN_BEHAVIORAL of IV_112 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity IV_111 is

   port( A : in std_logic;  Y : out std_logic);

end IV_111;

architecture SYN_BEHAVIORAL of IV_111 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity IV_110 is

   port( A : in std_logic;  Y : out std_logic);

end IV_110;

architecture SYN_BEHAVIORAL of IV_110 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity IV_109 is

   port( A : in std_logic;  Y : out std_logic);

end IV_109;

architecture SYN_BEHAVIORAL of IV_109 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity IV_108 is

   port( A : in std_logic;  Y : out std_logic);

end IV_108;

architecture SYN_BEHAVIORAL of IV_108 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity IV_107 is

   port( A : in std_logic;  Y : out std_logic);

end IV_107;

architecture SYN_BEHAVIORAL of IV_107 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity IV_106 is

   port( A : in std_logic;  Y : out std_logic);

end IV_106;

architecture SYN_BEHAVIORAL of IV_106 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity IV_105 is

   port( A : in std_logic;  Y : out std_logic);

end IV_105;

architecture SYN_BEHAVIORAL of IV_105 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity IV_104 is

   port( A : in std_logic;  Y : out std_logic);

end IV_104;

architecture SYN_BEHAVIORAL of IV_104 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity IV_103 is

   port( A : in std_logic;  Y : out std_logic);

end IV_103;

architecture SYN_BEHAVIORAL of IV_103 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity IV_102 is

   port( A : in std_logic;  Y : out std_logic);

end IV_102;

architecture SYN_BEHAVIORAL of IV_102 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity IV_101 is

   port( A : in std_logic;  Y : out std_logic);

end IV_101;

architecture SYN_BEHAVIORAL of IV_101 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity IV_100 is

   port( A : in std_logic;  Y : out std_logic);

end IV_100;

architecture SYN_BEHAVIORAL of IV_100 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity IV_99 is

   port( A : in std_logic;  Y : out std_logic);

end IV_99;

architecture SYN_BEHAVIORAL of IV_99 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity IV_98 is

   port( A : in std_logic;  Y : out std_logic);

end IV_98;

architecture SYN_BEHAVIORAL of IV_98 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity IV_97 is

   port( A : in std_logic;  Y : out std_logic);

end IV_97;

architecture SYN_BEHAVIORAL of IV_97 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity IV_96 is

   port( A : in std_logic;  Y : out std_logic);

end IV_96;

architecture SYN_BEHAVIORAL of IV_96 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity IV_95 is

   port( A : in std_logic;  Y : out std_logic);

end IV_95;

architecture SYN_BEHAVIORAL of IV_95 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity IV_94 is

   port( A : in std_logic;  Y : out std_logic);

end IV_94;

architecture SYN_BEHAVIORAL of IV_94 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity IV_93 is

   port( A : in std_logic;  Y : out std_logic);

end IV_93;

architecture SYN_BEHAVIORAL of IV_93 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity IV_92 is

   port( A : in std_logic;  Y : out std_logic);

end IV_92;

architecture SYN_BEHAVIORAL of IV_92 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity IV_91 is

   port( A : in std_logic;  Y : out std_logic);

end IV_91;

architecture SYN_BEHAVIORAL of IV_91 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity IV_90 is

   port( A : in std_logic;  Y : out std_logic);

end IV_90;

architecture SYN_BEHAVIORAL of IV_90 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity IV_89 is

   port( A : in std_logic;  Y : out std_logic);

end IV_89;

architecture SYN_BEHAVIORAL of IV_89 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity IV_88 is

   port( A : in std_logic;  Y : out std_logic);

end IV_88;

architecture SYN_BEHAVIORAL of IV_88 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity IV_87 is

   port( A : in std_logic;  Y : out std_logic);

end IV_87;

architecture SYN_BEHAVIORAL of IV_87 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity IV_86 is

   port( A : in std_logic;  Y : out std_logic);

end IV_86;

architecture SYN_BEHAVIORAL of IV_86 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity IV_85 is

   port( A : in std_logic;  Y : out std_logic);

end IV_85;

architecture SYN_BEHAVIORAL of IV_85 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity IV_84 is

   port( A : in std_logic;  Y : out std_logic);

end IV_84;

architecture SYN_BEHAVIORAL of IV_84 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity IV_83 is

   port( A : in std_logic;  Y : out std_logic);

end IV_83;

architecture SYN_BEHAVIORAL of IV_83 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity IV_82 is

   port( A : in std_logic;  Y : out std_logic);

end IV_82;

architecture SYN_BEHAVIORAL of IV_82 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity IV_81 is

   port( A : in std_logic;  Y : out std_logic);

end IV_81;

architecture SYN_BEHAVIORAL of IV_81 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity IV_80 is

   port( A : in std_logic;  Y : out std_logic);

end IV_80;

architecture SYN_BEHAVIORAL of IV_80 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity IV_79 is

   port( A : in std_logic;  Y : out std_logic);

end IV_79;

architecture SYN_BEHAVIORAL of IV_79 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity IV_78 is

   port( A : in std_logic;  Y : out std_logic);

end IV_78;

architecture SYN_BEHAVIORAL of IV_78 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity IV_77 is

   port( A : in std_logic;  Y : out std_logic);

end IV_77;

architecture SYN_BEHAVIORAL of IV_77 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity IV_76 is

   port( A : in std_logic;  Y : out std_logic);

end IV_76;

architecture SYN_BEHAVIORAL of IV_76 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity IV_75 is

   port( A : in std_logic;  Y : out std_logic);

end IV_75;

architecture SYN_BEHAVIORAL of IV_75 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity IV_74 is

   port( A : in std_logic;  Y : out std_logic);

end IV_74;

architecture SYN_BEHAVIORAL of IV_74 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity IV_73 is

   port( A : in std_logic;  Y : out std_logic);

end IV_73;

architecture SYN_BEHAVIORAL of IV_73 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity IV_72 is

   port( A : in std_logic;  Y : out std_logic);

end IV_72;

architecture SYN_BEHAVIORAL of IV_72 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity IV_71 is

   port( A : in std_logic;  Y : out std_logic);

end IV_71;

architecture SYN_BEHAVIORAL of IV_71 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity IV_70 is

   port( A : in std_logic;  Y : out std_logic);

end IV_70;

architecture SYN_BEHAVIORAL of IV_70 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity IV_69 is

   port( A : in std_logic;  Y : out std_logic);

end IV_69;

architecture SYN_BEHAVIORAL of IV_69 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity IV_68 is

   port( A : in std_logic;  Y : out std_logic);

end IV_68;

architecture SYN_BEHAVIORAL of IV_68 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity IV_67 is

   port( A : in std_logic;  Y : out std_logic);

end IV_67;

architecture SYN_BEHAVIORAL of IV_67 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity IV_66 is

   port( A : in std_logic;  Y : out std_logic);

end IV_66;

architecture SYN_BEHAVIORAL of IV_66 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity IV_65 is

   port( A : in std_logic;  Y : out std_logic);

end IV_65;

architecture SYN_BEHAVIORAL of IV_65 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1996 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1996;

architecture SYN_BEHAVIORAL of FA_1996 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n3, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U1 : INV_X1 port map( A => n2, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n3, B2 => Ci, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_2006 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2006;

architecture SYN_BEHAVIORAL of FA_2006 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n3, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U1 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n3, B2 => Ci, ZN => n2);
   U2 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_2010 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2010;

architecture SYN_BEHAVIORAL of FA_2010 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U1 : XOR2_X1 port map( A => Ci, B => n3, Z => S);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n3, B2 => Ci, ZN => n2);
   U3 : INV_X1 port map( A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_2047 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2047;

architecture SYN_BEHAVIORAL of FA_2047 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net63890, net83667, n3, n2, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => B, ZN => n7);
   U2 : AOI22_X1 port map( A1 => B, A2 => n6, B1 => Ci, B2 => n3, ZN => n2);
   U3 : INV_X1 port map( A => n2, ZN => Co);
   U4 : CLKBUF_X1 port map( A => A, Z => n6);
   U5 : CLKBUF_X1 port map( A => Ci, Z => net63890);
   U6 : XNOR2_X1 port map( A => A, B => n7, ZN => n3);
   U7 : CLKBUF_X1 port map( A => n3, Z => net83667);
   U8 : XOR2_X1 port map( A => net63890, B => net83667, Z => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity FA_1024 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1024;

architecture SYN_BEHAVIORAL of FA_1024 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net83665, net83535, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => B, ZN => net83535);
   U2 : AOI21_X1 port map( B1 => A, B2 => Ci, A => B, ZN => n6);
   U3 : NOR2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U4 : CLKBUF_X1 port map( A => A, Z => net83665);
   U5 : NOR2_X1 port map( A1 => net83665, A2 => Ci, ZN => n5);
   U6 : XNOR2_X1 port map( A => net83665, B => net83535, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity RCA_NbitRca64_31 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_NbitRca64_31;

architecture SYN_STRUCTURAL of RCA_NbitRca64_31 is

   component FA_1921
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1922
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1923
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1924
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1925
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1926
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1927
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1928
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1929
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1930
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1931
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1932
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1933
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1934
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1935
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1936
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1937
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1938
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1939
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1940
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1941
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1942
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1943
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1944
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1945
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1946
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1947
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1948
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1949
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1950
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1951
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1952
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1953
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1954
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1955
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1956
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1957
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1958
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1959
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1960
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1961
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1962
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1963
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1964
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1965
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1966
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1967
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1968
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1969
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1970
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1971
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1972
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1973
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1974
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1975
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1976
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1977
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1978
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1979
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1980
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1981
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1982
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1983
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1984
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_63_port, CTMP_62_port, CTMP_61_port, CTMP_60_port, CTMP_59_port,
      CTMP_58_port, CTMP_57_port, CTMP_56_port, CTMP_55_port, CTMP_54_port, 
      CTMP_53_port, CTMP_52_port, CTMP_51_port, CTMP_50_port, CTMP_49_port, 
      CTMP_48_port, CTMP_47_port, CTMP_46_port, CTMP_45_port, CTMP_44_port, 
      CTMP_43_port, CTMP_42_port, CTMP_41_port, CTMP_40_port, CTMP_39_port, 
      CTMP_38_port, CTMP_37_port, CTMP_36_port, CTMP_35_port, CTMP_34_port, 
      CTMP_33_port, CTMP_32_port, CTMP_31_port, CTMP_30_port, CTMP_29_port, 
      CTMP_28_port, CTMP_27_port, CTMP_26_port, CTMP_25_port, CTMP_24_port, 
      CTMP_23_port, CTMP_22_port, CTMP_21_port, CTMP_20_port, CTMP_19_port, 
      CTMP_18_port, CTMP_17_port, CTMP_16_port, CTMP_15_port, CTMP_14_port, 
      CTMP_13_port, CTMP_12_port, CTMP_11_port, CTMP_10_port, CTMP_9_port, 
      CTMP_8_port, CTMP_7_port, CTMP_6_port, CTMP_5_port, CTMP_4_port, 
      CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_1984 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_1983 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1)
                           , Co => CTMP_2_port);
   FAI_3 : FA_1982 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2)
                           , Co => CTMP_3_port);
   FAI_4 : FA_1981 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3)
                           , Co => CTMP_4_port);
   FAI_5 : FA_1980 port map( A => A(4), B => B(4), Ci => CTMP_4_port, S => S(4)
                           , Co => CTMP_5_port);
   FAI_6 : FA_1979 port map( A => A(5), B => B(5), Ci => CTMP_5_port, S => S(5)
                           , Co => CTMP_6_port);
   FAI_7 : FA_1978 port map( A => A(6), B => B(6), Ci => CTMP_6_port, S => S(6)
                           , Co => CTMP_7_port);
   FAI_8 : FA_1977 port map( A => A(7), B => B(7), Ci => CTMP_7_port, S => S(7)
                           , Co => CTMP_8_port);
   FAI_9 : FA_1976 port map( A => A(8), B => B(8), Ci => CTMP_8_port, S => S(8)
                           , Co => CTMP_9_port);
   FAI_10 : FA_1975 port map( A => A(9), B => B(9), Ci => CTMP_9_port, S => 
                           S(9), Co => CTMP_10_port);
   FAI_11 : FA_1974 port map( A => A(10), B => B(10), Ci => CTMP_10_port, S => 
                           S(10), Co => CTMP_11_port);
   FAI_12 : FA_1973 port map( A => A(11), B => B(11), Ci => CTMP_11_port, S => 
                           S(11), Co => CTMP_12_port);
   FAI_13 : FA_1972 port map( A => A(12), B => B(12), Ci => CTMP_12_port, S => 
                           S(12), Co => CTMP_13_port);
   FAI_14 : FA_1971 port map( A => A(13), B => B(13), Ci => CTMP_13_port, S => 
                           S(13), Co => CTMP_14_port);
   FAI_15 : FA_1970 port map( A => A(14), B => B(14), Ci => CTMP_14_port, S => 
                           S(14), Co => CTMP_15_port);
   FAI_16 : FA_1969 port map( A => A(15), B => B(15), Ci => CTMP_15_port, S => 
                           S(15), Co => CTMP_16_port);
   FAI_17 : FA_1968 port map( A => A(16), B => B(16), Ci => CTMP_16_port, S => 
                           S(16), Co => CTMP_17_port);
   FAI_18 : FA_1967 port map( A => A(17), B => B(17), Ci => CTMP_17_port, S => 
                           S(17), Co => CTMP_18_port);
   FAI_19 : FA_1966 port map( A => A(18), B => B(18), Ci => CTMP_18_port, S => 
                           S(18), Co => CTMP_19_port);
   FAI_20 : FA_1965 port map( A => A(19), B => B(19), Ci => CTMP_19_port, S => 
                           S(19), Co => CTMP_20_port);
   FAI_21 : FA_1964 port map( A => A(20), B => B(20), Ci => CTMP_20_port, S => 
                           S(20), Co => CTMP_21_port);
   FAI_22 : FA_1963 port map( A => A(21), B => B(21), Ci => CTMP_21_port, S => 
                           S(21), Co => CTMP_22_port);
   FAI_23 : FA_1962 port map( A => A(22), B => B(22), Ci => CTMP_22_port, S => 
                           S(22), Co => CTMP_23_port);
   FAI_24 : FA_1961 port map( A => A(23), B => B(23), Ci => CTMP_23_port, S => 
                           S(23), Co => CTMP_24_port);
   FAI_25 : FA_1960 port map( A => A(24), B => B(24), Ci => CTMP_24_port, S => 
                           S(24), Co => CTMP_25_port);
   FAI_26 : FA_1959 port map( A => A(25), B => B(25), Ci => CTMP_25_port, S => 
                           S(25), Co => CTMP_26_port);
   FAI_27 : FA_1958 port map( A => A(26), B => B(26), Ci => CTMP_26_port, S => 
                           S(26), Co => CTMP_27_port);
   FAI_28 : FA_1957 port map( A => A(27), B => B(27), Ci => CTMP_27_port, S => 
                           S(27), Co => CTMP_28_port);
   FAI_29 : FA_1956 port map( A => A(28), B => B(28), Ci => CTMP_28_port, S => 
                           S(28), Co => CTMP_29_port);
   FAI_30 : FA_1955 port map( A => A(29), B => B(29), Ci => CTMP_29_port, S => 
                           S(29), Co => CTMP_30_port);
   FAI_31 : FA_1954 port map( A => A(30), B => B(30), Ci => CTMP_30_port, S => 
                           S(30), Co => CTMP_31_port);
   FAI_32 : FA_1953 port map( A => A(31), B => B(31), Ci => CTMP_31_port, S => 
                           S(31), Co => CTMP_32_port);
   FAI_33 : FA_1952 port map( A => A(32), B => B(32), Ci => CTMP_32_port, S => 
                           S(32), Co => CTMP_33_port);
   FAI_34 : FA_1951 port map( A => A(33), B => B(33), Ci => CTMP_33_port, S => 
                           S(33), Co => CTMP_34_port);
   FAI_35 : FA_1950 port map( A => A(34), B => B(34), Ci => CTMP_34_port, S => 
                           S(34), Co => CTMP_35_port);
   FAI_36 : FA_1949 port map( A => A(35), B => B(35), Ci => CTMP_35_port, S => 
                           S(35), Co => CTMP_36_port);
   FAI_37 : FA_1948 port map( A => A(36), B => B(36), Ci => CTMP_36_port, S => 
                           S(36), Co => CTMP_37_port);
   FAI_38 : FA_1947 port map( A => A(37), B => B(37), Ci => CTMP_37_port, S => 
                           S(37), Co => CTMP_38_port);
   FAI_39 : FA_1946 port map( A => A(38), B => B(38), Ci => CTMP_38_port, S => 
                           S(38), Co => CTMP_39_port);
   FAI_40 : FA_1945 port map( A => A(39), B => B(39), Ci => CTMP_39_port, S => 
                           S(39), Co => CTMP_40_port);
   FAI_41 : FA_1944 port map( A => A(40), B => B(40), Ci => CTMP_40_port, S => 
                           S(40), Co => CTMP_41_port);
   FAI_42 : FA_1943 port map( A => A(41), B => B(41), Ci => CTMP_41_port, S => 
                           S(41), Co => CTMP_42_port);
   FAI_43 : FA_1942 port map( A => A(42), B => B(42), Ci => CTMP_42_port, S => 
                           S(42), Co => CTMP_43_port);
   FAI_44 : FA_1941 port map( A => A(43), B => B(43), Ci => CTMP_43_port, S => 
                           S(43), Co => CTMP_44_port);
   FAI_45 : FA_1940 port map( A => A(44), B => B(44), Ci => CTMP_44_port, S => 
                           S(44), Co => CTMP_45_port);
   FAI_46 : FA_1939 port map( A => A(45), B => B(45), Ci => CTMP_45_port, S => 
                           S(45), Co => CTMP_46_port);
   FAI_47 : FA_1938 port map( A => A(46), B => B(46), Ci => CTMP_46_port, S => 
                           S(46), Co => CTMP_47_port);
   FAI_48 : FA_1937 port map( A => A(47), B => B(47), Ci => CTMP_47_port, S => 
                           S(47), Co => CTMP_48_port);
   FAI_49 : FA_1936 port map( A => A(48), B => B(48), Ci => CTMP_48_port, S => 
                           S(48), Co => CTMP_49_port);
   FAI_50 : FA_1935 port map( A => A(49), B => B(49), Ci => CTMP_49_port, S => 
                           S(49), Co => CTMP_50_port);
   FAI_51 : FA_1934 port map( A => A(50), B => B(50), Ci => CTMP_50_port, S => 
                           S(50), Co => CTMP_51_port);
   FAI_52 : FA_1933 port map( A => A(51), B => B(51), Ci => CTMP_51_port, S => 
                           S(51), Co => CTMP_52_port);
   FAI_53 : FA_1932 port map( A => A(52), B => B(52), Ci => CTMP_52_port, S => 
                           S(52), Co => CTMP_53_port);
   FAI_54 : FA_1931 port map( A => A(53), B => B(53), Ci => CTMP_53_port, S => 
                           S(53), Co => CTMP_54_port);
   FAI_55 : FA_1930 port map( A => A(54), B => B(54), Ci => CTMP_54_port, S => 
                           S(54), Co => CTMP_55_port);
   FAI_56 : FA_1929 port map( A => A(55), B => B(55), Ci => CTMP_55_port, S => 
                           S(55), Co => CTMP_56_port);
   FAI_57 : FA_1928 port map( A => A(56), B => B(56), Ci => CTMP_56_port, S => 
                           S(56), Co => CTMP_57_port);
   FAI_58 : FA_1927 port map( A => A(57), B => B(57), Ci => CTMP_57_port, S => 
                           S(57), Co => CTMP_58_port);
   FAI_59 : FA_1926 port map( A => A(58), B => B(58), Ci => CTMP_58_port, S => 
                           S(58), Co => CTMP_59_port);
   FAI_60 : FA_1925 port map( A => A(59), B => B(59), Ci => CTMP_59_port, S => 
                           S(59), Co => CTMP_60_port);
   FAI_61 : FA_1924 port map( A => A(60), B => B(60), Ci => CTMP_60_port, S => 
                           S(60), Co => CTMP_61_port);
   FAI_62 : FA_1923 port map( A => A(61), B => B(61), Ci => CTMP_61_port, S => 
                           S(61), Co => CTMP_62_port);
   FAI_63 : FA_1922 port map( A => A(62), B => B(62), Ci => CTMP_62_port, S => 
                           S(62), Co => CTMP_63_port);
   FAI_64 : FA_1921 port map( A => A(63), B => B(63), Ci => CTMP_63_port, S => 
                           S(63), Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity MUX51_MuxNbit64_16 is

   port( zeroSignal, A_signal, A_neg, A_shifted, A_neg_shifted : in 
         std_logic_vector (63 downto 0);  Sel : in std_logic_vector (2 downto 
         0);  Y : out std_logic_vector (63 downto 0));

end MUX51_MuxNbit64_16;

architecture SYN_BEHAVIORAL_2 of MUX51_MuxNbit64_16 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X4
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X8
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n10, n11, n12, n13, n14, n16, n17, n18, n19, n20, n21, n22, 
      n23, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39
      , n40, n41, n42, n43, n44, n45, n46, n48, n49, n50, n51, n52, n53, n54, 
      n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70
      , n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, 
      n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99
      , n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
      n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, 
      n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, 
      net58758, net58748, net58746, net58744, net58776, net58772, net58770, 
      net58790, net58788, net58786, net58784, net58782, net58780, net58810, 
      net58808, net58806, net58804, net61182, net61181, net61179, net61178, 
      net58814, net58794, n68, net83887, net84205, net84185, net84181, net84175
      , net84173, net84171, net84116, net84113, n15, net84210, net84203, 
      net84177, net84169, net84167, net84222, net84186, net83612, net58792, 
      net58742, n9, n5, n25, n24, n141, n142, n143, n144, n145, n146, n147, 
      n148, n149, n150, n151, n152, n153 : std_logic;

begin
   
   U1 : NOR2_X1 port map( A1 => n143, A2 => n152, ZN => n91);
   U2 : NAND2_X1 port map( A1 => n153, A2 => net84185, ZN => n152);
   U3 : NAND2_X1 port map( A1 => n5, A2 => A_shifted(2), ZN => net84185);
   U4 : INV_X1 port map( A => A_shifted(3), ZN => net84171);
   U5 : INV_X1 port map( A => zeroSignal(4), ZN => net84175);
   U6 : INV_X1 port map( A => n147, ZN => n9);
   U7 : NAND2_X1 port map( A1 => n150, A2 => net84169, ZN => net84177);
   U8 : BUF_X2 port map( A => net58810, Z => net58806);
   U9 : BUF_X1 port map( A => net58814, Z => net58810);
   U10 : AND2_X1 port map( A1 => n145, A2 => net84116, ZN => n141);
   U11 : AND3_X1 port map( A1 => n146, A2 => net84113, A3 => Sel(1), ZN => n142
                           );
   U12 : INV_X1 port map( A => net84167, ZN => n5);
   U13 : BUF_X1 port map( A => net58742, Z => net61179);
   U14 : AND2_X1 port map( A1 => zeroSignal(2), A2 => net58746, ZN => n143);
   U15 : AND2_X1 port map( A1 => zeroSignal(3), A2 => net58748, ZN => n144);
   U16 : OR2_X1 port map( A1 => net84175, A2 => net84177, ZN => n145);
   U17 : NAND2_X1 port map( A1 => net84205, A2 => A_neg_shifted(2), ZN => n153)
                           ;
   U18 : NAND2_X1 port map( A1 => n24, A2 => n25, ZN => Y(5));
   U19 : AOI222_X1 port map( A1 => A_shifted(5), A2 => net58742, B1 => 
                           zeroSignal(5), B2 => net58758, C1 => 
                           A_neg_shifted(5), C2 => net58776, ZN => n25);
   U20 : INV_X2 port map( A => net84169, ZN => net58776);
   U21 : INV_X2 port map( A => net84177, ZN => net58758);
   U22 : BUF_X1 port map( A => n5, Z => net58742);
   U23 : CLKBUF_X1 port map( A => net58742, Z => net61178);
   U24 : NAND2_X1 port map( A1 => A_shifted(4), A2 => n5, ZN => net84116);
   U25 : AOI22_X1 port map( A1 => A_neg(5), A2 => net58788, B1 => A_signal(5), 
                           B2 => net83612, ZN => n24);
   U26 : CLKBUF_X1 port map( A => net58814, Z => net83612);
   U27 : BUF_X1 port map( A => n9, Z => net58814);
   U28 : AOI22_X1 port map( A1 => A_neg(3), A2 => net58784, B1 => A_signal(3), 
                           B2 => n9, ZN => n68);
   U29 : AOI22_X1 port map( A1 => A_neg(2), A2 => net58782, B1 => A_signal(2), 
                           B2 => n9, ZN => n90);
   U30 : NAND2_X1 port map( A1 => net84186, A2 => net84113, ZN => n147);
   U31 : INV_X1 port map( A => Sel(2), ZN => net84113);
   U32 : NOR2_X1 port map( A1 => n146, A2 => net84222, ZN => net84186);
   U33 : BUF_X1 port map( A => Sel(1), Z => net84222);
   U34 : INV_X1 port map( A => Sel(0), ZN => n146);
   U35 : INV_X1 port map( A => n146, ZN => net84203);
   U36 : BUF_X1 port map( A => net58792, Z => net58788);
   U37 : CLKBUF_X1 port map( A => n142, Z => net58792);
   U38 : BUF_X1 port map( A => net58792, Z => net58786);
   U39 : BUF_X1 port map( A => net58792, Z => net58790);
   U40 : BUF_X1 port map( A => n142, Z => net58794);
   U41 : NAND2_X1 port map( A1 => n149, A2 => net84210, ZN => net84169);
   U42 : OAI22_X1 port map( A1 => net84169, A2 => net84173, B1 => net84167, B2 
                           => net84171, ZN => net84181);
   U43 : INV_X1 port map( A => net84169, ZN => net84205);
   U44 : INV_X1 port map( A => net84113, ZN => net84210);
   U45 : NOR2_X1 port map( A1 => Sel(1), A2 => Sel(0), ZN => n149);
   U46 : OAI21_X1 port map( B1 => net84222, B2 => net84203, A => net84113, ZN 
                           => n150);
   U47 : NAND2_X1 port map( A1 => n148, A2 => net84113, ZN => net84167);
   U48 : AND2_X1 port map( A1 => Sel(0), A2 => Sel(1), ZN => n148);
   U49 : AOI222_X1 port map( A1 => A_shifted(6), A2 => net61179, B1 => 
                           zeroSignal(6), B2 => net58758, C1 => 
                           A_neg_shifted(6), C2 => net58776, ZN => n15);
   U50 : NAND2_X1 port map( A1 => n14, A2 => n15, ZN => Y(6));
   U51 : NAND3_X1 port map( A1 => n46, A2 => n151, A3 => n141, ZN => Y(4));
   U52 : NAND2_X1 port map( A1 => A_neg_shifted(4), A2 => net58776, ZN => n151)
                           ;
   U53 : INV_X1 port map( A => A_neg_shifted(3), ZN => net84173);
   U54 : CLKBUF_X1 port map( A => net58782, Z => net83887);
   U55 : NOR2_X1 port map( A1 => net84181, A2 => n144, ZN => n69);
   U56 : BUF_X2 port map( A => net58794, Z => net58782);
   U57 : CLKBUF_X1 port map( A => net58810, Z => net58808);
   U58 : CLKBUF_X1 port map( A => net58810, Z => net58804);
   U59 : BUF_X1 port map( A => net61178, Z => net61181);
   U60 : BUF_X8 port map( A => net61179, Z => net61182);
   U61 : BUF_X4 port map( A => net58776, Z => net58770);
   U62 : NAND2_X1 port map( A1 => n68, A2 => n69, ZN => Y(3));
   U63 : BUF_X2 port map( A => net58794, Z => net58784);
   U64 : CLKBUF_X1 port map( A => net58794, Z => net58780);
   U65 : CLKBUF_X1 port map( A => net58776, Z => net58772);
   U66 : BUF_X1 port map( A => net58758, Z => net58748);
   U67 : BUF_X1 port map( A => net58758, Z => net58746);
   U68 : BUF_X1 port map( A => net58758, Z => net58744);
   U69 : NAND2_X1 port map( A1 => n132, A2 => n133, ZN => Y(10));
   U70 : AOI22_X1 port map( A1 => A_neg(10), A2 => net58780, B1 => A_signal(10)
                           , B2 => net58808, ZN => n132);
   U71 : NAND2_X1 port map( A1 => n128, A2 => n129, ZN => Y(12));
   U72 : AOI222_X1 port map( A1 => A_shifted(12), A2 => net61182, B1 => 
                           zeroSignal(12), B2 => net58744, C1 => 
                           A_neg_shifted(12), C2 => net58776, ZN => n129);
   U73 : AOI222_X1 port map( A1 => A_shifted(11), A2 => net61182, B1 => 
                           zeroSignal(11), B2 => net58744, C1 => 
                           A_neg_shifted(11), C2 => net58770, ZN => n131);
   U74 : AOI222_X1 port map( A1 => A_shifted(13), A2 => net61182, B1 => 
                           zeroSignal(13), B2 => net58744, C1 => 
                           A_neg_shifted(13), C2 => net58772, ZN => n127);
   U75 : NAND2_X1 port map( A1 => n34, A2 => n35, ZN => Y(55));
   U76 : AOI222_X1 port map( A1 => A_shifted(55), A2 => net61182, B1 => 
                           zeroSignal(55), B2 => net58758, C1 => 
                           A_neg_shifted(55), C2 => net58770, ZN => n35);
   U77 : AOI22_X1 port map( A1 => A_neg(55), A2 => net58788, B1 => A_signal(55)
                           , B2 => net58804, ZN => n34);
   U78 : NAND2_X1 port map( A1 => n124, A2 => n125, ZN => Y(14));
   U79 : AOI222_X1 port map( A1 => A_shifted(14), A2 => net61182, B1 => 
                           zeroSignal(14), B2 => net58744, C1 => 
                           A_neg_shifted(14), C2 => net58770, ZN => n125);
   U80 : AOI222_X1 port map( A1 => A_shifted(37), A2 => net61182, B1 => 
                           zeroSignal(37), B2 => net58748, C1 => 
                           A_neg_shifted(37), C2 => net58770, ZN => n75);
   U81 : NAND2_X1 port map( A1 => n118, A2 => n119, ZN => Y(17));
   U82 : AOI222_X1 port map( A1 => A_shifted(17), A2 => net61182, B1 => 
                           zeroSignal(17), B2 => net58744, C1 => 
                           A_neg_shifted(17), C2 => net58770, ZN => n119);
   U83 : AOI222_X1 port map( A1 => A_shifted(16), A2 => net61182, B1 => 
                           zeroSignal(16), B2 => net58744, C1 => 
                           A_neg_shifted(16), C2 => net58770, ZN => n121);
   U84 : NAND2_X1 port map( A1 => n114, A2 => n115, ZN => Y(19));
   U85 : NAND2_X1 port map( A1 => n36, A2 => n37, ZN => Y(54));
   U86 : AOI22_X1 port map( A1 => A_neg(54), A2 => net58788, B1 => A_signal(54)
                           , B2 => net58808, ZN => n36);
   U87 : NAND2_X1 port map( A1 => n28, A2 => n29, ZN => Y(58));
   U88 : AOI222_X1 port map( A1 => A_shifted(58), A2 => net61182, B1 => 
                           zeroSignal(58), B2 => net58758, C1 => 
                           A_neg_shifted(58), C2 => net58776, ZN => n29);
   U89 : AOI22_X1 port map( A1 => A_neg(58), A2 => net58788, B1 => A_signal(58)
                           , B2 => net58806, ZN => n28);
   U90 : NAND2_X1 port map( A1 => n116, A2 => n117, ZN => Y(18));
   U91 : AOI222_X1 port map( A1 => A_shifted(18), A2 => net61182, B1 => 
                           zeroSignal(18), B2 => net58744, C1 => 
                           A_neg_shifted(18), C2 => net58770, ZN => n117);
   U92 : NAND2_X1 port map( A1 => n30, A2 => n31, ZN => Y(57));
   U93 : AOI222_X1 port map( A1 => A_shifted(57), A2 => net61182, B1 => 
                           zeroSignal(57), B2 => net58758, C1 => 
                           A_neg_shifted(57), C2 => net58772, ZN => n31);
   U94 : AOI22_X1 port map( A1 => A_neg(57), A2 => net58788, B1 => A_signal(57)
                           , B2 => net58808, ZN => n30);
   U95 : NAND2_X1 port map( A1 => n32, A2 => n33, ZN => Y(56));
   U96 : AOI222_X1 port map( A1 => A_shifted(56), A2 => net61181, B1 => 
                           zeroSignal(56), B2 => net58758, C1 => 
                           A_neg_shifted(56), C2 => net58776, ZN => n33);
   U97 : AOI22_X1 port map( A1 => A_neg(56), A2 => net58788, B1 => A_signal(56)
                           , B2 => net58806, ZN => n32);
   U98 : NAND2_X1 port map( A1 => n22, A2 => n23, ZN => Y(60));
   U99 : AOI222_X1 port map( A1 => A_shifted(60), A2 => net61182, B1 => 
                           zeroSignal(60), B2 => net58758, C1 => 
                           A_neg_shifted(60), C2 => net58772, ZN => n23);
   U100 : AOI22_X1 port map( A1 => A_neg(60), A2 => net58788, B1 => 
                           A_signal(60), B2 => net58804, ZN => n22);
   U101 : NAND2_X1 port map( A1 => n26, A2 => n27, ZN => Y(59));
   U102 : AOI222_X1 port map( A1 => A_shifted(59), A2 => net61181, B1 => 
                           zeroSignal(59), B2 => net58758, C1 => 
                           A_neg_shifted(59), C2 => net58770, ZN => n27);
   U103 : AOI22_X1 port map( A1 => A_neg(59), A2 => net58788, B1 => 
                           A_signal(59), B2 => net58804, ZN => n26);
   U104 : NAND2_X1 port map( A1 => n58, A2 => n59, ZN => Y(44));
   U105 : AOI222_X1 port map( A1 => A_shifted(44), A2 => net61182, B1 => 
                           zeroSignal(44), B2 => net58758, C1 => 
                           A_neg_shifted(44), C2 => net58772, ZN => n59);
   U106 : NAND2_X1 port map( A1 => n106, A2 => n107, ZN => Y(22));
   U107 : AOI222_X1 port map( A1 => A_shifted(22), A2 => net61182, B1 => 
                           zeroSignal(22), B2 => net58746, C1 => 
                           A_neg_shifted(22), C2 => net58770, ZN => n107);
   U108 : AOI22_X1 port map( A1 => A_neg(22), A2 => net58782, B1 => 
                           A_signal(22), B2 => net58806, ZN => n106);
   U109 : AOI222_X1 port map( A1 => A_shifted(20), A2 => net61182, B1 => 
                           zeroSignal(20), B2 => net58746, C1 => 
                           A_neg_shifted(20), C2 => net58770, ZN => n111);
   U110 : AOI222_X1 port map( A1 => A_shifted(21), A2 => net61182, B1 => 
                           zeroSignal(21), B2 => net58746, C1 => 
                           A_neg_shifted(21), C2 => net58770, ZN => n109);
   U111 : NAND2_X1 port map( A1 => n18, A2 => n19, ZN => Y(62));
   U112 : AOI222_X1 port map( A1 => A_shifted(62), A2 => net61181, B1 => 
                           zeroSignal(62), B2 => net58758, C1 => 
                           A_neg_shifted(62), C2 => net58772, ZN => n19);
   U113 : AOI22_X1 port map( A1 => A_neg(62), A2 => net58788, B1 => 
                           A_signal(62), B2 => net58806, ZN => n18);
   U114 : NAND2_X1 port map( A1 => n16, A2 => n17, ZN => Y(63));
   U115 : AOI222_X1 port map( A1 => A_shifted(63), A2 => net61181, B1 => 
                           zeroSignal(63), B2 => net58758, C1 => 
                           A_neg_shifted(63), C2 => net58776, ZN => n17);
   U116 : AOI22_X1 port map( A1 => A_neg(63), A2 => net58788, B1 => 
                           A_signal(63), B2 => net58804, ZN => n16);
   U117 : NAND2_X1 port map( A1 => n38, A2 => n39, ZN => Y(53));
   U118 : AOI222_X1 port map( A1 => A_shifted(53), A2 => net61182, B1 => 
                           zeroSignal(53), B2 => net58758, C1 => 
                           A_neg_shifted(53), C2 => net58772, ZN => n39);
   U119 : NAND2_X1 port map( A1 => n20, A2 => n21, ZN => Y(61));
   U120 : AOI222_X1 port map( A1 => A_shifted(61), A2 => net61181, B1 => 
                           zeroSignal(61), B2 => net58758, C1 => 
                           A_neg_shifted(61), C2 => net58770, ZN => n21);
   U121 : AOI22_X1 port map( A1 => A_neg(61), A2 => net58788, B1 => 
                           A_signal(61), B2 => net58808, ZN => n20);
   U122 : AOI222_X1 port map( A1 => A_shifted(41), A2 => net61182, B1 => 
                           zeroSignal(41), B2 => net58748, C1 => 
                           A_neg_shifted(41), C2 => net58770, ZN => n65);
   U123 : AOI222_X1 port map( A1 => A_shifted(23), A2 => net61182, B1 => 
                           zeroSignal(23), B2 => net58746, C1 => 
                           A_neg_shifted(23), C2 => net58770, ZN => n105);
   U124 : NAND2_X1 port map( A1 => n96, A2 => n97, ZN => Y(27));
   U125 : AOI222_X1 port map( A1 => A_shifted(27), A2 => net61182, B1 => 
                           zeroSignal(27), B2 => net58746, C1 => 
                           A_neg_shifted(27), C2 => net58770, ZN => n97);
   U126 : NAND2_X1 port map( A1 => n102, A2 => n103, ZN => Y(24));
   U127 : AOI222_X1 port map( A1 => A_shifted(24), A2 => net61182, B1 => 
                           zeroSignal(24), B2 => net58746, C1 => 
                           A_neg_shifted(24), C2 => net58770, ZN => n103);
   U128 : NAND2_X1 port map( A1 => n98, A2 => n99, ZN => Y(26));
   U129 : AOI222_X1 port map( A1 => A_shifted(26), A2 => net61182, B1 => 
                           zeroSignal(26), B2 => net58746, C1 => 
                           A_neg_shifted(26), C2 => net58770, ZN => n99);
   U130 : AOI22_X1 port map( A1 => A_neg(26), A2 => net58782, B1 => 
                           A_signal(26), B2 => net58806, ZN => n98);
   U131 : NAND2_X1 port map( A1 => n60, A2 => n61, ZN => Y(43));
   U132 : AOI222_X1 port map( A1 => A_shifted(43), A2 => net61182, B1 => 
                           zeroSignal(43), B2 => net58758, C1 => 
                           A_neg_shifted(43), C2 => net58772, ZN => n61);
   U133 : NAND2_X1 port map( A1 => n54, A2 => n55, ZN => Y(46));
   U134 : AOI222_X1 port map( A1 => A_shifted(46), A2 => net61181, B1 => 
                           zeroSignal(46), B2 => net58758, C1 => 
                           A_neg_shifted(46), C2 => net58770, ZN => n55);
   U135 : NAND2_X1 port map( A1 => n56, A2 => n57, ZN => Y(45));
   U136 : NAND2_X1 port map( A1 => n52, A2 => n53, ZN => Y(47));
   U137 : NAND2_X1 port map( A1 => n82, A2 => n83, ZN => Y(33));
   U138 : AOI222_X1 port map( A1 => A_shifted(33), A2 => net61182, B1 => 
                           zeroSignal(33), B2 => net58748, C1 => 
                           A_neg_shifted(33), C2 => net58770, ZN => n83);
   U139 : NAND2_X1 port map( A1 => n50, A2 => n51, ZN => Y(48));
   U140 : NAND2_X1 port map( A1 => n62, A2 => n63, ZN => Y(42));
   U141 : AOI22_X1 port map( A1 => A_neg(42), A2 => net58786, B1 => 
                           A_signal(42), B2 => net58804, ZN => n62);
   U142 : AOI222_X1 port map( A1 => A_shifted(42), A2 => net61182, B1 => 
                           zeroSignal(42), B2 => net58758, C1 => 
                           A_neg_shifted(42), C2 => net58772, ZN => n63);
   U143 : NAND2_X1 port map( A1 => n44, A2 => n45, ZN => Y(50));
   U144 : AOI222_X1 port map( A1 => A_shifted(50), A2 => net61182, B1 => 
                           zeroSignal(50), B2 => net58758, C1 => 
                           A_neg_shifted(50), C2 => net58776, ZN => n45);
   U145 : NAND2_X1 port map( A1 => n94, A2 => n95, ZN => Y(28));
   U146 : AOI222_X1 port map( A1 => A_shifted(28), A2 => net61182, B1 => 
                           zeroSignal(28), B2 => net58746, C1 => 
                           A_neg_shifted(28), C2 => net58772, ZN => n95);
   U147 : NAND2_X1 port map( A1 => n92, A2 => n93, ZN => Y(29));
   U148 : AOI222_X1 port map( A1 => A_shifted(29), A2 => net61182, B1 => 
                           zeroSignal(29), B2 => net58746, C1 => 
                           A_neg_shifted(29), C2 => net58770, ZN => n93);
   U149 : AOI22_X1 port map( A1 => A_neg(29), A2 => net83887, B1 => 
                           A_signal(29), B2 => net58804, ZN => n92);
   U150 : NAND2_X1 port map( A1 => n88, A2 => n89, ZN => Y(30));
   U151 : AOI222_X1 port map( A1 => A_shifted(30), A2 => net61182, B1 => 
                           zeroSignal(30), B2 => net58746, C1 => 
                           A_neg_shifted(30), C2 => net58772, ZN => n89);
   U152 : AOI22_X1 port map( A1 => A_neg(30), A2 => net83887, B1 => 
                           A_signal(30), B2 => net58806, ZN => n88);
   U153 : NAND2_X1 port map( A1 => n40, A2 => n41, ZN => Y(52));
   U154 : AOI222_X1 port map( A1 => A_shifted(52), A2 => net61181, B1 => 
                           zeroSignal(52), B2 => net58758, C1 => 
                           A_neg_shifted(52), C2 => net58776, ZN => n41);
   U155 : AOI22_X1 port map( A1 => A_neg(52), A2 => net58786, B1 => 
                           A_signal(52), B2 => net58804, ZN => n40);
   U156 : NAND2_X1 port map( A1 => n42, A2 => n43, ZN => Y(51));
   U157 : AOI22_X1 port map( A1 => A_neg(51), A2 => net58786, B1 => 
                           A_signal(51), B2 => net58806, ZN => n42);
   U158 : AOI222_X1 port map( A1 => A_shifted(31), A2 => net61182, B1 => 
                           zeroSignal(31), B2 => net58748, C1 => 
                           A_neg_shifted(31), C2 => net58770, ZN => n87);
   U159 : NAND2_X1 port map( A1 => n48, A2 => n49, ZN => Y(49));
   U160 : AOI22_X1 port map( A1 => A_neg(49), A2 => net58786, B1 => 
                           A_signal(49), B2 => net58806, ZN => n48);
   U161 : AOI222_X1 port map( A1 => A_shifted(32), A2 => net61182, B1 => 
                           zeroSignal(32), B2 => net58748, C1 => 
                           A_neg_shifted(32), C2 => net58772, ZN => n85);
   U162 : AOI22_X1 port map( A1 => A_neg(32), A2 => net58784, B1 => 
                           A_signal(32), B2 => net58806, ZN => n84);
   U163 : AOI222_X1 port map( A1 => A_shifted(34), A2 => net61182, B1 => 
                           zeroSignal(34), B2 => net58748, C1 => 
                           A_neg_shifted(34), C2 => net58772, ZN => n81);
   U164 : AOI22_X1 port map( A1 => A_neg(34), A2 => net58784, B1 => 
                           A_signal(34), B2 => net58806, ZN => n80);
   U165 : NAND2_X1 port map( A1 => n78, A2 => n79, ZN => Y(35));
   U166 : AOI222_X1 port map( A1 => A_shifted(35), A2 => net61182, B1 => 
                           zeroSignal(35), B2 => net58748, C1 => 
                           A_neg_shifted(35), C2 => net58770, ZN => n79);
   U167 : AOI22_X1 port map( A1 => A_neg(35), A2 => net58784, B1 => 
                           A_signal(35), B2 => net58804, ZN => n78);
   U168 : NAND2_X1 port map( A1 => n72, A2 => n73, ZN => Y(38));
   U169 : AOI22_X1 port map( A1 => A_neg(38), A2 => net58784, B1 => 
                           A_signal(38), B2 => net58806, ZN => n72);
   U170 : NAND2_X1 port map( A1 => n70, A2 => n71, ZN => Y(39));
   U171 : AOI222_X1 port map( A1 => A_shifted(39), A2 => net61182, B1 => 
                           zeroSignal(39), B2 => net58748, C1 => 
                           A_neg_shifted(39), C2 => net58770, ZN => n71);
   U172 : AOI22_X1 port map( A1 => A_neg(39), A2 => net58784, B1 => 
                           A_signal(39), B2 => net58804, ZN => n70);
   U173 : NAND2_X1 port map( A1 => n76, A2 => n77, ZN => Y(36));
   U174 : AOI222_X1 port map( A1 => A_shifted(36), A2 => net61182, B1 => 
                           zeroSignal(36), B2 => net58748, C1 => 
                           A_neg_shifted(36), C2 => net58772, ZN => n77);
   U175 : AOI22_X1 port map( A1 => A_neg(36), A2 => net58784, B1 => 
                           A_signal(36), B2 => net58806, ZN => n76);
   U176 : NAND2_X1 port map( A1 => n66, A2 => n67, ZN => Y(40));
   U177 : AOI222_X1 port map( A1 => A_shifted(40), A2 => net61182, B1 => 
                           zeroSignal(40), B2 => net58748, C1 => 
                           A_neg_shifted(40), C2 => net58772, ZN => n67);
   U178 : AOI22_X1 port map( A1 => A_neg(40), A2 => net58784, B1 => 
                           A_signal(40), B2 => net58806, ZN => n66);
   U179 : AOI22_X1 port map( A1 => A_neg(1), A2 => net58780, B1 => A_signal(1),
                           B2 => net58808, ZN => n112);
   U180 : AOI222_X1 port map( A1 => A_shifted(0), A2 => net61181, B1 => 
                           zeroSignal(0), B2 => net58744, C1 => 
                           A_neg_shifted(0), C2 => net58770, ZN => n135);
   U181 : AOI222_X1 port map( A1 => A_shifted(9), A2 => net61181, B1 => 
                           zeroSignal(9), B2 => net58758, C1 => 
                           A_neg_shifted(9), C2 => net58770, ZN => n4);
   U182 : AOI222_X1 port map( A1 => A_shifted(51), A2 => net61182, B1 => 
                           zeroSignal(51), B2 => net58758, C1 => 
                           A_neg_shifted(51), C2 => net58770, ZN => n43);
   U183 : AOI22_X1 port map( A1 => A_neg(50), A2 => net58786, B1 => 
                           A_signal(50), B2 => net58804, ZN => n44);
   U184 : AOI222_X1 port map( A1 => A_shifted(54), A2 => net61181, B1 => 
                           zeroSignal(54), B2 => net58758, C1 => 
                           A_neg_shifted(54), C2 => net58776, ZN => n37);
   U185 : AOI22_X1 port map( A1 => A_neg(53), A2 => net58788, B1 => 
                           A_signal(53), B2 => net58806, ZN => n38);
   U186 : AOI222_X1 port map( A1 => A_shifted(49), A2 => net61181, B1 => 
                           zeroSignal(49), B2 => net58758, C1 => 
                           A_neg_shifted(49), C2 => net58772, ZN => n49);
   U187 : AOI22_X1 port map( A1 => A_neg(48), A2 => net58786, B1 => 
                           A_signal(48), B2 => net58804, ZN => n50);
   U188 : AOI222_X1 port map( A1 => A_shifted(47), A2 => net61182, B1 => 
                           zeroSignal(47), B2 => net58758, C1 => 
                           A_neg_shifted(47), C2 => net58772, ZN => n53);
   U189 : AOI22_X1 port map( A1 => A_neg(46), A2 => net58786, B1 => 
                           A_signal(46), B2 => net58804, ZN => n54);
   U190 : AOI222_X1 port map( A1 => A_shifted(48), A2 => net61182, B1 => 
                           zeroSignal(48), B2 => net58758, C1 => 
                           A_neg_shifted(48), C2 => net58770, ZN => n51);
   U191 : AOI22_X1 port map( A1 => A_neg(47), A2 => net58786, B1 => 
                           A_signal(47), B2 => net58806, ZN => n52);
   U192 : AOI222_X1 port map( A1 => A_shifted(45), A2 => net61182, B1 => 
                           zeroSignal(45), B2 => net58758, C1 => 
                           A_neg_shifted(45), C2 => net58770, ZN => n57);
   U193 : AOI22_X1 port map( A1 => A_neg(44), A2 => net58786, B1 => 
                           A_signal(44), B2 => net58804, ZN => n58);
   U194 : NAND2_X1 port map( A1 => n112, A2 => n113, ZN => Y(1));
   U195 : NAND2_X1 port map( A1 => n134, A2 => n135, ZN => Y(0));
   U196 : AOI22_X1 port map( A1 => A_neg(0), A2 => net58780, B1 => A_signal(0),
                           B2 => net58806, ZN => n134);
   U197 : AOI222_X1 port map( A1 => A_shifted(1), A2 => net61182, B1 => 
                           zeroSignal(1), B2 => net58744, C1 => 
                           A_neg_shifted(1), C2 => net58776, ZN => n113);
   U198 : NAND2_X1 port map( A1 => n3, A2 => n4, ZN => Y(9));
   U199 : AOI222_X1 port map( A1 => A_shifted(10), A2 => net61182, B1 => 
                           zeroSignal(10), B2 => net58744, C1 => 
                           A_neg_shifted(10), C2 => net58770, ZN => n133);
   U200 : NAND2_X1 port map( A1 => n86, A2 => n87, ZN => Y(31));
   U201 : AOI22_X1 port map( A1 => A_neg(31), A2 => net58784, B1 => 
                           A_signal(31), B2 => net58804, ZN => n86);
   U202 : NAND2_X1 port map( A1 => n10, A2 => n11, ZN => Y(8));
   U203 : AOI22_X1 port map( A1 => A_neg(45), A2 => net58786, B1 => 
                           A_signal(45), B2 => net58806, ZN => n56);
   U204 : AOI22_X1 port map( A1 => A_neg(43), A2 => net58786, B1 => 
                           A_signal(43), B2 => net58806, ZN => n60);
   U205 : NAND2_X1 port map( A1 => n80, A2 => n81, ZN => Y(34));
   U206 : AOI222_X1 port map( A1 => A_shifted(8), A2 => net61179, B1 => 
                           zeroSignal(8), B2 => net58758, C1 => 
                           A_neg_shifted(8), C2 => net58770, ZN => n11);
   U207 : NAND2_X1 port map( A1 => n12, A2 => n13, ZN => Y(7));
   U208 : AOI22_X1 port map( A1 => A_neg(33), A2 => net58784, B1 => 
                           A_signal(33), B2 => net58804, ZN => n82);
   U209 : NAND2_X1 port map( A1 => n84, A2 => n85, ZN => Y(32));
   U210 : AOI222_X1 port map( A1 => A_shifted(7), A2 => net61178, B1 => 
                           zeroSignal(7), B2 => net58758, C1 => 
                           A_neg_shifted(7), C2 => net58770, ZN => n13);
   U211 : AOI222_X1 port map( A1 => A_shifted(38), A2 => net61182, B1 => 
                           zeroSignal(38), B2 => net58748, C1 => 
                           A_neg_shifted(38), C2 => net58772, ZN => n73);
   U212 : NAND2_X1 port map( A1 => n64, A2 => n65, ZN => Y(41));
   U213 : AOI22_X1 port map( A1 => A_neg(41), A2 => net58784, B1 => 
                           A_signal(41), B2 => net58804, ZN => n64);
   U214 : AOI22_X1 port map( A1 => A_neg(28), A2 => net58782, B1 => 
                           A_signal(28), B2 => net58804, ZN => n94);
   U215 : NAND2_X1 port map( A1 => n74, A2 => n75, ZN => Y(37));
   U216 : AOI22_X1 port map( A1 => A_neg(27), A2 => net58782, B1 => 
                           A_signal(27), B2 => net58806, ZN => n96);
   U217 : AOI22_X1 port map( A1 => A_neg(25), A2 => net58782, B1 => 
                           A_signal(25), B2 => net58806, ZN => n100);
   U218 : NAND2_X1 port map( A1 => n100, A2 => n101, ZN => Y(25));
   U219 : AOI222_X1 port map( A1 => A_shifted(25), A2 => net61182, B1 => 
                           zeroSignal(25), B2 => net58746, C1 => 
                           A_neg_shifted(25), C2 => net58770, ZN => n101);
   U220 : AOI22_X1 port map( A1 => A_neg(24), A2 => net58782, B1 => 
                           A_signal(24), B2 => net58806, ZN => n102);
   U221 : AOI22_X1 port map( A1 => A_neg(23), A2 => net58782, B1 => 
                           A_signal(23), B2 => net58806, ZN => n104);
   U222 : NAND2_X1 port map( A1 => n104, A2 => n105, ZN => Y(23));
   U223 : AOI22_X1 port map( A1 => A_neg(20), A2 => net58782, B1 => 
                           A_signal(20), B2 => net58806, ZN => n110);
   U224 : NAND2_X1 port map( A1 => n110, A2 => n111, ZN => Y(20));
   U225 : AOI22_X1 port map( A1 => A_neg(21), A2 => net58782, B1 => 
                           A_signal(21), B2 => net58806, ZN => n108);
   U226 : NAND2_X1 port map( A1 => n108, A2 => n109, ZN => Y(21));
   U227 : AOI22_X1 port map( A1 => A_neg(19), A2 => net58780, B1 => 
                           A_signal(19), B2 => net58806, ZN => n114);
   U228 : AOI222_X1 port map( A1 => A_shifted(19), A2 => net61182, B1 => 
                           zeroSignal(19), B2 => net58744, C1 => 
                           A_neg_shifted(19), C2 => net58770, ZN => n115);
   U229 : AOI22_X1 port map( A1 => A_neg(18), A2 => net58780, B1 => 
                           A_signal(18), B2 => net58806, ZN => n116);
   U230 : NAND2_X1 port map( A1 => n90, A2 => n91, ZN => Y(2));
   U231 : AOI22_X1 port map( A1 => A_neg(15), A2 => net58780, B1 => 
                           A_signal(15), B2 => net58806, ZN => n122);
   U232 : NAND2_X1 port map( A1 => n122, A2 => n123, ZN => Y(15));
   U233 : AOI22_X1 port map( A1 => A_neg(17), A2 => net58780, B1 => 
                           A_signal(17), B2 => net58806, ZN => n118);
   U234 : AOI22_X1 port map( A1 => A_neg(16), A2 => net58780, B1 => 
                           A_signal(16), B2 => net58806, ZN => n120);
   U235 : NAND2_X1 port map( A1 => n120, A2 => n121, ZN => Y(16));
   U236 : AOI222_X1 port map( A1 => A_shifted(15), A2 => net61182, B1 => 
                           zeroSignal(15), B2 => net58744, C1 => 
                           A_neg_shifted(15), C2 => net58770, ZN => n123);
   U237 : AOI22_X1 port map( A1 => A_neg(14), A2 => net58780, B1 => 
                           A_signal(14), B2 => net58806, ZN => n124);
   U238 : AOI22_X1 port map( A1 => A_neg(11), A2 => net58780, B1 => 
                           A_signal(11), B2 => net58808, ZN => n130);
   U239 : NAND2_X1 port map( A1 => n130, A2 => n131, ZN => Y(11));
   U240 : AOI22_X1 port map( A1 => A_neg(13), A2 => net58780, B1 => 
                           A_signal(13), B2 => net58804, ZN => n126);
   U241 : AOI22_X1 port map( A1 => A_neg(12), A2 => net58780, B1 => 
                           A_signal(12), B2 => net58808, ZN => n128);
   U242 : AOI22_X1 port map( A1 => A_neg(9), A2 => net58790, B1 => A_signal(9),
                           B2 => net58808, ZN => n3);
   U243 : NAND2_X1 port map( A1 => n126, A2 => n127, ZN => Y(13));
   U244 : AOI22_X1 port map( A1 => A_neg(7), A2 => net58790, B1 => A_signal(7),
                           B2 => net58810, ZN => n12);
   U245 : AOI22_X1 port map( A1 => A_neg(8), A2 => net58790, B1 => A_signal(8),
                           B2 => net58810, ZN => n10);
   U246 : AOI22_X1 port map( A1 => A_neg(6), A2 => net58790, B1 => A_signal(6),
                           B2 => net58810, ZN => n14);
   U247 : AOI22_X1 port map( A1 => A_neg(4), A2 => net58786, B1 => A_signal(4),
                           B2 => net58814, ZN => n46);
   U248 : AOI22_X1 port map( A1 => A_neg(37), A2 => net58784, B1 => 
                           A_signal(37), B2 => net58804, ZN => n74);

end SYN_BEHAVIORAL_2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity encoder_16 is

   port( pieceofB : in std_logic_vector (2 downto 0);  sel : out 
         std_logic_vector (2 downto 0));

end encoder_16;

architecture SYN_behavioral of encoder_16 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => pieceofB(1), A2 => pieceofB(0), ZN => n2);
   U4 : NOR3_X1 port map( A1 => n1, A2 => pieceofB(1), A3 => pieceofB(0), ZN =>
                           sel(2));
   U5 : OAI21_X1 port map( B1 => pieceofB(1), B2 => pieceofB(0), A => n2, ZN =>
                           n4);
   U6 : INV_X1 port map( A => pieceofB(2), ZN => n1);
   U7 : AOI21_X1 port map( B1 => n4, B2 => n2, A => pieceofB(2), ZN => sel(0));
   U8 : OAI21_X1 port map( B1 => pieceofB(1), B2 => pieceofB(0), A => n2, ZN =>
                           n3);
   U9 : OAI22_X1 port map( A1 => n1, A2 => n3, B1 => pieceofB(2), B2 => n2, ZN 
                           => sel(1));

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity leftshifter_NbitShifter64_63 is

   port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
         std_logic_vector (63 downto 0));

end leftshifter_NbitShifter64_63;

architecture SYN_behavioral of leftshifter_NbitShifter64_63 is

signal X_Logic0_port : std_logic;

begin
   shift_out <= ( shift_in(62), shift_in(61), shift_in(60), shift_in(59), 
      shift_in(58), shift_in(57), shift_in(56), shift_in(55), shift_in(54), 
      shift_in(53), shift_in(52), shift_in(51), shift_in(50), shift_in(49), 
      shift_in(48), shift_in(47), shift_in(46), shift_in(45), shift_in(44), 
      shift_in(43), shift_in(42), shift_in(41), shift_in(40), shift_in(39), 
      shift_in(38), shift_in(37), shift_in(36), shift_in(35), shift_in(34), 
      shift_in(33), shift_in(32), shift_in(31), shift_in(30), shift_in(29), 
      shift_in(28), shift_in(27), shift_in(26), shift_in(25), shift_in(24), 
      shift_in(23), shift_in(22), shift_in(21), shift_in(20), shift_in(19), 
      shift_in(18), shift_in(17), shift_in(16), shift_in(15), shift_in(14), 
      shift_in(13), shift_in(12), shift_in(11), shift_in(10), shift_in(9), 
      shift_in(8), shift_in(7), shift_in(6), shift_in(5), shift_in(4), 
      shift_in(3), shift_in(2), shift_in(1), shift_in(0), X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity RCA_NbitRca64_16 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_NbitRca64_16;

architecture SYN_STRUCTURAL of RCA_NbitRca64_16 is

   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component FA_1985
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1986
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1987
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1988
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1989
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1990
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1991
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1992
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1993
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1994
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1995
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1996
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1997
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1998
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1999
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_2000
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_2001
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_2002
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_2003
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_2004
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_2005
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_2006
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_2007
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_2008
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_2009
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_2010
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_2011
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_2012
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_2013
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_2014
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_2015
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_2016
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_2017
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_2018
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_2019
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_2020
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_2021
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_2022
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_2023
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_2024
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_2025
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_2026
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_2027
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_2028
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_2029
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_2030
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_2031
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_2032
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_2033
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_2034
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_2035
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_2036
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_2037
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_2038
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_2039
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_2040
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_2041
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_2042
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_2043
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_2044
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_2045
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_2046
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_2047
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1024
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n2, CTMP_63_port, CTMP_62_port, CTMP_61_port, CTMP_60_port, 
      CTMP_59_port, CTMP_58_port, CTMP_57_port, CTMP_56_port, CTMP_55_port, 
      CTMP_54_port, CTMP_53_port, CTMP_52_port, CTMP_51_port, CTMP_50_port, 
      CTMP_49_port, CTMP_48_port, CTMP_47_port, CTMP_46_port, CTMP_45_port, 
      CTMP_44_port, CTMP_43_port, CTMP_42_port, CTMP_41_port, CTMP_40_port, 
      CTMP_39_port, CTMP_38_port, CTMP_37_port, CTMP_36_port, CTMP_35_port, 
      CTMP_34_port, CTMP_33_port, CTMP_32_port, CTMP_31_port, CTMP_30_port, 
      CTMP_29_port, CTMP_28_port, CTMP_27_port, CTMP_26_port, CTMP_25_port, 
      CTMP_24_port, CTMP_23_port, CTMP_22_port, CTMP_21_port, CTMP_20_port, 
      CTMP_19_port, CTMP_18_port, CTMP_17_port, CTMP_16_port, CTMP_15_port, 
      CTMP_14_port, CTMP_13_port, CTMP_12_port, CTMP_11_port, CTMP_10_port, 
      CTMP_9_port, CTMP_8_port, CTMP_7_port, CTMP_6_port, CTMP_5_port, 
      CTMP_4_port, CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_1024 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_2047 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1)
                           , Co => CTMP_2_port);
   FAI_3 : FA_2046 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2)
                           , Co => CTMP_3_port);
   FAI_4 : FA_2045 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3)
                           , Co => CTMP_4_port);
   FAI_5 : FA_2044 port map( A => A(4), B => B(4), Ci => CTMP_4_port, S => S(4)
                           , Co => CTMP_5_port);
   FAI_6 : FA_2043 port map( A => A(5), B => B(5), Ci => CTMP_5_port, S => S(5)
                           , Co => CTMP_6_port);
   FAI_7 : FA_2042 port map( A => A(6), B => B(6), Ci => CTMP_6_port, S => S(6)
                           , Co => CTMP_7_port);
   FAI_8 : FA_2041 port map( A => A(7), B => B(7), Ci => CTMP_7_port, S => S(7)
                           , Co => CTMP_8_port);
   FAI_9 : FA_2040 port map( A => A(8), B => B(8), Ci => CTMP_8_port, S => S(8)
                           , Co => CTMP_9_port);
   FAI_10 : FA_2039 port map( A => A(9), B => B(9), Ci => CTMP_9_port, S => 
                           S(9), Co => CTMP_10_port);
   FAI_11 : FA_2038 port map( A => A(10), B => B(10), Ci => CTMP_10_port, S => 
                           S(10), Co => CTMP_11_port);
   FAI_12 : FA_2037 port map( A => A(11), B => B(11), Ci => CTMP_11_port, S => 
                           S(11), Co => CTMP_12_port);
   FAI_13 : FA_2036 port map( A => A(12), B => B(12), Ci => CTMP_12_port, S => 
                           S(12), Co => CTMP_13_port);
   FAI_14 : FA_2035 port map( A => A(13), B => B(13), Ci => CTMP_13_port, S => 
                           S(13), Co => CTMP_14_port);
   FAI_15 : FA_2034 port map( A => A(14), B => B(14), Ci => CTMP_14_port, S => 
                           S(14), Co => CTMP_15_port);
   FAI_16 : FA_2033 port map( A => A(15), B => B(15), Ci => CTMP_15_port, S => 
                           S(15), Co => CTMP_16_port);
   FAI_17 : FA_2032 port map( A => A(16), B => B(16), Ci => CTMP_16_port, S => 
                           S(16), Co => CTMP_17_port);
   FAI_18 : FA_2031 port map( A => A(17), B => B(17), Ci => CTMP_17_port, S => 
                           S(17), Co => CTMP_18_port);
   FAI_19 : FA_2030 port map( A => A(18), B => B(18), Ci => CTMP_18_port, S => 
                           S(18), Co => CTMP_19_port);
   FAI_20 : FA_2029 port map( A => A(19), B => B(19), Ci => CTMP_19_port, S => 
                           S(19), Co => CTMP_20_port);
   FAI_21 : FA_2028 port map( A => A(20), B => B(20), Ci => CTMP_20_port, S => 
                           S(20), Co => CTMP_21_port);
   FAI_22 : FA_2027 port map( A => A(21), B => B(21), Ci => CTMP_21_port, S => 
                           S(21), Co => CTMP_22_port);
   FAI_23 : FA_2026 port map( A => A(22), B => B(22), Ci => CTMP_22_port, S => 
                           S(22), Co => CTMP_23_port);
   FAI_24 : FA_2025 port map( A => A(23), B => B(23), Ci => CTMP_23_port, S => 
                           S(23), Co => CTMP_24_port);
   FAI_25 : FA_2024 port map( A => A(24), B => B(24), Ci => CTMP_24_port, S => 
                           S(24), Co => CTMP_25_port);
   FAI_26 : FA_2023 port map( A => A(25), B => B(25), Ci => CTMP_25_port, S => 
                           S(25), Co => CTMP_26_port);
   FAI_27 : FA_2022 port map( A => A(26), B => B(26), Ci => CTMP_26_port, S => 
                           S(26), Co => CTMP_27_port);
   FAI_28 : FA_2021 port map( A => A(27), B => B(27), Ci => CTMP_27_port, S => 
                           S(27), Co => CTMP_28_port);
   FAI_29 : FA_2020 port map( A => A(28), B => B(28), Ci => CTMP_28_port, S => 
                           S(28), Co => CTMP_29_port);
   FAI_30 : FA_2019 port map( A => A(29), B => B(29), Ci => CTMP_29_port, S => 
                           S(29), Co => CTMP_30_port);
   FAI_31 : FA_2018 port map( A => A(30), B => B(30), Ci => CTMP_30_port, S => 
                           S(30), Co => CTMP_31_port);
   FAI_32 : FA_2017 port map( A => A(31), B => B(31), Ci => CTMP_31_port, S => 
                           S(31), Co => CTMP_32_port);
   FAI_33 : FA_2016 port map( A => A(32), B => B(32), Ci => CTMP_32_port, S => 
                           S(32), Co => CTMP_33_port);
   FAI_34 : FA_2015 port map( A => A(33), B => B(33), Ci => CTMP_33_port, S => 
                           S(33), Co => CTMP_34_port);
   FAI_35 : FA_2014 port map( A => A(34), B => B(34), Ci => CTMP_34_port, S => 
                           S(34), Co => CTMP_35_port);
   FAI_36 : FA_2013 port map( A => A(35), B => B(35), Ci => CTMP_35_port, S => 
                           S(35), Co => CTMP_36_port);
   FAI_37 : FA_2012 port map( A => A(36), B => B(36), Ci => CTMP_36_port, S => 
                           S(36), Co => CTMP_37_port);
   FAI_38 : FA_2011 port map( A => A(37), B => B(37), Ci => CTMP_37_port, S => 
                           S(37), Co => CTMP_38_port);
   FAI_39 : FA_2010 port map( A => A(38), B => B(38), Ci => CTMP_38_port, S => 
                           S(38), Co => CTMP_39_port);
   FAI_40 : FA_2009 port map( A => A(39), B => B(39), Ci => CTMP_39_port, S => 
                           S(39), Co => CTMP_40_port);
   FAI_41 : FA_2008 port map( A => A(40), B => B(40), Ci => CTMP_40_port, S => 
                           S(40), Co => CTMP_41_port);
   FAI_42 : FA_2007 port map( A => A(41), B => B(41), Ci => CTMP_41_port, S => 
                           S(41), Co => CTMP_42_port);
   FAI_43 : FA_2006 port map( A => A(42), B => B(42), Ci => CTMP_42_port, S => 
                           n2, Co => CTMP_43_port);
   FAI_44 : FA_2005 port map( A => A(43), B => B(43), Ci => CTMP_43_port, S => 
                           S(43), Co => CTMP_44_port);
   FAI_45 : FA_2004 port map( A => A(44), B => B(44), Ci => CTMP_44_port, S => 
                           S(44), Co => CTMP_45_port);
   FAI_46 : FA_2003 port map( A => A(45), B => B(45), Ci => CTMP_45_port, S => 
                           S(45), Co => CTMP_46_port);
   FAI_47 : FA_2002 port map( A => A(46), B => B(46), Ci => CTMP_46_port, S => 
                           S(46), Co => CTMP_47_port);
   FAI_48 : FA_2001 port map( A => A(47), B => B(47), Ci => CTMP_47_port, S => 
                           S(47), Co => CTMP_48_port);
   FAI_49 : FA_2000 port map( A => A(48), B => B(48), Ci => CTMP_48_port, S => 
                           S(48), Co => CTMP_49_port);
   FAI_50 : FA_1999 port map( A => A(49), B => B(49), Ci => CTMP_49_port, S => 
                           S(49), Co => CTMP_50_port);
   FAI_51 : FA_1998 port map( A => A(50), B => B(50), Ci => CTMP_50_port, S => 
                           S(50), Co => CTMP_51_port);
   FAI_52 : FA_1997 port map( A => A(51), B => B(51), Ci => CTMP_51_port, S => 
                           S(51), Co => CTMP_52_port);
   FAI_53 : FA_1996 port map( A => A(52), B => B(52), Ci => CTMP_52_port, S => 
                           S(52), Co => CTMP_53_port);
   FAI_54 : FA_1995 port map( A => A(53), B => B(53), Ci => CTMP_53_port, S => 
                           S(53), Co => CTMP_54_port);
   FAI_55 : FA_1994 port map( A => A(54), B => B(54), Ci => CTMP_54_port, S => 
                           S(54), Co => CTMP_55_port);
   FAI_56 : FA_1993 port map( A => A(55), B => B(55), Ci => CTMP_55_port, S => 
                           S(55), Co => CTMP_56_port);
   FAI_57 : FA_1992 port map( A => A(56), B => B(56), Ci => CTMP_56_port, S => 
                           S(56), Co => CTMP_57_port);
   FAI_58 : FA_1991 port map( A => A(57), B => B(57), Ci => CTMP_57_port, S => 
                           S(57), Co => CTMP_58_port);
   FAI_59 : FA_1990 port map( A => A(58), B => B(58), Ci => CTMP_58_port, S => 
                           S(58), Co => CTMP_59_port);
   FAI_60 : FA_1989 port map( A => A(59), B => B(59), Ci => CTMP_59_port, S => 
                           S(59), Co => CTMP_60_port);
   FAI_61 : FA_1988 port map( A => A(60), B => B(60), Ci => CTMP_60_port, S => 
                           S(60), Co => CTMP_61_port);
   FAI_62 : FA_1987 port map( A => A(61), B => B(61), Ci => CTMP_61_port, S => 
                           S(61), Co => CTMP_62_port);
   FAI_63 : FA_1986 port map( A => A(62), B => B(62), Ci => CTMP_62_port, S => 
                           S(62), Co => CTMP_63_port);
   FAI_64 : FA_1985 port map( A => A(63), B => B(63), Ci => CTMP_63_port, S => 
                           S(63), Co => Co);
   U1 : BUF_X2 port map( A => n2, Z => S(42));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity IV_64 is

   port( A : in std_logic;  Y : out std_logic);

end IV_64;

architecture SYN_BEHAVIORAL of IV_64 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_1.all;

entity BOOTHMUL_1 is

   port( A, B : in std_logic_vector (31 downto 0);  P : out std_logic_vector 
         (63 downto 0));

end BOOTHMUL_1;

architecture SYN_STRUCTURAL of BOOTHMUL_1 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component RCA_NbitRca64_17
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NbitRca64_18
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NbitRca64_19
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NbitRca64_20
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NbitRca64_21
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NbitRca64_22
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NbitRca64_23
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NbitRca64_24
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NbitRca64_25
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NbitRca64_26
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NbitRca64_27
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NbitRca64_28
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NbitRca64_29
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NbitRca64_30
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NbitRca64_31
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component MUX51_MuxNbit64_17
      port( zeroSignal, A_signal, A_neg, A_shifted, A_neg_shifted : in 
            std_logic_vector (63 downto 0);  Sel : in std_logic_vector (2 
            downto 0);  Y : out std_logic_vector (63 downto 0));
   end component;
   
   component encoder_17
      port( pieceofB : in std_logic_vector (2 downto 0);  sel : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component MUX51_MuxNbit64_18
      port( zeroSignal, A_signal, A_neg, A_shifted, A_neg_shifted : in 
            std_logic_vector (63 downto 0);  Sel : in std_logic_vector (2 
            downto 0);  Y : out std_logic_vector (63 downto 0));
   end component;
   
   component encoder_18
      port( pieceofB : in std_logic_vector (2 downto 0);  sel : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component MUX51_MuxNbit64_19
      port( zeroSignal, A_signal, A_neg, A_shifted, A_neg_shifted : in 
            std_logic_vector (63 downto 0);  Sel : in std_logic_vector (2 
            downto 0);  Y : out std_logic_vector (63 downto 0));
   end component;
   
   component encoder_19
      port( pieceofB : in std_logic_vector (2 downto 0);  sel : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component MUX51_MuxNbit64_20
      port( zeroSignal, A_signal, A_neg, A_shifted, A_neg_shifted : in 
            std_logic_vector (63 downto 0);  Sel : in std_logic_vector (2 
            downto 0);  Y : out std_logic_vector (63 downto 0));
   end component;
   
   component encoder_20
      port( pieceofB : in std_logic_vector (2 downto 0);  sel : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component MUX51_MuxNbit64_21
      port( zeroSignal, A_signal, A_neg, A_shifted, A_neg_shifted : in 
            std_logic_vector (63 downto 0);  Sel : in std_logic_vector (2 
            downto 0);  Y : out std_logic_vector (63 downto 0));
   end component;
   
   component encoder_21
      port( pieceofB : in std_logic_vector (2 downto 0);  sel : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component MUX51_MuxNbit64_22
      port( zeroSignal, A_signal, A_neg, A_shifted, A_neg_shifted : in 
            std_logic_vector (63 downto 0);  Sel : in std_logic_vector (2 
            downto 0);  Y : out std_logic_vector (63 downto 0));
   end component;
   
   component encoder_22
      port( pieceofB : in std_logic_vector (2 downto 0);  sel : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component MUX51_MuxNbit64_23
      port( zeroSignal, A_signal, A_neg, A_shifted, A_neg_shifted : in 
            std_logic_vector (63 downto 0);  Sel : in std_logic_vector (2 
            downto 0);  Y : out std_logic_vector (63 downto 0));
   end component;
   
   component encoder_23
      port( pieceofB : in std_logic_vector (2 downto 0);  sel : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component MUX51_MuxNbit64_24
      port( zeroSignal, A_signal, A_neg, A_shifted, A_neg_shifted : in 
            std_logic_vector (63 downto 0);  Sel : in std_logic_vector (2 
            downto 0);  Y : out std_logic_vector (63 downto 0));
   end component;
   
   component encoder_24
      port( pieceofB : in std_logic_vector (2 downto 0);  sel : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component MUX51_MuxNbit64_25
      port( zeroSignal, A_signal, A_neg, A_shifted, A_neg_shifted : in 
            std_logic_vector (63 downto 0);  Sel : in std_logic_vector (2 
            downto 0);  Y : out std_logic_vector (63 downto 0));
   end component;
   
   component encoder_25
      port( pieceofB : in std_logic_vector (2 downto 0);  sel : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component MUX51_MuxNbit64_26
      port( zeroSignal, A_signal, A_neg, A_shifted, A_neg_shifted : in 
            std_logic_vector (63 downto 0);  Sel : in std_logic_vector (2 
            downto 0);  Y : out std_logic_vector (63 downto 0));
   end component;
   
   component encoder_26
      port( pieceofB : in std_logic_vector (2 downto 0);  sel : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component MUX51_MuxNbit64_27
      port( zeroSignal, A_signal, A_neg, A_shifted, A_neg_shifted : in 
            std_logic_vector (63 downto 0);  Sel : in std_logic_vector (2 
            downto 0);  Y : out std_logic_vector (63 downto 0));
   end component;
   
   component encoder_27
      port( pieceofB : in std_logic_vector (2 downto 0);  sel : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component MUX51_MuxNbit64_28
      port( zeroSignal, A_signal, A_neg, A_shifted, A_neg_shifted : in 
            std_logic_vector (63 downto 0);  Sel : in std_logic_vector (2 
            downto 0);  Y : out std_logic_vector (63 downto 0));
   end component;
   
   component encoder_28
      port( pieceofB : in std_logic_vector (2 downto 0);  sel : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component MUX51_MuxNbit64_29
      port( zeroSignal, A_signal, A_neg, A_shifted, A_neg_shifted : in 
            std_logic_vector (63 downto 0);  Sel : in std_logic_vector (2 
            downto 0);  Y : out std_logic_vector (63 downto 0));
   end component;
   
   component encoder_29
      port( pieceofB : in std_logic_vector (2 downto 0);  sel : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component MUX51_MuxNbit64_30
      port( zeroSignal, A_signal, A_neg, A_shifted, A_neg_shifted : in 
            std_logic_vector (63 downto 0);  Sel : in std_logic_vector (2 
            downto 0);  Y : out std_logic_vector (63 downto 0));
   end component;
   
   component encoder_30
      port( pieceofB : in std_logic_vector (2 downto 0);  sel : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component MUX51_MuxNbit64_31
      port( zeroSignal, A_signal, A_neg, A_shifted, A_neg_shifted : in 
            std_logic_vector (63 downto 0);  Sel : in std_logic_vector (2 
            downto 0);  Y : out std_logic_vector (63 downto 0));
   end component;
   
   component encoder_31
      port( pieceofB : in std_logic_vector (2 downto 0);  sel : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component MUX51_MuxNbit64_16
      port( zeroSignal, A_signal, A_neg, A_shifted, A_neg_shifted : in 
            std_logic_vector (63 downto 0);  Sel : in std_logic_vector (2 
            downto 0);  Y : out std_logic_vector (63 downto 0));
   end component;
   
   component encoder_16
      port( pieceofB : in std_logic_vector (2 downto 0);  sel : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_64
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_65
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_66
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_67
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_68
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_69
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_70
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_71
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_72
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_73
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_74
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_75
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_76
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_77
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_78
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_79
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_80
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_81
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_82
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_83
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_84
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_85
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_86
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_87
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_88
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_89
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_90
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_91
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_92
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_93
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_94
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_95
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_96
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_97
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_98
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_99
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_100
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_101
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_102
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_103
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_104
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_105
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_106
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_107
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_108
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_109
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_110
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_111
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_112
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_113
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_114
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_115
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_116
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_117
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_118
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_119
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_120
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_121
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_122
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_123
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_124
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_125
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component leftshifter_NbitShifter64_63
      port( shift_in : in std_logic_vector (63 downto 0);  shift_out : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component RCA_NbitRca64_16
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component IV_65
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_66
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_67
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_68
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_69
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_70
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_71
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_72
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_73
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_74
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_75
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_76
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_77
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_78
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_79
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_80
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_81
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_82
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_83
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_84
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_85
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_86
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_87
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_88
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_89
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_90
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_91
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_92
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_93
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_94
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_95
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_96
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_97
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_98
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_99
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_100
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_101
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_102
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_103
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_104
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_105
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_106
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_107
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_108
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_109
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_110
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_111
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_112
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_113
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_114
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_115
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_116
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_117
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_118
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_119
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_120
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_121
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_122
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_123
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_124
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_125
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_126
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_127
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_64
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, A_complement_63_port, 
      A_complement_62_port, A_complement_61_port, A_complement_60_port, 
      A_complement_59_port, A_complement_58_port, A_complement_57_port, 
      A_complement_56_port, A_complement_55_port, A_complement_54_port, 
      A_complement_53_port, A_complement_52_port, A_complement_51_port, 
      A_complement_50_port, A_complement_49_port, A_complement_48_port, 
      A_complement_47_port, A_complement_46_port, A_complement_45_port, 
      A_complement_44_port, A_complement_43_port, A_complement_42_port, 
      A_complement_41_port, A_complement_40_port, A_complement_39_port, 
      A_complement_38_port, A_complement_37_port, A_complement_36_port, 
      A_complement_35_port, A_complement_34_port, A_complement_33_port, 
      A_complement_32_port, A_complement_31_port, A_complement_30_port, 
      A_complement_29_port, A_complement_28_port, A_complement_27_port, 
      A_complement_26_port, A_complement_25_port, A_complement_24_port, 
      A_complement_23_port, A_complement_22_port, A_complement_21_port, 
      A_complement_20_port, A_complement_19_port, A_complement_18_port, 
      A_complement_17_port, A_complement_16_port, A_complement_15_port, 
      A_complement_14_port, A_complement_13_port, A_complement_12_port, 
      A_complement_11_port, A_complement_10_port, A_complement_9_port, 
      A_complement_8_port, A_complement_7_port, A_complement_6_port, 
      A_complement_5_port, A_complement_4_port, A_complement_3_port, 
      A_complement_2_port, A_complement_1_port, A_complement_0_port, 
      negative_inputs_0_63_port, negative_inputs_0_62_port, 
      negative_inputs_0_61_port, negative_inputs_0_60_port, 
      negative_inputs_0_59_port, negative_inputs_0_58_port, 
      negative_inputs_0_57_port, negative_inputs_0_56_port, 
      negative_inputs_0_55_port, negative_inputs_0_54_port, 
      negative_inputs_0_53_port, negative_inputs_0_52_port, 
      negative_inputs_0_51_port, negative_inputs_0_50_port, 
      negative_inputs_0_49_port, negative_inputs_0_48_port, 
      negative_inputs_0_47_port, negative_inputs_0_46_port, 
      negative_inputs_0_45_port, negative_inputs_0_44_port, 
      negative_inputs_0_43_port, negative_inputs_0_42_port, 
      negative_inputs_0_41_port, negative_inputs_0_40_port, 
      negative_inputs_0_39_port, negative_inputs_0_38_port, 
      negative_inputs_0_37_port, negative_inputs_0_36_port, 
      negative_inputs_0_35_port, negative_inputs_0_34_port, 
      negative_inputs_0_33_port, negative_inputs_0_32_port, 
      negative_inputs_0_31_port, negative_inputs_0_30_port, 
      negative_inputs_0_29_port, negative_inputs_0_28_port, 
      negative_inputs_0_27_port, negative_inputs_0_26_port, 
      negative_inputs_0_25_port, negative_inputs_0_24_port, 
      negative_inputs_0_23_port, negative_inputs_0_22_port, 
      negative_inputs_0_21_port, negative_inputs_0_20_port, 
      negative_inputs_0_19_port, negative_inputs_0_18_port, 
      negative_inputs_0_17_port, negative_inputs_0_16_port, 
      negative_inputs_0_15_port, negative_inputs_0_14_port, 
      negative_inputs_0_13_port, negative_inputs_0_12_port, 
      negative_inputs_0_11_port, negative_inputs_0_10_port, 
      negative_inputs_0_9_port, negative_inputs_0_8_port, 
      negative_inputs_0_7_port, negative_inputs_0_6_port, 
      negative_inputs_0_5_port, negative_inputs_0_4_port, 
      negative_inputs_0_3_port, negative_inputs_0_2_port, 
      negative_inputs_0_1_port, negative_inputs_0_0_port, 
      positive_inputs_8_63_port, positive_inputs_8_62_port, 
      positive_inputs_8_61_port, positive_inputs_8_60_port, 
      positive_inputs_8_59_port, positive_inputs_8_58_port, 
      positive_inputs_8_57_port, positive_inputs_8_56_port, 
      positive_inputs_8_55_port, positive_inputs_8_54_port, 
      positive_inputs_8_53_port, positive_inputs_8_52_port, 
      positive_inputs_8_51_port, positive_inputs_8_50_port, 
      positive_inputs_8_49_port, positive_inputs_8_48_port, 
      positive_inputs_8_47_port, positive_inputs_8_46_port, 
      positive_inputs_8_45_port, positive_inputs_8_44_port, 
      positive_inputs_8_43_port, positive_inputs_8_42_port, 
      positive_inputs_8_41_port, positive_inputs_8_40_port, 
      positive_inputs_8_39_port, positive_inputs_8_38_port, 
      positive_inputs_8_37_port, positive_inputs_8_36_port, 
      positive_inputs_8_35_port, positive_inputs_8_34_port, 
      positive_inputs_8_33_port, positive_inputs_8_32_port, 
      positive_inputs_8_31_port, positive_inputs_8_30_port, 
      positive_inputs_8_29_port, positive_inputs_8_28_port, 
      positive_inputs_8_27_port, positive_inputs_8_26_port, 
      positive_inputs_8_25_port, positive_inputs_8_24_port, 
      positive_inputs_8_23_port, positive_inputs_8_22_port, 
      positive_inputs_8_21_port, positive_inputs_8_20_port, 
      positive_inputs_8_19_port, positive_inputs_8_18_port, 
      positive_inputs_8_17_port, positive_inputs_8_16_port, 
      positive_inputs_8_15_port, positive_inputs_8_14_port, 
      positive_inputs_8_13_port, positive_inputs_8_12_port, 
      positive_inputs_8_11_port, positive_inputs_8_10_port, 
      positive_inputs_8_9_port, positive_inputs_8_8_port, 
      positive_inputs_8_7_port, positive_inputs_8_6_port, 
      positive_inputs_8_5_port, positive_inputs_8_4_port, 
      positive_inputs_8_3_port, positive_inputs_8_2_port, 
      positive_inputs_8_1_port, positive_inputs_7_63_port, 
      positive_inputs_7_62_port, positive_inputs_7_61_port, 
      positive_inputs_7_60_port, positive_inputs_7_59_port, 
      positive_inputs_7_58_port, positive_inputs_7_57_port, 
      positive_inputs_7_56_port, positive_inputs_7_55_port, 
      positive_inputs_7_54_port, positive_inputs_7_53_port, 
      positive_inputs_7_52_port, positive_inputs_7_51_port, 
      positive_inputs_7_50_port, positive_inputs_7_49_port, 
      positive_inputs_7_48_port, positive_inputs_7_47_port, 
      positive_inputs_7_46_port, positive_inputs_7_45_port, 
      positive_inputs_7_44_port, positive_inputs_7_43_port, 
      positive_inputs_7_42_port, positive_inputs_7_41_port, 
      positive_inputs_7_40_port, positive_inputs_7_39_port, 
      positive_inputs_7_38_port, positive_inputs_7_37_port, 
      positive_inputs_7_36_port, positive_inputs_7_35_port, 
      positive_inputs_7_34_port, positive_inputs_7_33_port, 
      positive_inputs_7_32_port, positive_inputs_7_31_port, 
      positive_inputs_7_30_port, positive_inputs_7_29_port, 
      positive_inputs_7_28_port, positive_inputs_7_27_port, 
      positive_inputs_7_26_port, positive_inputs_7_25_port, 
      positive_inputs_7_24_port, positive_inputs_7_23_port, 
      positive_inputs_7_22_port, positive_inputs_7_21_port, 
      positive_inputs_7_20_port, positive_inputs_7_19_port, 
      positive_inputs_7_18_port, positive_inputs_7_17_port, 
      positive_inputs_7_16_port, positive_inputs_7_15_port, 
      positive_inputs_7_14_port, positive_inputs_7_13_port, 
      positive_inputs_7_12_port, positive_inputs_7_11_port, 
      positive_inputs_7_10_port, positive_inputs_7_9_port, 
      positive_inputs_7_8_port, positive_inputs_7_7_port, 
      positive_inputs_7_6_port, positive_inputs_7_5_port, 
      positive_inputs_7_4_port, positive_inputs_7_3_port, 
      positive_inputs_7_2_port, positive_inputs_7_1_port, 
      positive_inputs_6_63_port, positive_inputs_6_62_port, 
      positive_inputs_6_61_port, positive_inputs_6_60_port, 
      positive_inputs_6_59_port, positive_inputs_6_58_port, 
      positive_inputs_6_57_port, positive_inputs_6_56_port, 
      positive_inputs_6_55_port, positive_inputs_6_54_port, 
      positive_inputs_6_53_port, positive_inputs_6_52_port, 
      positive_inputs_6_51_port, positive_inputs_6_50_port, 
      positive_inputs_6_49_port, positive_inputs_6_48_port, 
      positive_inputs_6_47_port, positive_inputs_6_46_port, 
      positive_inputs_6_45_port, positive_inputs_6_44_port, 
      positive_inputs_6_43_port, positive_inputs_6_42_port, 
      positive_inputs_6_41_port, positive_inputs_6_40_port, 
      positive_inputs_6_39_port, positive_inputs_6_38_port, 
      positive_inputs_6_37_port, positive_inputs_6_36_port, 
      positive_inputs_6_35_port, positive_inputs_6_34_port, 
      positive_inputs_6_33_port, positive_inputs_6_32_port, 
      positive_inputs_6_31_port, positive_inputs_6_30_port, 
      positive_inputs_6_29_port, positive_inputs_6_28_port, 
      positive_inputs_6_27_port, positive_inputs_6_26_port, 
      positive_inputs_6_25_port, positive_inputs_6_24_port, 
      positive_inputs_6_23_port, positive_inputs_6_22_port, 
      positive_inputs_6_21_port, positive_inputs_6_20_port, 
      positive_inputs_6_19_port, positive_inputs_6_18_port, 
      positive_inputs_6_17_port, positive_inputs_6_16_port, 
      positive_inputs_6_15_port, positive_inputs_6_14_port, 
      positive_inputs_6_13_port, positive_inputs_6_12_port, 
      positive_inputs_6_11_port, positive_inputs_6_10_port, 
      positive_inputs_6_9_port, positive_inputs_6_8_port, 
      positive_inputs_6_7_port, positive_inputs_6_6_port, 
      positive_inputs_6_5_port, positive_inputs_6_4_port, 
      positive_inputs_6_3_port, positive_inputs_6_2_port, 
      positive_inputs_6_1_port, positive_inputs_5_63_port, 
      positive_inputs_5_62_port, positive_inputs_5_61_port, 
      positive_inputs_5_60_port, positive_inputs_5_59_port, 
      positive_inputs_5_58_port, positive_inputs_5_57_port, 
      positive_inputs_5_56_port, positive_inputs_5_55_port, 
      positive_inputs_5_54_port, positive_inputs_5_53_port, 
      positive_inputs_5_52_port, positive_inputs_5_51_port, 
      positive_inputs_5_50_port, positive_inputs_5_49_port, 
      positive_inputs_5_48_port, positive_inputs_5_47_port, 
      positive_inputs_5_46_port, positive_inputs_5_45_port, 
      positive_inputs_5_44_port, positive_inputs_5_43_port, 
      positive_inputs_5_42_port, positive_inputs_5_41_port, 
      positive_inputs_5_40_port, positive_inputs_5_39_port, 
      positive_inputs_5_38_port, positive_inputs_5_37_port, 
      positive_inputs_5_36_port, positive_inputs_5_35_port, 
      positive_inputs_5_34_port, positive_inputs_5_33_port, 
      positive_inputs_5_32_port, positive_inputs_5_31_port, 
      positive_inputs_5_30_port, positive_inputs_5_29_port, 
      positive_inputs_5_28_port, positive_inputs_5_27_port, 
      positive_inputs_5_26_port, positive_inputs_5_25_port, 
      positive_inputs_5_24_port, positive_inputs_5_23_port, 
      positive_inputs_5_22_port, positive_inputs_5_21_port, 
      positive_inputs_5_20_port, positive_inputs_5_19_port, 
      positive_inputs_5_18_port, positive_inputs_5_17_port, 
      positive_inputs_5_16_port, positive_inputs_5_15_port, 
      positive_inputs_5_14_port, positive_inputs_5_13_port, 
      positive_inputs_5_12_port, positive_inputs_5_11_port, 
      positive_inputs_5_10_port, positive_inputs_5_9_port, 
      positive_inputs_5_8_port, positive_inputs_5_7_port, 
      positive_inputs_5_6_port, positive_inputs_5_5_port, 
      positive_inputs_5_4_port, positive_inputs_5_3_port, 
      positive_inputs_5_2_port, positive_inputs_5_1_port, 
      positive_inputs_4_63_port, positive_inputs_4_62_port, 
      positive_inputs_4_61_port, positive_inputs_4_60_port, 
      positive_inputs_4_59_port, positive_inputs_4_58_port, 
      positive_inputs_4_57_port, positive_inputs_4_56_port, 
      positive_inputs_4_55_port, positive_inputs_4_54_port, 
      positive_inputs_4_53_port, positive_inputs_4_52_port, 
      positive_inputs_4_51_port, positive_inputs_4_50_port, 
      positive_inputs_4_49_port, positive_inputs_4_48_port, 
      positive_inputs_4_47_port, positive_inputs_4_46_port, 
      positive_inputs_4_45_port, positive_inputs_4_44_port, 
      positive_inputs_4_43_port, positive_inputs_4_42_port, 
      positive_inputs_4_41_port, positive_inputs_4_40_port, 
      positive_inputs_4_39_port, positive_inputs_4_38_port, 
      positive_inputs_4_37_port, positive_inputs_4_36_port, 
      positive_inputs_4_35_port, positive_inputs_4_34_port, 
      positive_inputs_4_33_port, positive_inputs_4_32_port, 
      positive_inputs_4_31_port, positive_inputs_4_30_port, 
      positive_inputs_4_29_port, positive_inputs_4_28_port, 
      positive_inputs_4_27_port, positive_inputs_4_26_port, 
      positive_inputs_4_25_port, positive_inputs_4_24_port, 
      positive_inputs_4_23_port, positive_inputs_4_22_port, 
      positive_inputs_4_21_port, positive_inputs_4_20_port, 
      positive_inputs_4_19_port, positive_inputs_4_18_port, 
      positive_inputs_4_17_port, positive_inputs_4_16_port, 
      positive_inputs_4_15_port, positive_inputs_4_14_port, 
      positive_inputs_4_13_port, positive_inputs_4_12_port, 
      positive_inputs_4_11_port, positive_inputs_4_10_port, 
      positive_inputs_4_9_port, positive_inputs_4_8_port, 
      positive_inputs_4_7_port, positive_inputs_4_6_port, 
      positive_inputs_4_5_port, positive_inputs_4_4_port, 
      positive_inputs_4_3_port, positive_inputs_4_2_port, 
      positive_inputs_4_1_port, positive_inputs_3_63_port, 
      positive_inputs_3_62_port, positive_inputs_3_61_port, 
      positive_inputs_3_60_port, positive_inputs_3_59_port, 
      positive_inputs_3_58_port, positive_inputs_3_57_port, 
      positive_inputs_3_56_port, positive_inputs_3_55_port, 
      positive_inputs_3_54_port, positive_inputs_3_53_port, 
      positive_inputs_3_52_port, positive_inputs_3_51_port, 
      positive_inputs_3_50_port, positive_inputs_3_49_port, 
      positive_inputs_3_48_port, positive_inputs_3_47_port, 
      positive_inputs_3_46_port, positive_inputs_3_45_port, 
      positive_inputs_3_44_port, positive_inputs_3_43_port, 
      positive_inputs_3_42_port, positive_inputs_3_41_port, 
      positive_inputs_3_40_port, positive_inputs_3_39_port, 
      positive_inputs_3_38_port, positive_inputs_3_37_port, 
      positive_inputs_3_36_port, positive_inputs_3_35_port, 
      positive_inputs_3_34_port, positive_inputs_3_33_port, 
      positive_inputs_3_32_port, positive_inputs_3_31_port, 
      positive_inputs_3_30_port, positive_inputs_3_29_port, 
      positive_inputs_3_28_port, positive_inputs_3_27_port, 
      positive_inputs_3_26_port, positive_inputs_3_25_port, 
      positive_inputs_3_24_port, positive_inputs_3_23_port, 
      positive_inputs_3_22_port, positive_inputs_3_21_port, 
      positive_inputs_3_20_port, positive_inputs_3_19_port, 
      positive_inputs_3_18_port, positive_inputs_3_17_port, 
      positive_inputs_3_16_port, positive_inputs_3_15_port, 
      positive_inputs_3_14_port, positive_inputs_3_13_port, 
      positive_inputs_3_12_port, positive_inputs_3_11_port, 
      positive_inputs_3_10_port, positive_inputs_3_9_port, 
      positive_inputs_3_8_port, positive_inputs_3_7_port, 
      positive_inputs_3_6_port, positive_inputs_3_5_port, 
      positive_inputs_3_4_port, positive_inputs_3_3_port, 
      positive_inputs_3_2_port, positive_inputs_3_1_port, 
      positive_inputs_2_63_port, positive_inputs_2_62_port, 
      positive_inputs_2_61_port, positive_inputs_2_60_port, 
      positive_inputs_2_59_port, positive_inputs_2_58_port, 
      positive_inputs_2_57_port, positive_inputs_2_56_port, 
      positive_inputs_2_55_port, positive_inputs_2_54_port, 
      positive_inputs_2_53_port, positive_inputs_2_52_port, 
      positive_inputs_2_51_port, positive_inputs_2_50_port, 
      positive_inputs_2_49_port, positive_inputs_2_48_port, 
      positive_inputs_2_47_port, positive_inputs_2_46_port, 
      positive_inputs_2_45_port, positive_inputs_2_44_port, 
      positive_inputs_2_43_port, positive_inputs_2_42_port, 
      positive_inputs_2_41_port, positive_inputs_2_40_port, 
      positive_inputs_2_39_port, positive_inputs_2_38_port, 
      positive_inputs_2_37_port, positive_inputs_2_36_port, 
      positive_inputs_2_35_port, positive_inputs_2_34_port, 
      positive_inputs_2_33_port, positive_inputs_2_32_port, 
      positive_inputs_2_31_port, positive_inputs_2_30_port, 
      positive_inputs_2_29_port, positive_inputs_2_28_port, 
      positive_inputs_2_27_port, positive_inputs_2_26_port, 
      positive_inputs_2_25_port, positive_inputs_2_24_port, 
      positive_inputs_2_23_port, positive_inputs_2_22_port, 
      positive_inputs_2_21_port, positive_inputs_2_20_port, 
      positive_inputs_2_19_port, positive_inputs_2_18_port, 
      positive_inputs_2_17_port, positive_inputs_2_16_port, 
      positive_inputs_2_15_port, positive_inputs_2_14_port, 
      positive_inputs_2_13_port, positive_inputs_2_12_port, 
      positive_inputs_2_11_port, positive_inputs_2_10_port, 
      positive_inputs_2_9_port, positive_inputs_2_8_port, 
      positive_inputs_2_7_port, positive_inputs_2_6_port, 
      positive_inputs_2_5_port, positive_inputs_2_4_port, 
      positive_inputs_2_3_port, positive_inputs_2_2_port, 
      positive_inputs_2_1_port, positive_inputs_1_63_port, 
      positive_inputs_1_62_port, positive_inputs_1_61_port, 
      positive_inputs_1_60_port, positive_inputs_1_59_port, 
      positive_inputs_1_58_port, positive_inputs_1_57_port, 
      positive_inputs_1_56_port, positive_inputs_1_55_port, 
      positive_inputs_1_54_port, positive_inputs_1_53_port, 
      positive_inputs_1_52_port, positive_inputs_1_51_port, 
      positive_inputs_1_50_port, positive_inputs_1_49_port, 
      positive_inputs_1_48_port, positive_inputs_1_47_port, 
      positive_inputs_1_46_port, positive_inputs_1_45_port, 
      positive_inputs_1_44_port, positive_inputs_1_43_port, 
      positive_inputs_1_42_port, positive_inputs_1_41_port, 
      positive_inputs_1_40_port, positive_inputs_1_39_port, 
      positive_inputs_1_38_port, positive_inputs_1_37_port, 
      positive_inputs_1_36_port, positive_inputs_1_35_port, 
      positive_inputs_1_34_port, positive_inputs_1_33_port, 
      positive_inputs_1_32_port, positive_inputs_1_31_port, 
      positive_inputs_1_30_port, positive_inputs_1_29_port, 
      positive_inputs_1_28_port, positive_inputs_1_27_port, 
      positive_inputs_1_26_port, positive_inputs_1_25_port, 
      positive_inputs_1_24_port, positive_inputs_1_23_port, 
      positive_inputs_1_22_port, positive_inputs_1_21_port, 
      positive_inputs_1_20_port, positive_inputs_1_19_port, 
      positive_inputs_1_18_port, positive_inputs_1_17_port, 
      positive_inputs_1_16_port, positive_inputs_1_15_port, 
      positive_inputs_1_14_port, positive_inputs_1_13_port, 
      positive_inputs_1_12_port, positive_inputs_1_11_port, 
      positive_inputs_1_10_port, positive_inputs_1_9_port, 
      positive_inputs_1_8_port, positive_inputs_1_7_port, 
      positive_inputs_1_6_port, positive_inputs_1_5_port, 
      positive_inputs_1_4_port, positive_inputs_1_3_port, 
      positive_inputs_1_2_port, positive_inputs_1_1_port, 
      positive_inputs_16_63_port, positive_inputs_16_62_port, 
      positive_inputs_16_61_port, positive_inputs_16_60_port, 
      positive_inputs_16_59_port, positive_inputs_16_58_port, 
      positive_inputs_16_57_port, positive_inputs_16_56_port, 
      positive_inputs_16_55_port, positive_inputs_16_54_port, 
      positive_inputs_16_53_port, positive_inputs_16_52_port, 
      positive_inputs_16_51_port, positive_inputs_16_50_port, 
      positive_inputs_16_49_port, positive_inputs_16_48_port, 
      positive_inputs_16_47_port, positive_inputs_16_46_port, 
      positive_inputs_16_45_port, positive_inputs_16_44_port, 
      positive_inputs_16_43_port, positive_inputs_16_42_port, 
      positive_inputs_16_41_port, positive_inputs_16_40_port, 
      positive_inputs_16_39_port, positive_inputs_16_38_port, 
      positive_inputs_16_37_port, positive_inputs_16_36_port, 
      positive_inputs_16_35_port, positive_inputs_16_34_port, 
      positive_inputs_16_33_port, positive_inputs_16_32_port, 
      positive_inputs_16_31_port, positive_inputs_16_30_port, 
      positive_inputs_16_29_port, positive_inputs_16_28_port, 
      positive_inputs_16_27_port, positive_inputs_16_26_port, 
      positive_inputs_16_25_port, positive_inputs_16_24_port, 
      positive_inputs_16_23_port, positive_inputs_16_22_port, 
      positive_inputs_16_21_port, positive_inputs_16_20_port, 
      positive_inputs_16_19_port, positive_inputs_16_18_port, 
      positive_inputs_16_17_port, positive_inputs_16_16_port, 
      positive_inputs_16_15_port, positive_inputs_16_14_port, 
      positive_inputs_16_13_port, positive_inputs_16_12_port, 
      positive_inputs_16_11_port, positive_inputs_16_10_port, 
      positive_inputs_16_9_port, positive_inputs_16_8_port, 
      positive_inputs_16_7_port, positive_inputs_16_6_port, 
      positive_inputs_16_5_port, positive_inputs_16_4_port, 
      positive_inputs_16_3_port, positive_inputs_16_2_port, 
      positive_inputs_16_1_port, positive_inputs_15_63_port, 
      positive_inputs_15_62_port, positive_inputs_15_61_port, 
      positive_inputs_15_60_port, positive_inputs_15_59_port, 
      positive_inputs_15_58_port, positive_inputs_15_57_port, 
      positive_inputs_15_56_port, positive_inputs_15_55_port, 
      positive_inputs_15_54_port, positive_inputs_15_53_port, 
      positive_inputs_15_52_port, positive_inputs_15_51_port, 
      positive_inputs_15_50_port, positive_inputs_15_49_port, 
      positive_inputs_15_48_port, positive_inputs_15_47_port, 
      positive_inputs_15_46_port, positive_inputs_15_45_port, 
      positive_inputs_15_44_port, positive_inputs_15_43_port, 
      positive_inputs_15_42_port, positive_inputs_15_41_port, 
      positive_inputs_15_40_port, positive_inputs_15_39_port, 
      positive_inputs_15_38_port, positive_inputs_15_37_port, 
      positive_inputs_15_36_port, positive_inputs_15_35_port, 
      positive_inputs_15_34_port, positive_inputs_15_33_port, 
      positive_inputs_15_32_port, positive_inputs_15_31_port, 
      positive_inputs_15_30_port, positive_inputs_15_29_port, 
      positive_inputs_15_28_port, positive_inputs_15_27_port, 
      positive_inputs_15_26_port, positive_inputs_15_25_port, 
      positive_inputs_15_24_port, positive_inputs_15_23_port, 
      positive_inputs_15_22_port, positive_inputs_15_21_port, 
      positive_inputs_15_20_port, positive_inputs_15_19_port, 
      positive_inputs_15_18_port, positive_inputs_15_17_port, 
      positive_inputs_15_16_port, positive_inputs_15_15_port, 
      positive_inputs_15_14_port, positive_inputs_15_13_port, 
      positive_inputs_15_12_port, positive_inputs_15_11_port, 
      positive_inputs_15_10_port, positive_inputs_15_9_port, 
      positive_inputs_15_8_port, positive_inputs_15_7_port, 
      positive_inputs_15_6_port, positive_inputs_15_5_port, 
      positive_inputs_15_4_port, positive_inputs_15_3_port, 
      positive_inputs_15_2_port, positive_inputs_15_1_port, 
      positive_inputs_14_63_port, positive_inputs_14_62_port, 
      positive_inputs_14_61_port, positive_inputs_14_60_port, 
      positive_inputs_14_59_port, positive_inputs_14_58_port, 
      positive_inputs_14_57_port, positive_inputs_14_56_port, 
      positive_inputs_14_55_port, positive_inputs_14_54_port, 
      positive_inputs_14_53_port, positive_inputs_14_52_port, 
      positive_inputs_14_51_port, positive_inputs_14_50_port, 
      positive_inputs_14_49_port, positive_inputs_14_48_port, 
      positive_inputs_14_47_port, positive_inputs_14_46_port, 
      positive_inputs_14_45_port, positive_inputs_14_44_port, 
      positive_inputs_14_43_port, positive_inputs_14_42_port, 
      positive_inputs_14_41_port, positive_inputs_14_40_port, 
      positive_inputs_14_39_port, positive_inputs_14_38_port, 
      positive_inputs_14_37_port, positive_inputs_14_36_port, 
      positive_inputs_14_35_port, positive_inputs_14_34_port, 
      positive_inputs_14_33_port, positive_inputs_14_32_port, 
      positive_inputs_14_31_port, positive_inputs_14_30_port, 
      positive_inputs_14_29_port, positive_inputs_14_28_port, 
      positive_inputs_14_27_port, positive_inputs_14_26_port, 
      positive_inputs_14_25_port, positive_inputs_14_24_port, 
      positive_inputs_14_23_port, positive_inputs_14_22_port, 
      positive_inputs_14_21_port, positive_inputs_14_20_port, 
      positive_inputs_14_19_port, positive_inputs_14_18_port, 
      positive_inputs_14_17_port, positive_inputs_14_16_port, 
      positive_inputs_14_15_port, positive_inputs_14_14_port, 
      positive_inputs_14_13_port, positive_inputs_14_12_port, 
      positive_inputs_14_11_port, positive_inputs_14_10_port, 
      positive_inputs_14_9_port, positive_inputs_14_8_port, 
      positive_inputs_14_7_port, positive_inputs_14_6_port, 
      positive_inputs_14_5_port, positive_inputs_14_4_port, 
      positive_inputs_14_3_port, positive_inputs_14_2_port, 
      positive_inputs_14_1_port, positive_inputs_13_63_port, 
      positive_inputs_13_62_port, positive_inputs_13_61_port, 
      positive_inputs_13_60_port, positive_inputs_13_59_port, 
      positive_inputs_13_58_port, positive_inputs_13_57_port, 
      positive_inputs_13_56_port, positive_inputs_13_55_port, 
      positive_inputs_13_54_port, positive_inputs_13_53_port, 
      positive_inputs_13_52_port, positive_inputs_13_51_port, 
      positive_inputs_13_50_port, positive_inputs_13_49_port, 
      positive_inputs_13_48_port, positive_inputs_13_47_port, 
      positive_inputs_13_46_port, positive_inputs_13_45_port, 
      positive_inputs_13_44_port, positive_inputs_13_43_port, 
      positive_inputs_13_42_port, positive_inputs_13_41_port, 
      positive_inputs_13_40_port, positive_inputs_13_39_port, 
      positive_inputs_13_38_port, positive_inputs_13_37_port, 
      positive_inputs_13_36_port, positive_inputs_13_35_port, 
      positive_inputs_13_34_port, positive_inputs_13_33_port, 
      positive_inputs_13_32_port, positive_inputs_13_31_port, 
      positive_inputs_13_30_port, positive_inputs_13_29_port, 
      positive_inputs_13_28_port, positive_inputs_13_27_port, 
      positive_inputs_13_26_port, positive_inputs_13_25_port, 
      positive_inputs_13_24_port, positive_inputs_13_23_port, 
      positive_inputs_13_22_port, positive_inputs_13_21_port, 
      positive_inputs_13_20_port, positive_inputs_13_19_port, 
      positive_inputs_13_18_port, positive_inputs_13_17_port, 
      positive_inputs_13_16_port, positive_inputs_13_15_port, 
      positive_inputs_13_14_port, positive_inputs_13_13_port, 
      positive_inputs_13_12_port, positive_inputs_13_11_port, 
      positive_inputs_13_10_port, positive_inputs_13_9_port, 
      positive_inputs_13_8_port, positive_inputs_13_7_port, 
      positive_inputs_13_6_port, positive_inputs_13_5_port, 
      positive_inputs_13_4_port, positive_inputs_13_3_port, 
      positive_inputs_13_2_port, positive_inputs_13_1_port, 
      positive_inputs_12_63_port, positive_inputs_12_62_port, 
      positive_inputs_12_61_port, positive_inputs_12_60_port, 
      positive_inputs_12_59_port, positive_inputs_12_58_port, 
      positive_inputs_12_57_port, positive_inputs_12_56_port, 
      positive_inputs_12_55_port, positive_inputs_12_54_port, 
      positive_inputs_12_53_port, positive_inputs_12_52_port, 
      positive_inputs_12_51_port, positive_inputs_12_50_port, 
      positive_inputs_12_49_port, positive_inputs_12_48_port, 
      positive_inputs_12_47_port, positive_inputs_12_46_port, 
      positive_inputs_12_45_port, positive_inputs_12_44_port, 
      positive_inputs_12_43_port, positive_inputs_12_42_port, 
      positive_inputs_12_41_port, positive_inputs_12_40_port, 
      positive_inputs_12_39_port, positive_inputs_12_38_port, 
      positive_inputs_12_37_port, positive_inputs_12_36_port, 
      positive_inputs_12_35_port, positive_inputs_12_34_port, 
      positive_inputs_12_33_port, positive_inputs_12_32_port, 
      positive_inputs_12_31_port, positive_inputs_12_30_port, 
      positive_inputs_12_29_port, positive_inputs_12_28_port, 
      positive_inputs_12_27_port, positive_inputs_12_26_port, 
      positive_inputs_12_25_port, positive_inputs_12_24_port, 
      positive_inputs_12_23_port, positive_inputs_12_22_port, 
      positive_inputs_12_21_port, positive_inputs_12_20_port, 
      positive_inputs_12_19_port, positive_inputs_12_18_port, 
      positive_inputs_12_17_port, positive_inputs_12_16_port, 
      positive_inputs_12_15_port, positive_inputs_12_14_port, 
      positive_inputs_12_13_port, positive_inputs_12_12_port, 
      positive_inputs_12_11_port, positive_inputs_12_10_port, 
      positive_inputs_12_9_port, positive_inputs_12_8_port, 
      positive_inputs_12_7_port, positive_inputs_12_6_port, 
      positive_inputs_12_5_port, positive_inputs_12_4_port, 
      positive_inputs_12_3_port, positive_inputs_12_2_port, 
      positive_inputs_12_1_port, positive_inputs_11_63_port, 
      positive_inputs_11_62_port, positive_inputs_11_61_port, 
      positive_inputs_11_60_port, positive_inputs_11_59_port, 
      positive_inputs_11_58_port, positive_inputs_11_57_port, 
      positive_inputs_11_56_port, positive_inputs_11_55_port, 
      positive_inputs_11_54_port, positive_inputs_11_53_port, 
      positive_inputs_11_52_port, positive_inputs_11_51_port, 
      positive_inputs_11_50_port, positive_inputs_11_49_port, 
      positive_inputs_11_48_port, positive_inputs_11_47_port, 
      positive_inputs_11_46_port, positive_inputs_11_45_port, 
      positive_inputs_11_44_port, positive_inputs_11_43_port, 
      positive_inputs_11_42_port, positive_inputs_11_41_port, 
      positive_inputs_11_40_port, positive_inputs_11_39_port, 
      positive_inputs_11_38_port, positive_inputs_11_37_port, 
      positive_inputs_11_36_port, positive_inputs_11_35_port, 
      positive_inputs_11_34_port, positive_inputs_11_33_port, 
      positive_inputs_11_32_port, positive_inputs_11_31_port, 
      positive_inputs_11_30_port, positive_inputs_11_29_port, 
      positive_inputs_11_28_port, positive_inputs_11_27_port, 
      positive_inputs_11_26_port, positive_inputs_11_25_port, 
      positive_inputs_11_24_port, positive_inputs_11_23_port, 
      positive_inputs_11_22_port, positive_inputs_11_21_port, 
      positive_inputs_11_20_port, positive_inputs_11_19_port, 
      positive_inputs_11_18_port, positive_inputs_11_17_port, 
      positive_inputs_11_16_port, positive_inputs_11_15_port, 
      positive_inputs_11_14_port, positive_inputs_11_13_port, 
      positive_inputs_11_12_port, positive_inputs_11_11_port, 
      positive_inputs_11_10_port, positive_inputs_11_9_port, 
      positive_inputs_11_8_port, positive_inputs_11_7_port, 
      positive_inputs_11_6_port, positive_inputs_11_5_port, 
      positive_inputs_11_4_port, positive_inputs_11_3_port, 
      positive_inputs_11_2_port, positive_inputs_11_1_port, 
      positive_inputs_10_63_port, positive_inputs_10_62_port, 
      positive_inputs_10_61_port, positive_inputs_10_60_port, 
      positive_inputs_10_59_port, positive_inputs_10_58_port, 
      positive_inputs_10_57_port, positive_inputs_10_56_port, 
      positive_inputs_10_55_port, positive_inputs_10_54_port, 
      positive_inputs_10_53_port, positive_inputs_10_52_port, 
      positive_inputs_10_51_port, positive_inputs_10_50_port, 
      positive_inputs_10_49_port, positive_inputs_10_48_port, 
      positive_inputs_10_47_port, positive_inputs_10_46_port, 
      positive_inputs_10_45_port, positive_inputs_10_44_port, 
      positive_inputs_10_43_port, positive_inputs_10_42_port, 
      positive_inputs_10_41_port, positive_inputs_10_40_port, 
      positive_inputs_10_39_port, positive_inputs_10_38_port, 
      positive_inputs_10_37_port, positive_inputs_10_36_port, 
      positive_inputs_10_35_port, positive_inputs_10_34_port, 
      positive_inputs_10_33_port, positive_inputs_10_32_port, 
      positive_inputs_10_31_port, positive_inputs_10_30_port, 
      positive_inputs_10_29_port, positive_inputs_10_28_port, 
      positive_inputs_10_27_port, positive_inputs_10_26_port, 
      positive_inputs_10_25_port, positive_inputs_10_24_port, 
      positive_inputs_10_23_port, positive_inputs_10_22_port, 
      positive_inputs_10_21_port, positive_inputs_10_20_port, 
      positive_inputs_10_19_port, positive_inputs_10_18_port, 
      positive_inputs_10_17_port, positive_inputs_10_16_port, 
      positive_inputs_10_15_port, positive_inputs_10_14_port, 
      positive_inputs_10_13_port, positive_inputs_10_12_port, 
      positive_inputs_10_11_port, positive_inputs_10_10_port, 
      positive_inputs_10_9_port, positive_inputs_10_8_port, 
      positive_inputs_10_7_port, positive_inputs_10_6_port, 
      positive_inputs_10_5_port, positive_inputs_10_4_port, 
      positive_inputs_10_3_port, positive_inputs_10_2_port, 
      positive_inputs_10_1_port, positive_inputs_9_63_port, 
      positive_inputs_9_62_port, positive_inputs_9_61_port, 
      positive_inputs_9_60_port, positive_inputs_9_59_port, 
      positive_inputs_9_58_port, positive_inputs_9_57_port, 
      positive_inputs_9_56_port, positive_inputs_9_55_port, 
      positive_inputs_9_54_port, positive_inputs_9_53_port, 
      positive_inputs_9_52_port, positive_inputs_9_51_port, 
      positive_inputs_9_50_port, positive_inputs_9_49_port, 
      positive_inputs_9_48_port, positive_inputs_9_47_port, 
      positive_inputs_9_46_port, positive_inputs_9_45_port, 
      positive_inputs_9_44_port, positive_inputs_9_43_port, 
      positive_inputs_9_42_port, positive_inputs_9_41_port, 
      positive_inputs_9_40_port, positive_inputs_9_39_port, 
      positive_inputs_9_38_port, positive_inputs_9_37_port, 
      positive_inputs_9_36_port, positive_inputs_9_35_port, 
      positive_inputs_9_34_port, positive_inputs_9_33_port, 
      positive_inputs_9_32_port, positive_inputs_9_31_port, 
      positive_inputs_9_30_port, positive_inputs_9_29_port, 
      positive_inputs_9_28_port, positive_inputs_9_27_port, 
      positive_inputs_9_26_port, positive_inputs_9_25_port, 
      positive_inputs_9_24_port, positive_inputs_9_23_port, 
      positive_inputs_9_22_port, positive_inputs_9_21_port, 
      positive_inputs_9_20_port, positive_inputs_9_19_port, 
      positive_inputs_9_18_port, positive_inputs_9_17_port, 
      positive_inputs_9_16_port, positive_inputs_9_15_port, 
      positive_inputs_9_14_port, positive_inputs_9_13_port, 
      positive_inputs_9_12_port, positive_inputs_9_11_port, 
      positive_inputs_9_10_port, positive_inputs_9_9_port, 
      positive_inputs_9_8_port, positive_inputs_9_7_port, 
      positive_inputs_9_6_port, positive_inputs_9_5_port, 
      positive_inputs_9_4_port, positive_inputs_9_3_port, 
      positive_inputs_9_2_port, positive_inputs_9_1_port, 
      positive_inputs_24_63_port, positive_inputs_24_62_port, 
      positive_inputs_24_61_port, positive_inputs_24_60_port, 
      positive_inputs_24_59_port, positive_inputs_24_58_port, 
      positive_inputs_24_57_port, positive_inputs_24_56_port, 
      positive_inputs_24_55_port, positive_inputs_24_54_port, 
      positive_inputs_24_53_port, positive_inputs_24_52_port, 
      positive_inputs_24_51_port, positive_inputs_24_50_port, 
      positive_inputs_24_49_port, positive_inputs_24_48_port, 
      positive_inputs_24_47_port, positive_inputs_24_46_port, 
      positive_inputs_24_45_port, positive_inputs_24_44_port, 
      positive_inputs_24_43_port, positive_inputs_24_42_port, 
      positive_inputs_24_41_port, positive_inputs_24_40_port, 
      positive_inputs_24_39_port, positive_inputs_24_38_port, 
      positive_inputs_24_37_port, positive_inputs_24_36_port, 
      positive_inputs_24_35_port, positive_inputs_24_34_port, 
      positive_inputs_24_33_port, positive_inputs_24_32_port, 
      positive_inputs_24_31_port, positive_inputs_24_30_port, 
      positive_inputs_24_29_port, positive_inputs_24_28_port, 
      positive_inputs_24_27_port, positive_inputs_24_26_port, 
      positive_inputs_24_25_port, positive_inputs_24_24_port, 
      positive_inputs_24_23_port, positive_inputs_24_22_port, 
      positive_inputs_24_21_port, positive_inputs_24_20_port, 
      positive_inputs_24_19_port, positive_inputs_24_18_port, 
      positive_inputs_24_17_port, positive_inputs_24_16_port, 
      positive_inputs_24_15_port, positive_inputs_24_14_port, 
      positive_inputs_24_13_port, positive_inputs_24_12_port, 
      positive_inputs_24_11_port, positive_inputs_24_10_port, 
      positive_inputs_24_9_port, positive_inputs_24_8_port, 
      positive_inputs_24_7_port, positive_inputs_24_6_port, 
      positive_inputs_24_5_port, positive_inputs_24_4_port, 
      positive_inputs_24_3_port, positive_inputs_24_2_port, 
      positive_inputs_24_1_port, positive_inputs_23_63_port, 
      positive_inputs_23_62_port, positive_inputs_23_61_port, 
      positive_inputs_23_60_port, positive_inputs_23_59_port, 
      positive_inputs_23_58_port, positive_inputs_23_57_port, 
      positive_inputs_23_56_port, positive_inputs_23_55_port, 
      positive_inputs_23_54_port, positive_inputs_23_53_port, 
      positive_inputs_23_52_port, positive_inputs_23_51_port, 
      positive_inputs_23_50_port, positive_inputs_23_49_port, 
      positive_inputs_23_48_port, positive_inputs_23_47_port, 
      positive_inputs_23_46_port, positive_inputs_23_45_port, 
      positive_inputs_23_44_port, positive_inputs_23_43_port, 
      positive_inputs_23_42_port, positive_inputs_23_41_port, 
      positive_inputs_23_40_port, positive_inputs_23_39_port, 
      positive_inputs_23_38_port, positive_inputs_23_37_port, 
      positive_inputs_23_36_port, positive_inputs_23_35_port, 
      positive_inputs_23_34_port, positive_inputs_23_33_port, 
      positive_inputs_23_32_port, positive_inputs_23_31_port, 
      positive_inputs_23_30_port, positive_inputs_23_29_port, 
      positive_inputs_23_28_port, positive_inputs_23_27_port, 
      positive_inputs_23_26_port, positive_inputs_23_25_port, 
      positive_inputs_23_24_port, positive_inputs_23_23_port, 
      positive_inputs_23_22_port, positive_inputs_23_21_port, 
      positive_inputs_23_20_port, positive_inputs_23_19_port, 
      positive_inputs_23_18_port, positive_inputs_23_17_port, 
      positive_inputs_23_16_port, positive_inputs_23_15_port, 
      positive_inputs_23_14_port, positive_inputs_23_13_port, 
      positive_inputs_23_12_port, positive_inputs_23_11_port, 
      positive_inputs_23_10_port, positive_inputs_23_9_port, 
      positive_inputs_23_8_port, positive_inputs_23_7_port, 
      positive_inputs_23_6_port, positive_inputs_23_5_port, 
      positive_inputs_23_4_port, positive_inputs_23_3_port, 
      positive_inputs_23_2_port, positive_inputs_23_1_port, 
      positive_inputs_22_63_port, positive_inputs_22_62_port, 
      positive_inputs_22_61_port, positive_inputs_22_60_port, 
      positive_inputs_22_59_port, positive_inputs_22_58_port, 
      positive_inputs_22_57_port, positive_inputs_22_56_port, 
      positive_inputs_22_55_port, positive_inputs_22_54_port, 
      positive_inputs_22_53_port, positive_inputs_22_52_port, 
      positive_inputs_22_51_port, positive_inputs_22_50_port, 
      positive_inputs_22_49_port, positive_inputs_22_48_port, 
      positive_inputs_22_47_port, positive_inputs_22_46_port, 
      positive_inputs_22_45_port, positive_inputs_22_44_port, 
      positive_inputs_22_43_port, positive_inputs_22_42_port, 
      positive_inputs_22_41_port, positive_inputs_22_40_port, 
      positive_inputs_22_39_port, positive_inputs_22_38_port, 
      positive_inputs_22_37_port, positive_inputs_22_36_port, 
      positive_inputs_22_35_port, positive_inputs_22_34_port, 
      positive_inputs_22_33_port, positive_inputs_22_32_port, 
      positive_inputs_22_31_port, positive_inputs_22_30_port, 
      positive_inputs_22_29_port, positive_inputs_22_28_port, 
      positive_inputs_22_27_port, positive_inputs_22_26_port, 
      positive_inputs_22_25_port, positive_inputs_22_24_port, 
      positive_inputs_22_23_port, positive_inputs_22_22_port, 
      positive_inputs_22_21_port, positive_inputs_22_20_port, 
      positive_inputs_22_19_port, positive_inputs_22_18_port, 
      positive_inputs_22_17_port, positive_inputs_22_16_port, 
      positive_inputs_22_15_port, positive_inputs_22_14_port, 
      positive_inputs_22_13_port, positive_inputs_22_12_port, 
      positive_inputs_22_11_port, positive_inputs_22_10_port, 
      positive_inputs_22_9_port, positive_inputs_22_8_port, 
      positive_inputs_22_7_port, positive_inputs_22_6_port, 
      positive_inputs_22_5_port, positive_inputs_22_4_port, 
      positive_inputs_22_3_port, positive_inputs_22_2_port, 
      positive_inputs_22_1_port, positive_inputs_21_63_port, 
      positive_inputs_21_62_port, positive_inputs_21_61_port, 
      positive_inputs_21_60_port, positive_inputs_21_59_port, 
      positive_inputs_21_58_port, positive_inputs_21_57_port, 
      positive_inputs_21_56_port, positive_inputs_21_55_port, 
      positive_inputs_21_54_port, positive_inputs_21_53_port, 
      positive_inputs_21_52_port, positive_inputs_21_51_port, 
      positive_inputs_21_50_port, positive_inputs_21_49_port, 
      positive_inputs_21_48_port, positive_inputs_21_47_port, 
      positive_inputs_21_46_port, positive_inputs_21_45_port, 
      positive_inputs_21_44_port, positive_inputs_21_43_port, 
      positive_inputs_21_42_port, positive_inputs_21_41_port, 
      positive_inputs_21_40_port, positive_inputs_21_39_port, 
      positive_inputs_21_38_port, positive_inputs_21_37_port, 
      positive_inputs_21_36_port, positive_inputs_21_35_port, 
      positive_inputs_21_34_port, positive_inputs_21_33_port, 
      positive_inputs_21_32_port, positive_inputs_21_31_port, 
      positive_inputs_21_30_port, positive_inputs_21_29_port, 
      positive_inputs_21_28_port, positive_inputs_21_27_port, 
      positive_inputs_21_26_port, positive_inputs_21_25_port, 
      positive_inputs_21_24_port, positive_inputs_21_23_port, 
      positive_inputs_21_22_port, positive_inputs_21_21_port, 
      positive_inputs_21_20_port, positive_inputs_21_19_port, 
      positive_inputs_21_18_port, positive_inputs_21_17_port, 
      positive_inputs_21_16_port, positive_inputs_21_15_port, 
      positive_inputs_21_14_port, positive_inputs_21_13_port, 
      positive_inputs_21_12_port, positive_inputs_21_11_port, 
      positive_inputs_21_10_port, positive_inputs_21_9_port, 
      positive_inputs_21_8_port, positive_inputs_21_7_port, 
      positive_inputs_21_6_port, positive_inputs_21_5_port, 
      positive_inputs_21_4_port, positive_inputs_21_3_port, 
      positive_inputs_21_2_port, positive_inputs_21_1_port, 
      positive_inputs_20_63_port, positive_inputs_20_62_port, 
      positive_inputs_20_61_port, positive_inputs_20_60_port, 
      positive_inputs_20_59_port, positive_inputs_20_58_port, 
      positive_inputs_20_57_port, positive_inputs_20_56_port, 
      positive_inputs_20_55_port, positive_inputs_20_54_port, 
      positive_inputs_20_53_port, positive_inputs_20_52_port, 
      positive_inputs_20_51_port, positive_inputs_20_50_port, 
      positive_inputs_20_49_port, positive_inputs_20_48_port, 
      positive_inputs_20_47_port, positive_inputs_20_46_port, 
      positive_inputs_20_45_port, positive_inputs_20_44_port, 
      positive_inputs_20_43_port, positive_inputs_20_42_port, 
      positive_inputs_20_41_port, positive_inputs_20_40_port, 
      positive_inputs_20_39_port, positive_inputs_20_38_port, 
      positive_inputs_20_37_port, positive_inputs_20_36_port, 
      positive_inputs_20_35_port, positive_inputs_20_34_port, 
      positive_inputs_20_33_port, positive_inputs_20_32_port, 
      positive_inputs_20_31_port, positive_inputs_20_30_port, 
      positive_inputs_20_29_port, positive_inputs_20_28_port, 
      positive_inputs_20_27_port, positive_inputs_20_26_port, 
      positive_inputs_20_25_port, positive_inputs_20_24_port, 
      positive_inputs_20_23_port, positive_inputs_20_22_port, 
      positive_inputs_20_21_port, positive_inputs_20_20_port, 
      positive_inputs_20_19_port, positive_inputs_20_18_port, 
      positive_inputs_20_17_port, positive_inputs_20_16_port, 
      positive_inputs_20_15_port, positive_inputs_20_14_port, 
      positive_inputs_20_13_port, positive_inputs_20_12_port, 
      positive_inputs_20_11_port, positive_inputs_20_10_port, 
      positive_inputs_20_9_port, positive_inputs_20_8_port, 
      positive_inputs_20_7_port, positive_inputs_20_6_port, 
      positive_inputs_20_5_port, positive_inputs_20_4_port, 
      positive_inputs_20_3_port, positive_inputs_20_2_port, 
      positive_inputs_20_1_port, positive_inputs_19_63_port, 
      positive_inputs_19_62_port, positive_inputs_19_61_port, 
      positive_inputs_19_60_port, positive_inputs_19_59_port, 
      positive_inputs_19_58_port, positive_inputs_19_57_port, 
      positive_inputs_19_56_port, positive_inputs_19_55_port, 
      positive_inputs_19_54_port, positive_inputs_19_53_port, 
      positive_inputs_19_52_port, positive_inputs_19_51_port, 
      positive_inputs_19_50_port, positive_inputs_19_49_port, 
      positive_inputs_19_48_port, positive_inputs_19_47_port, 
      positive_inputs_19_46_port, positive_inputs_19_45_port, 
      positive_inputs_19_44_port, positive_inputs_19_43_port, 
      positive_inputs_19_42_port, positive_inputs_19_41_port, 
      positive_inputs_19_40_port, positive_inputs_19_39_port, 
      positive_inputs_19_38_port, positive_inputs_19_37_port, 
      positive_inputs_19_36_port, positive_inputs_19_35_port, 
      positive_inputs_19_34_port, positive_inputs_19_33_port, 
      positive_inputs_19_32_port, positive_inputs_19_31_port, 
      positive_inputs_19_30_port, positive_inputs_19_29_port, 
      positive_inputs_19_28_port, positive_inputs_19_27_port, 
      positive_inputs_19_26_port, positive_inputs_19_25_port, 
      positive_inputs_19_24_port, positive_inputs_19_23_port, 
      positive_inputs_19_22_port, positive_inputs_19_21_port, 
      positive_inputs_19_20_port, positive_inputs_19_19_port, 
      positive_inputs_19_18_port, positive_inputs_19_17_port, 
      positive_inputs_19_16_port, positive_inputs_19_15_port, 
      positive_inputs_19_14_port, positive_inputs_19_13_port, 
      positive_inputs_19_12_port, positive_inputs_19_11_port, 
      positive_inputs_19_10_port, positive_inputs_19_9_port, 
      positive_inputs_19_8_port, positive_inputs_19_7_port, 
      positive_inputs_19_6_port, positive_inputs_19_5_port, 
      positive_inputs_19_4_port, positive_inputs_19_3_port, 
      positive_inputs_19_2_port, positive_inputs_19_1_port, 
      positive_inputs_18_63_port, positive_inputs_18_62_port, 
      positive_inputs_18_61_port, positive_inputs_18_60_port, 
      positive_inputs_18_59_port, positive_inputs_18_58_port, 
      positive_inputs_18_57_port, positive_inputs_18_56_port, 
      positive_inputs_18_55_port, positive_inputs_18_54_port, 
      positive_inputs_18_53_port, positive_inputs_18_52_port, 
      positive_inputs_18_51_port, positive_inputs_18_50_port, 
      positive_inputs_18_49_port, positive_inputs_18_48_port, 
      positive_inputs_18_47_port, positive_inputs_18_46_port, 
      positive_inputs_18_45_port, positive_inputs_18_44_port, 
      positive_inputs_18_43_port, positive_inputs_18_42_port, 
      positive_inputs_18_41_port, positive_inputs_18_40_port, 
      positive_inputs_18_39_port, positive_inputs_18_38_port, 
      positive_inputs_18_37_port, positive_inputs_18_36_port, 
      positive_inputs_18_35_port, positive_inputs_18_34_port, 
      positive_inputs_18_33_port, positive_inputs_18_32_port, 
      positive_inputs_18_31_port, positive_inputs_18_30_port, 
      positive_inputs_18_29_port, positive_inputs_18_28_port, 
      positive_inputs_18_27_port, positive_inputs_18_26_port, 
      positive_inputs_18_25_port, positive_inputs_18_24_port, 
      positive_inputs_18_23_port, positive_inputs_18_22_port, 
      positive_inputs_18_21_port, positive_inputs_18_20_port, 
      positive_inputs_18_19_port, positive_inputs_18_18_port, 
      positive_inputs_18_17_port, positive_inputs_18_16_port, 
      positive_inputs_18_15_port, positive_inputs_18_14_port, 
      positive_inputs_18_13_port, positive_inputs_18_12_port, 
      positive_inputs_18_11_port, positive_inputs_18_10_port, 
      positive_inputs_18_9_port, positive_inputs_18_8_port, 
      positive_inputs_18_7_port, positive_inputs_18_6_port, 
      positive_inputs_18_5_port, positive_inputs_18_4_port, 
      positive_inputs_18_3_port, positive_inputs_18_2_port, 
      positive_inputs_18_1_port, positive_inputs_17_63_port, 
      positive_inputs_17_62_port, positive_inputs_17_61_port, 
      positive_inputs_17_60_port, positive_inputs_17_59_port, 
      positive_inputs_17_58_port, positive_inputs_17_57_port, 
      positive_inputs_17_56_port, positive_inputs_17_55_port, 
      positive_inputs_17_54_port, positive_inputs_17_53_port, 
      positive_inputs_17_52_port, positive_inputs_17_51_port, 
      positive_inputs_17_50_port, positive_inputs_17_49_port, 
      positive_inputs_17_48_port, positive_inputs_17_47_port, 
      positive_inputs_17_46_port, positive_inputs_17_45_port, 
      positive_inputs_17_44_port, positive_inputs_17_43_port, 
      positive_inputs_17_42_port, positive_inputs_17_41_port, 
      positive_inputs_17_40_port, positive_inputs_17_39_port, 
      positive_inputs_17_38_port, positive_inputs_17_37_port, 
      positive_inputs_17_36_port, positive_inputs_17_35_port, 
      positive_inputs_17_34_port, positive_inputs_17_33_port, 
      positive_inputs_17_32_port, positive_inputs_17_31_port, 
      positive_inputs_17_30_port, positive_inputs_17_29_port, 
      positive_inputs_17_28_port, positive_inputs_17_27_port, 
      positive_inputs_17_26_port, positive_inputs_17_25_port, 
      positive_inputs_17_24_port, positive_inputs_17_23_port, 
      positive_inputs_17_22_port, positive_inputs_17_21_port, 
      positive_inputs_17_20_port, positive_inputs_17_19_port, 
      positive_inputs_17_18_port, positive_inputs_17_17_port, 
      positive_inputs_17_16_port, positive_inputs_17_15_port, 
      positive_inputs_17_14_port, positive_inputs_17_13_port, 
      positive_inputs_17_12_port, positive_inputs_17_11_port, 
      positive_inputs_17_10_port, positive_inputs_17_9_port, 
      positive_inputs_17_8_port, positive_inputs_17_7_port, 
      positive_inputs_17_6_port, positive_inputs_17_5_port, 
      positive_inputs_17_4_port, positive_inputs_17_3_port, 
      positive_inputs_17_2_port, positive_inputs_17_1_port, 
      positive_inputs_31_63_port, positive_inputs_31_62_port, 
      positive_inputs_31_61_port, positive_inputs_31_60_port, 
      positive_inputs_31_59_port, positive_inputs_31_58_port, 
      positive_inputs_31_57_port, positive_inputs_31_56_port, 
      positive_inputs_31_55_port, positive_inputs_31_54_port, 
      positive_inputs_31_53_port, positive_inputs_31_52_port, 
      positive_inputs_31_51_port, positive_inputs_31_50_port, 
      positive_inputs_31_49_port, positive_inputs_31_48_port, 
      positive_inputs_31_47_port, positive_inputs_31_46_port, 
      positive_inputs_31_45_port, positive_inputs_31_44_port, 
      positive_inputs_31_43_port, positive_inputs_31_42_port, 
      positive_inputs_31_41_port, positive_inputs_31_40_port, 
      positive_inputs_31_39_port, positive_inputs_31_38_port, 
      positive_inputs_31_37_port, positive_inputs_31_36_port, 
      positive_inputs_31_35_port, positive_inputs_31_34_port, 
      positive_inputs_31_33_port, positive_inputs_31_32_port, 
      positive_inputs_31_31_port, positive_inputs_31_30_port, 
      positive_inputs_31_29_port, positive_inputs_31_28_port, 
      positive_inputs_31_27_port, positive_inputs_31_26_port, 
      positive_inputs_31_25_port, positive_inputs_31_24_port, 
      positive_inputs_31_23_port, positive_inputs_31_22_port, 
      positive_inputs_31_21_port, positive_inputs_31_20_port, 
      positive_inputs_31_19_port, positive_inputs_31_18_port, 
      positive_inputs_31_17_port, positive_inputs_31_16_port, 
      positive_inputs_31_15_port, positive_inputs_31_14_port, 
      positive_inputs_31_13_port, positive_inputs_31_12_port, 
      positive_inputs_31_11_port, positive_inputs_31_10_port, 
      positive_inputs_31_9_port, positive_inputs_31_8_port, 
      positive_inputs_31_7_port, positive_inputs_31_6_port, 
      positive_inputs_31_5_port, positive_inputs_31_4_port, 
      positive_inputs_31_3_port, positive_inputs_31_2_port, 
      positive_inputs_31_1_port, positive_inputs_30_63_port, 
      positive_inputs_30_62_port, positive_inputs_30_61_port, 
      positive_inputs_30_60_port, positive_inputs_30_59_port, 
      positive_inputs_30_58_port, positive_inputs_30_57_port, 
      positive_inputs_30_56_port, positive_inputs_30_55_port, 
      positive_inputs_30_54_port, positive_inputs_30_53_port, 
      positive_inputs_30_52_port, positive_inputs_30_51_port, 
      positive_inputs_30_50_port, positive_inputs_30_49_port, 
      positive_inputs_30_48_port, positive_inputs_30_47_port, 
      positive_inputs_30_46_port, positive_inputs_30_45_port, 
      positive_inputs_30_44_port, positive_inputs_30_43_port, 
      positive_inputs_30_42_port, positive_inputs_30_41_port, 
      positive_inputs_30_40_port, positive_inputs_30_39_port, 
      positive_inputs_30_38_port, positive_inputs_30_37_port, 
      positive_inputs_30_36_port, positive_inputs_30_35_port, 
      positive_inputs_30_34_port, positive_inputs_30_33_port, 
      positive_inputs_30_32_port, positive_inputs_30_31_port, 
      positive_inputs_30_30_port, positive_inputs_30_29_port, 
      positive_inputs_30_28_port, positive_inputs_30_27_port, 
      positive_inputs_30_26_port, positive_inputs_30_25_port, 
      positive_inputs_30_24_port, positive_inputs_30_23_port, 
      positive_inputs_30_22_port, positive_inputs_30_21_port, 
      positive_inputs_30_20_port, positive_inputs_30_19_port, 
      positive_inputs_30_18_port, positive_inputs_30_17_port, 
      positive_inputs_30_16_port, positive_inputs_30_15_port, 
      positive_inputs_30_14_port, positive_inputs_30_13_port, 
      positive_inputs_30_12_port, positive_inputs_30_11_port, 
      positive_inputs_30_10_port, positive_inputs_30_9_port, 
      positive_inputs_30_8_port, positive_inputs_30_7_port, 
      positive_inputs_30_6_port, positive_inputs_30_5_port, 
      positive_inputs_30_4_port, positive_inputs_30_3_port, 
      positive_inputs_30_2_port, positive_inputs_30_1_port, 
      positive_inputs_29_63_port, positive_inputs_29_62_port, 
      positive_inputs_29_61_port, positive_inputs_29_60_port, 
      positive_inputs_29_59_port, positive_inputs_29_58_port, 
      positive_inputs_29_57_port, positive_inputs_29_56_port, 
      positive_inputs_29_55_port, positive_inputs_29_54_port, 
      positive_inputs_29_53_port, positive_inputs_29_52_port, 
      positive_inputs_29_51_port, positive_inputs_29_50_port, 
      positive_inputs_29_49_port, positive_inputs_29_48_port, 
      positive_inputs_29_47_port, positive_inputs_29_46_port, 
      positive_inputs_29_45_port, positive_inputs_29_44_port, 
      positive_inputs_29_43_port, positive_inputs_29_42_port, 
      positive_inputs_29_41_port, positive_inputs_29_40_port, 
      positive_inputs_29_39_port, positive_inputs_29_38_port, 
      positive_inputs_29_37_port, positive_inputs_29_36_port, 
      positive_inputs_29_35_port, positive_inputs_29_34_port, 
      positive_inputs_29_33_port, positive_inputs_29_32_port, 
      positive_inputs_29_31_port, positive_inputs_29_30_port, 
      positive_inputs_29_29_port, positive_inputs_29_28_port, 
      positive_inputs_29_27_port, positive_inputs_29_26_port, 
      positive_inputs_29_25_port, positive_inputs_29_24_port, 
      positive_inputs_29_23_port, positive_inputs_29_22_port, 
      positive_inputs_29_21_port, positive_inputs_29_20_port, 
      positive_inputs_29_19_port, positive_inputs_29_18_port, 
      positive_inputs_29_17_port, positive_inputs_29_16_port, 
      positive_inputs_29_15_port, positive_inputs_29_14_port, 
      positive_inputs_29_13_port, positive_inputs_29_12_port, 
      positive_inputs_29_11_port, positive_inputs_29_10_port, 
      positive_inputs_29_9_port, positive_inputs_29_8_port, 
      positive_inputs_29_7_port, positive_inputs_29_6_port, 
      positive_inputs_29_5_port, positive_inputs_29_4_port, 
      positive_inputs_29_3_port, positive_inputs_29_2_port, 
      positive_inputs_29_1_port, positive_inputs_28_63_port, 
      positive_inputs_28_62_port, positive_inputs_28_61_port, 
      positive_inputs_28_60_port, positive_inputs_28_59_port, 
      positive_inputs_28_58_port, positive_inputs_28_57_port, 
      positive_inputs_28_56_port, positive_inputs_28_55_port, 
      positive_inputs_28_54_port, positive_inputs_28_53_port, 
      positive_inputs_28_52_port, positive_inputs_28_51_port, 
      positive_inputs_28_50_port, positive_inputs_28_49_port, 
      positive_inputs_28_48_port, positive_inputs_28_47_port, 
      positive_inputs_28_46_port, positive_inputs_28_45_port, 
      positive_inputs_28_44_port, positive_inputs_28_43_port, 
      positive_inputs_28_42_port, positive_inputs_28_41_port, 
      positive_inputs_28_40_port, positive_inputs_28_39_port, 
      positive_inputs_28_38_port, positive_inputs_28_37_port, 
      positive_inputs_28_36_port, positive_inputs_28_35_port, 
      positive_inputs_28_34_port, positive_inputs_28_33_port, 
      positive_inputs_28_32_port, positive_inputs_28_31_port, 
      positive_inputs_28_30_port, positive_inputs_28_29_port, 
      positive_inputs_28_28_port, positive_inputs_28_27_port, 
      positive_inputs_28_26_port, positive_inputs_28_25_port, 
      positive_inputs_28_24_port, positive_inputs_28_23_port, 
      positive_inputs_28_22_port, positive_inputs_28_21_port, 
      positive_inputs_28_20_port, positive_inputs_28_19_port, 
      positive_inputs_28_18_port, positive_inputs_28_17_port, 
      positive_inputs_28_16_port, positive_inputs_28_15_port, 
      positive_inputs_28_14_port, positive_inputs_28_13_port, 
      positive_inputs_28_12_port, positive_inputs_28_11_port, 
      positive_inputs_28_10_port, positive_inputs_28_9_port, 
      positive_inputs_28_8_port, positive_inputs_28_7_port, 
      positive_inputs_28_6_port, positive_inputs_28_5_port, 
      positive_inputs_28_4_port, positive_inputs_28_3_port, 
      positive_inputs_28_2_port, positive_inputs_28_1_port, 
      positive_inputs_27_63_port, positive_inputs_27_62_port, 
      positive_inputs_27_61_port, positive_inputs_27_60_port, 
      positive_inputs_27_59_port, positive_inputs_27_58_port, 
      positive_inputs_27_57_port, positive_inputs_27_56_port, 
      positive_inputs_27_55_port, positive_inputs_27_54_port, 
      positive_inputs_27_53_port, positive_inputs_27_52_port, 
      positive_inputs_27_51_port, positive_inputs_27_50_port, 
      positive_inputs_27_49_port, positive_inputs_27_48_port, 
      positive_inputs_27_47_port, positive_inputs_27_46_port, 
      positive_inputs_27_45_port, positive_inputs_27_44_port, 
      positive_inputs_27_43_port, positive_inputs_27_42_port, 
      positive_inputs_27_41_port, positive_inputs_27_40_port, 
      positive_inputs_27_39_port, positive_inputs_27_38_port, 
      positive_inputs_27_37_port, positive_inputs_27_36_port, 
      positive_inputs_27_35_port, positive_inputs_27_34_port, 
      positive_inputs_27_33_port, positive_inputs_27_32_port, 
      positive_inputs_27_31_port, positive_inputs_27_30_port, 
      positive_inputs_27_29_port, positive_inputs_27_28_port, 
      positive_inputs_27_27_port, positive_inputs_27_26_port, 
      positive_inputs_27_25_port, positive_inputs_27_24_port, 
      positive_inputs_27_23_port, positive_inputs_27_22_port, 
      positive_inputs_27_21_port, positive_inputs_27_20_port, 
      positive_inputs_27_19_port, positive_inputs_27_18_port, 
      positive_inputs_27_17_port, positive_inputs_27_16_port, 
      positive_inputs_27_15_port, positive_inputs_27_14_port, 
      positive_inputs_27_13_port, positive_inputs_27_12_port, 
      positive_inputs_27_11_port, positive_inputs_27_10_port, 
      positive_inputs_27_9_port, positive_inputs_27_8_port, 
      positive_inputs_27_7_port, positive_inputs_27_6_port, 
      positive_inputs_27_5_port, positive_inputs_27_4_port, 
      positive_inputs_27_3_port, positive_inputs_27_2_port, 
      positive_inputs_27_1_port, positive_inputs_26_63_port, 
      positive_inputs_26_62_port, positive_inputs_26_61_port, 
      positive_inputs_26_60_port, positive_inputs_26_59_port, 
      positive_inputs_26_58_port, positive_inputs_26_57_port, 
      positive_inputs_26_56_port, positive_inputs_26_55_port, 
      positive_inputs_26_54_port, positive_inputs_26_53_port, 
      positive_inputs_26_52_port, positive_inputs_26_51_port, 
      positive_inputs_26_50_port, positive_inputs_26_49_port, 
      positive_inputs_26_48_port, positive_inputs_26_47_port, 
      positive_inputs_26_46_port, positive_inputs_26_45_port, 
      positive_inputs_26_44_port, positive_inputs_26_43_port, 
      positive_inputs_26_42_port, positive_inputs_26_41_port, 
      positive_inputs_26_40_port, positive_inputs_26_39_port, 
      positive_inputs_26_38_port, positive_inputs_26_37_port, 
      positive_inputs_26_36_port, positive_inputs_26_35_port, 
      positive_inputs_26_34_port, positive_inputs_26_33_port, 
      positive_inputs_26_32_port, positive_inputs_26_31_port, 
      positive_inputs_26_30_port, positive_inputs_26_29_port, 
      positive_inputs_26_28_port, positive_inputs_26_27_port, 
      positive_inputs_26_26_port, positive_inputs_26_25_port, 
      positive_inputs_26_24_port, positive_inputs_26_23_port, 
      positive_inputs_26_22_port, positive_inputs_26_21_port, 
      positive_inputs_26_20_port, positive_inputs_26_19_port, 
      positive_inputs_26_18_port, positive_inputs_26_17_port, 
      positive_inputs_26_16_port, positive_inputs_26_15_port, 
      positive_inputs_26_14_port, positive_inputs_26_13_port, 
      positive_inputs_26_12_port, positive_inputs_26_11_port, 
      positive_inputs_26_10_port, positive_inputs_26_9_port, 
      positive_inputs_26_8_port, positive_inputs_26_7_port, 
      positive_inputs_26_6_port, positive_inputs_26_5_port, 
      positive_inputs_26_4_port, positive_inputs_26_3_port, 
      positive_inputs_26_2_port, positive_inputs_26_1_port, 
      positive_inputs_25_63_port, positive_inputs_25_62_port, 
      positive_inputs_25_61_port, positive_inputs_25_60_port, 
      positive_inputs_25_59_port, positive_inputs_25_58_port, 
      positive_inputs_25_57_port, positive_inputs_25_56_port, 
      positive_inputs_25_55_port, positive_inputs_25_54_port, 
      positive_inputs_25_53_port, positive_inputs_25_52_port, 
      positive_inputs_25_51_port, positive_inputs_25_50_port, 
      positive_inputs_25_49_port, positive_inputs_25_48_port, 
      positive_inputs_25_47_port, positive_inputs_25_46_port, 
      positive_inputs_25_45_port, positive_inputs_25_44_port, 
      positive_inputs_25_43_port, positive_inputs_25_42_port, 
      positive_inputs_25_41_port, positive_inputs_25_40_port, 
      positive_inputs_25_39_port, positive_inputs_25_38_port, 
      positive_inputs_25_37_port, positive_inputs_25_36_port, 
      positive_inputs_25_35_port, positive_inputs_25_34_port, 
      positive_inputs_25_33_port, positive_inputs_25_32_port, 
      positive_inputs_25_31_port, positive_inputs_25_30_port, 
      positive_inputs_25_29_port, positive_inputs_25_28_port, 
      positive_inputs_25_27_port, positive_inputs_25_26_port, 
      positive_inputs_25_25_port, positive_inputs_25_24_port, 
      positive_inputs_25_23_port, positive_inputs_25_22_port, 
      positive_inputs_25_21_port, positive_inputs_25_20_port, 
      positive_inputs_25_19_port, positive_inputs_25_18_port, 
      positive_inputs_25_17_port, positive_inputs_25_16_port, 
      positive_inputs_25_15_port, positive_inputs_25_14_port, 
      positive_inputs_25_13_port, positive_inputs_25_12_port, 
      positive_inputs_25_11_port, positive_inputs_25_10_port, 
      positive_inputs_25_9_port, positive_inputs_25_8_port, 
      positive_inputs_25_7_port, positive_inputs_25_6_port, 
      positive_inputs_25_5_port, positive_inputs_25_4_port, 
      positive_inputs_25_3_port, positive_inputs_25_2_port, 
      positive_inputs_25_1_port, negative_inputs_8_63_port, 
      negative_inputs_8_62_port, negative_inputs_8_61_port, 
      negative_inputs_8_60_port, negative_inputs_8_59_port, 
      negative_inputs_8_58_port, negative_inputs_8_57_port, 
      negative_inputs_8_56_port, negative_inputs_8_55_port, 
      negative_inputs_8_54_port, negative_inputs_8_53_port, 
      negative_inputs_8_52_port, negative_inputs_8_51_port, 
      negative_inputs_8_50_port, negative_inputs_8_49_port, 
      negative_inputs_8_48_port, negative_inputs_8_47_port, 
      negative_inputs_8_46_port, negative_inputs_8_45_port, 
      negative_inputs_8_44_port, negative_inputs_8_43_port, 
      negative_inputs_8_42_port, negative_inputs_8_41_port, 
      negative_inputs_8_40_port, negative_inputs_8_39_port, 
      negative_inputs_8_38_port, negative_inputs_8_37_port, 
      negative_inputs_8_36_port, negative_inputs_8_35_port, 
      negative_inputs_8_34_port, negative_inputs_8_33_port, 
      negative_inputs_8_32_port, negative_inputs_8_31_port, 
      negative_inputs_8_30_port, negative_inputs_8_29_port, 
      negative_inputs_8_28_port, negative_inputs_8_27_port, 
      negative_inputs_8_26_port, negative_inputs_8_25_port, 
      negative_inputs_8_24_port, negative_inputs_8_23_port, 
      negative_inputs_8_22_port, negative_inputs_8_21_port, 
      negative_inputs_8_20_port, negative_inputs_8_19_port, 
      negative_inputs_8_18_port, negative_inputs_8_17_port, 
      negative_inputs_8_16_port, negative_inputs_8_15_port, 
      negative_inputs_8_14_port, negative_inputs_8_13_port, 
      negative_inputs_8_12_port, negative_inputs_8_11_port, 
      negative_inputs_8_10_port, negative_inputs_8_9_port, 
      negative_inputs_8_8_port, negative_inputs_8_7_port, 
      negative_inputs_8_6_port, negative_inputs_8_5_port, 
      negative_inputs_8_4_port, negative_inputs_8_3_port, 
      negative_inputs_8_2_port, negative_inputs_8_1_port, 
      negative_inputs_7_63_port, negative_inputs_7_62_port, 
      negative_inputs_7_61_port, negative_inputs_7_60_port, 
      negative_inputs_7_59_port, negative_inputs_7_58_port, 
      negative_inputs_7_57_port, negative_inputs_7_56_port, 
      negative_inputs_7_55_port, negative_inputs_7_54_port, 
      negative_inputs_7_53_port, negative_inputs_7_52_port, 
      negative_inputs_7_51_port, negative_inputs_7_50_port, 
      negative_inputs_7_49_port, negative_inputs_7_48_port, 
      negative_inputs_7_47_port, negative_inputs_7_46_port, 
      negative_inputs_7_45_port, negative_inputs_7_44_port, 
      negative_inputs_7_43_port, negative_inputs_7_42_port, 
      negative_inputs_7_41_port, negative_inputs_7_40_port, 
      negative_inputs_7_39_port, negative_inputs_7_38_port, 
      negative_inputs_7_37_port, negative_inputs_7_36_port, 
      negative_inputs_7_35_port, negative_inputs_7_34_port, 
      negative_inputs_7_33_port, negative_inputs_7_32_port, 
      negative_inputs_7_31_port, negative_inputs_7_30_port, 
      negative_inputs_7_29_port, negative_inputs_7_28_port, 
      negative_inputs_7_27_port, negative_inputs_7_26_port, 
      negative_inputs_7_25_port, negative_inputs_7_24_port, 
      negative_inputs_7_23_port, negative_inputs_7_22_port, 
      negative_inputs_7_21_port, negative_inputs_7_20_port, 
      negative_inputs_7_19_port, negative_inputs_7_18_port, 
      negative_inputs_7_17_port, negative_inputs_7_16_port, 
      negative_inputs_7_15_port, negative_inputs_7_14_port, 
      negative_inputs_7_13_port, negative_inputs_7_12_port, 
      negative_inputs_7_11_port, negative_inputs_7_10_port, 
      negative_inputs_7_9_port, negative_inputs_7_8_port, 
      negative_inputs_7_7_port, negative_inputs_7_6_port, 
      negative_inputs_7_5_port, negative_inputs_7_4_port, 
      negative_inputs_7_3_port, negative_inputs_7_2_port, 
      negative_inputs_7_1_port, negative_inputs_6_63_port, 
      negative_inputs_6_62_port, negative_inputs_6_61_port, 
      negative_inputs_6_60_port, negative_inputs_6_59_port, 
      negative_inputs_6_58_port, negative_inputs_6_57_port, 
      negative_inputs_6_56_port, negative_inputs_6_55_port, 
      negative_inputs_6_54_port, negative_inputs_6_53_port, 
      negative_inputs_6_52_port, negative_inputs_6_51_port, 
      negative_inputs_6_50_port, negative_inputs_6_49_port, 
      negative_inputs_6_48_port, negative_inputs_6_47_port, 
      negative_inputs_6_46_port, negative_inputs_6_45_port, 
      negative_inputs_6_44_port, negative_inputs_6_43_port, 
      negative_inputs_6_42_port, negative_inputs_6_41_port, 
      negative_inputs_6_40_port, negative_inputs_6_39_port, 
      negative_inputs_6_38_port, negative_inputs_6_37_port, 
      negative_inputs_6_36_port, negative_inputs_6_35_port, 
      negative_inputs_6_34_port, negative_inputs_6_33_port, 
      negative_inputs_6_32_port, negative_inputs_6_31_port, 
      negative_inputs_6_30_port, negative_inputs_6_29_port, 
      negative_inputs_6_28_port, negative_inputs_6_27_port, 
      negative_inputs_6_26_port, negative_inputs_6_25_port, 
      negative_inputs_6_24_port, negative_inputs_6_23_port, 
      negative_inputs_6_22_port, negative_inputs_6_21_port, 
      negative_inputs_6_20_port, negative_inputs_6_19_port, 
      negative_inputs_6_18_port, negative_inputs_6_17_port, 
      negative_inputs_6_16_port, negative_inputs_6_15_port, 
      negative_inputs_6_14_port, negative_inputs_6_13_port, 
      negative_inputs_6_12_port, negative_inputs_6_11_port, 
      negative_inputs_6_10_port, negative_inputs_6_9_port, 
      negative_inputs_6_8_port, negative_inputs_6_7_port, 
      negative_inputs_6_6_port, negative_inputs_6_5_port, 
      negative_inputs_6_4_port, negative_inputs_6_3_port, 
      negative_inputs_6_2_port, negative_inputs_6_1_port, 
      negative_inputs_5_63_port, negative_inputs_5_62_port, 
      negative_inputs_5_61_port, negative_inputs_5_60_port, 
      negative_inputs_5_59_port, negative_inputs_5_58_port, 
      negative_inputs_5_57_port, negative_inputs_5_56_port, 
      negative_inputs_5_55_port, negative_inputs_5_54_port, 
      negative_inputs_5_53_port, negative_inputs_5_52_port, 
      negative_inputs_5_51_port, negative_inputs_5_50_port, 
      negative_inputs_5_49_port, negative_inputs_5_48_port, 
      negative_inputs_5_47_port, negative_inputs_5_46_port, 
      negative_inputs_5_45_port, negative_inputs_5_44_port, 
      negative_inputs_5_43_port, negative_inputs_5_42_port, 
      negative_inputs_5_41_port, negative_inputs_5_40_port, 
      negative_inputs_5_39_port, negative_inputs_5_38_port, 
      negative_inputs_5_37_port, negative_inputs_5_36_port, 
      negative_inputs_5_35_port, negative_inputs_5_34_port, 
      negative_inputs_5_33_port, negative_inputs_5_32_port, 
      negative_inputs_5_31_port, negative_inputs_5_30_port, 
      negative_inputs_5_29_port, negative_inputs_5_28_port, 
      negative_inputs_5_27_port, negative_inputs_5_26_port, 
      negative_inputs_5_25_port, negative_inputs_5_24_port, 
      negative_inputs_5_23_port, negative_inputs_5_22_port, 
      negative_inputs_5_21_port, negative_inputs_5_20_port, 
      negative_inputs_5_19_port, negative_inputs_5_18_port, 
      negative_inputs_5_17_port, negative_inputs_5_16_port, 
      negative_inputs_5_15_port, negative_inputs_5_14_port, 
      negative_inputs_5_13_port, negative_inputs_5_12_port, 
      negative_inputs_5_11_port, negative_inputs_5_10_port, 
      negative_inputs_5_9_port, negative_inputs_5_8_port, 
      negative_inputs_5_7_port, negative_inputs_5_6_port, 
      negative_inputs_5_5_port, negative_inputs_5_4_port, 
      negative_inputs_5_3_port, negative_inputs_5_2_port, 
      negative_inputs_5_1_port, negative_inputs_4_63_port, 
      negative_inputs_4_62_port, negative_inputs_4_61_port, 
      negative_inputs_4_60_port, negative_inputs_4_59_port, 
      negative_inputs_4_58_port, negative_inputs_4_57_port, 
      negative_inputs_4_56_port, negative_inputs_4_55_port, 
      negative_inputs_4_54_port, negative_inputs_4_53_port, 
      negative_inputs_4_52_port, negative_inputs_4_51_port, 
      negative_inputs_4_50_port, negative_inputs_4_49_port, 
      negative_inputs_4_48_port, negative_inputs_4_47_port, 
      negative_inputs_4_46_port, negative_inputs_4_45_port, 
      negative_inputs_4_44_port, negative_inputs_4_43_port, 
      negative_inputs_4_42_port, negative_inputs_4_41_port, 
      negative_inputs_4_40_port, negative_inputs_4_39_port, 
      negative_inputs_4_38_port, negative_inputs_4_37_port, 
      negative_inputs_4_36_port, negative_inputs_4_35_port, 
      negative_inputs_4_34_port, negative_inputs_4_33_port, 
      negative_inputs_4_32_port, negative_inputs_4_31_port, 
      negative_inputs_4_30_port, negative_inputs_4_29_port, 
      negative_inputs_4_28_port, negative_inputs_4_27_port, 
      negative_inputs_4_26_port, negative_inputs_4_25_port, 
      negative_inputs_4_24_port, negative_inputs_4_23_port, 
      negative_inputs_4_22_port, negative_inputs_4_21_port, 
      negative_inputs_4_20_port, negative_inputs_4_19_port, 
      negative_inputs_4_18_port, negative_inputs_4_17_port, 
      negative_inputs_4_16_port, negative_inputs_4_15_port, 
      negative_inputs_4_14_port, negative_inputs_4_13_port, 
      negative_inputs_4_12_port, negative_inputs_4_11_port, 
      negative_inputs_4_10_port, negative_inputs_4_9_port, 
      negative_inputs_4_8_port, negative_inputs_4_7_port, 
      negative_inputs_4_6_port, negative_inputs_4_5_port, 
      negative_inputs_4_4_port, negative_inputs_4_3_port, 
      negative_inputs_4_2_port, negative_inputs_4_1_port, 
      negative_inputs_3_63_port, negative_inputs_3_62_port, 
      negative_inputs_3_61_port, negative_inputs_3_60_port, 
      negative_inputs_3_59_port, negative_inputs_3_58_port, 
      negative_inputs_3_57_port, negative_inputs_3_56_port, 
      negative_inputs_3_55_port, negative_inputs_3_54_port, 
      negative_inputs_3_53_port, negative_inputs_3_52_port, 
      negative_inputs_3_51_port, negative_inputs_3_50_port, 
      negative_inputs_3_49_port, negative_inputs_3_48_port, 
      negative_inputs_3_47_port, negative_inputs_3_46_port, 
      negative_inputs_3_45_port, negative_inputs_3_44_port, 
      negative_inputs_3_43_port, negative_inputs_3_42_port, 
      negative_inputs_3_41_port, negative_inputs_3_40_port, 
      negative_inputs_3_39_port, negative_inputs_3_38_port, 
      negative_inputs_3_37_port, negative_inputs_3_36_port, 
      negative_inputs_3_35_port, negative_inputs_3_34_port, 
      negative_inputs_3_33_port, negative_inputs_3_32_port, 
      negative_inputs_3_31_port, negative_inputs_3_30_port, 
      negative_inputs_3_29_port, negative_inputs_3_28_port, 
      negative_inputs_3_27_port, negative_inputs_3_26_port, 
      negative_inputs_3_25_port, negative_inputs_3_24_port, 
      negative_inputs_3_23_port, negative_inputs_3_22_port, 
      negative_inputs_3_21_port, negative_inputs_3_20_port, 
      negative_inputs_3_19_port, negative_inputs_3_18_port, 
      negative_inputs_3_17_port, negative_inputs_3_16_port, 
      negative_inputs_3_15_port, negative_inputs_3_14_port, 
      negative_inputs_3_13_port, negative_inputs_3_12_port, 
      negative_inputs_3_11_port, negative_inputs_3_10_port, 
      negative_inputs_3_9_port, negative_inputs_3_8_port, 
      negative_inputs_3_7_port, negative_inputs_3_6_port, 
      negative_inputs_3_5_port, negative_inputs_3_4_port, 
      negative_inputs_3_3_port, negative_inputs_3_2_port, 
      negative_inputs_3_1_port, negative_inputs_2_63_port, 
      negative_inputs_2_62_port, negative_inputs_2_61_port, 
      negative_inputs_2_60_port, negative_inputs_2_59_port, 
      negative_inputs_2_58_port, negative_inputs_2_57_port, 
      negative_inputs_2_56_port, negative_inputs_2_55_port, 
      negative_inputs_2_54_port, negative_inputs_2_53_port, 
      negative_inputs_2_52_port, negative_inputs_2_51_port, 
      negative_inputs_2_50_port, negative_inputs_2_49_port, 
      negative_inputs_2_48_port, negative_inputs_2_47_port, 
      negative_inputs_2_46_port, negative_inputs_2_45_port, 
      negative_inputs_2_44_port, negative_inputs_2_43_port, 
      negative_inputs_2_42_port, negative_inputs_2_41_port, 
      negative_inputs_2_40_port, negative_inputs_2_39_port, 
      negative_inputs_2_38_port, negative_inputs_2_37_port, 
      negative_inputs_2_36_port, negative_inputs_2_35_port, 
      negative_inputs_2_34_port, negative_inputs_2_33_port, 
      negative_inputs_2_32_port, negative_inputs_2_31_port, 
      negative_inputs_2_30_port, negative_inputs_2_29_port, 
      negative_inputs_2_28_port, negative_inputs_2_27_port, 
      negative_inputs_2_26_port, negative_inputs_2_25_port, 
      negative_inputs_2_24_port, negative_inputs_2_23_port, 
      negative_inputs_2_22_port, negative_inputs_2_21_port, 
      negative_inputs_2_20_port, negative_inputs_2_19_port, 
      negative_inputs_2_18_port, negative_inputs_2_17_port, 
      negative_inputs_2_16_port, negative_inputs_2_15_port, 
      negative_inputs_2_14_port, negative_inputs_2_13_port, 
      negative_inputs_2_12_port, negative_inputs_2_11_port, 
      negative_inputs_2_10_port, negative_inputs_2_9_port, 
      negative_inputs_2_8_port, negative_inputs_2_7_port, 
      negative_inputs_2_6_port, negative_inputs_2_5_port, 
      negative_inputs_2_4_port, negative_inputs_2_3_port, 
      negative_inputs_2_2_port, negative_inputs_2_1_port, 
      negative_inputs_1_63_port, negative_inputs_1_62_port, 
      negative_inputs_1_61_port, negative_inputs_1_60_port, 
      negative_inputs_1_59_port, negative_inputs_1_58_port, 
      negative_inputs_1_57_port, negative_inputs_1_56_port, 
      negative_inputs_1_55_port, negative_inputs_1_54_port, 
      negative_inputs_1_53_port, negative_inputs_1_52_port, 
      negative_inputs_1_51_port, negative_inputs_1_50_port, 
      negative_inputs_1_49_port, negative_inputs_1_48_port, 
      negative_inputs_1_47_port, negative_inputs_1_46_port, 
      negative_inputs_1_45_port, negative_inputs_1_44_port, 
      negative_inputs_1_43_port, negative_inputs_1_42_port, 
      negative_inputs_1_41_port, negative_inputs_1_40_port, 
      negative_inputs_1_39_port, negative_inputs_1_38_port, 
      negative_inputs_1_37_port, negative_inputs_1_36_port, 
      negative_inputs_1_35_port, negative_inputs_1_34_port, 
      negative_inputs_1_33_port, negative_inputs_1_32_port, 
      negative_inputs_1_31_port, negative_inputs_1_30_port, 
      negative_inputs_1_29_port, negative_inputs_1_28_port, 
      negative_inputs_1_27_port, negative_inputs_1_26_port, 
      negative_inputs_1_25_port, negative_inputs_1_24_port, 
      negative_inputs_1_23_port, negative_inputs_1_22_port, 
      negative_inputs_1_21_port, negative_inputs_1_20_port, 
      negative_inputs_1_19_port, negative_inputs_1_18_port, 
      negative_inputs_1_17_port, negative_inputs_1_16_port, 
      negative_inputs_1_15_port, negative_inputs_1_14_port, 
      negative_inputs_1_13_port, negative_inputs_1_12_port, 
      negative_inputs_1_11_port, negative_inputs_1_10_port, 
      negative_inputs_1_9_port, negative_inputs_1_8_port, 
      negative_inputs_1_7_port, negative_inputs_1_6_port, 
      negative_inputs_1_5_port, negative_inputs_1_4_port, 
      negative_inputs_1_3_port, negative_inputs_1_2_port, 
      negative_inputs_1_1_port, negative_inputs_16_63_port, 
      negative_inputs_16_62_port, negative_inputs_16_61_port, 
      negative_inputs_16_60_port, negative_inputs_16_59_port, 
      negative_inputs_16_58_port, negative_inputs_16_57_port, 
      negative_inputs_16_56_port, negative_inputs_16_55_port, 
      negative_inputs_16_54_port, negative_inputs_16_53_port, 
      negative_inputs_16_52_port, negative_inputs_16_51_port, 
      negative_inputs_16_50_port, negative_inputs_16_49_port, 
      negative_inputs_16_48_port, negative_inputs_16_47_port, 
      negative_inputs_16_46_port, negative_inputs_16_45_port, 
      negative_inputs_16_44_port, negative_inputs_16_43_port, 
      negative_inputs_16_42_port, negative_inputs_16_41_port, 
      negative_inputs_16_40_port, negative_inputs_16_39_port, 
      negative_inputs_16_38_port, negative_inputs_16_37_port, 
      negative_inputs_16_36_port, negative_inputs_16_35_port, 
      negative_inputs_16_34_port, negative_inputs_16_33_port, 
      negative_inputs_16_32_port, negative_inputs_16_31_port, 
      negative_inputs_16_30_port, negative_inputs_16_29_port, 
      negative_inputs_16_28_port, negative_inputs_16_27_port, 
      negative_inputs_16_26_port, negative_inputs_16_25_port, 
      negative_inputs_16_24_port, negative_inputs_16_23_port, 
      negative_inputs_16_22_port, negative_inputs_16_21_port, 
      negative_inputs_16_20_port, negative_inputs_16_19_port, 
      negative_inputs_16_18_port, negative_inputs_16_17_port, 
      negative_inputs_16_16_port, negative_inputs_16_15_port, 
      negative_inputs_16_14_port, negative_inputs_16_13_port, 
      negative_inputs_16_12_port, negative_inputs_16_11_port, 
      negative_inputs_16_10_port, negative_inputs_16_9_port, 
      negative_inputs_16_8_port, negative_inputs_16_7_port, 
      negative_inputs_16_6_port, negative_inputs_16_5_port, 
      negative_inputs_16_4_port, negative_inputs_16_3_port, 
      negative_inputs_16_2_port, negative_inputs_16_1_port, 
      negative_inputs_15_63_port, negative_inputs_15_62_port, 
      negative_inputs_15_61_port, negative_inputs_15_60_port, 
      negative_inputs_15_59_port, negative_inputs_15_58_port, 
      negative_inputs_15_57_port, negative_inputs_15_56_port, 
      negative_inputs_15_55_port, negative_inputs_15_54_port, 
      negative_inputs_15_53_port, negative_inputs_15_52_port, 
      negative_inputs_15_51_port, negative_inputs_15_50_port, 
      negative_inputs_15_49_port, negative_inputs_15_48_port, 
      negative_inputs_15_47_port, negative_inputs_15_46_port, 
      negative_inputs_15_45_port, negative_inputs_15_44_port, 
      negative_inputs_15_43_port, negative_inputs_15_42_port, 
      negative_inputs_15_41_port, negative_inputs_15_40_port, 
      negative_inputs_15_39_port, negative_inputs_15_38_port, 
      negative_inputs_15_37_port, negative_inputs_15_36_port, 
      negative_inputs_15_35_port, negative_inputs_15_34_port, 
      negative_inputs_15_33_port, negative_inputs_15_32_port, 
      negative_inputs_15_31_port, negative_inputs_15_30_port, 
      negative_inputs_15_29_port, negative_inputs_15_28_port, 
      negative_inputs_15_27_port, negative_inputs_15_26_port, 
      negative_inputs_15_25_port, negative_inputs_15_24_port, 
      negative_inputs_15_23_port, negative_inputs_15_22_port, 
      negative_inputs_15_21_port, negative_inputs_15_20_port, 
      negative_inputs_15_19_port, negative_inputs_15_18_port, 
      negative_inputs_15_17_port, negative_inputs_15_16_port, 
      negative_inputs_15_15_port, negative_inputs_15_14_port, 
      negative_inputs_15_13_port, negative_inputs_15_12_port, 
      negative_inputs_15_11_port, negative_inputs_15_10_port, 
      negative_inputs_15_9_port, negative_inputs_15_8_port, 
      negative_inputs_15_7_port, negative_inputs_15_6_port, 
      negative_inputs_15_5_port, negative_inputs_15_4_port, 
      negative_inputs_15_3_port, negative_inputs_15_2_port, 
      negative_inputs_15_1_port, negative_inputs_14_63_port, 
      negative_inputs_14_62_port, negative_inputs_14_61_port, 
      negative_inputs_14_60_port, negative_inputs_14_59_port, 
      negative_inputs_14_58_port, negative_inputs_14_57_port, 
      negative_inputs_14_56_port, negative_inputs_14_55_port, 
      negative_inputs_14_54_port, negative_inputs_14_53_port, 
      negative_inputs_14_52_port, negative_inputs_14_51_port, 
      negative_inputs_14_50_port, negative_inputs_14_49_port, 
      negative_inputs_14_48_port, negative_inputs_14_47_port, 
      negative_inputs_14_46_port, negative_inputs_14_45_port, 
      negative_inputs_14_44_port, negative_inputs_14_43_port, 
      negative_inputs_14_42_port, negative_inputs_14_41_port, 
      negative_inputs_14_40_port, negative_inputs_14_39_port, 
      negative_inputs_14_38_port, negative_inputs_14_37_port, 
      negative_inputs_14_36_port, negative_inputs_14_35_port, 
      negative_inputs_14_34_port, negative_inputs_14_33_port, 
      negative_inputs_14_32_port, negative_inputs_14_31_port, 
      negative_inputs_14_30_port, negative_inputs_14_29_port, 
      negative_inputs_14_28_port, negative_inputs_14_27_port, 
      negative_inputs_14_26_port, negative_inputs_14_25_port, 
      negative_inputs_14_24_port, negative_inputs_14_23_port, 
      negative_inputs_14_22_port, negative_inputs_14_21_port, 
      negative_inputs_14_20_port, negative_inputs_14_19_port, 
      negative_inputs_14_18_port, negative_inputs_14_17_port, 
      negative_inputs_14_16_port, negative_inputs_14_15_port, 
      negative_inputs_14_14_port, negative_inputs_14_13_port, 
      negative_inputs_14_12_port, negative_inputs_14_11_port, 
      negative_inputs_14_10_port, negative_inputs_14_9_port, 
      negative_inputs_14_8_port, negative_inputs_14_7_port, 
      negative_inputs_14_6_port, negative_inputs_14_5_port, 
      negative_inputs_14_4_port, negative_inputs_14_3_port, 
      negative_inputs_14_2_port, negative_inputs_14_1_port, 
      negative_inputs_13_63_port, negative_inputs_13_62_port, 
      negative_inputs_13_61_port, negative_inputs_13_60_port, 
      negative_inputs_13_59_port, negative_inputs_13_58_port, 
      negative_inputs_13_57_port, negative_inputs_13_56_port, 
      negative_inputs_13_55_port, negative_inputs_13_54_port, 
      negative_inputs_13_53_port, negative_inputs_13_52_port, 
      negative_inputs_13_51_port, negative_inputs_13_50_port, 
      negative_inputs_13_49_port, negative_inputs_13_48_port, 
      negative_inputs_13_47_port, negative_inputs_13_46_port, 
      negative_inputs_13_45_port, negative_inputs_13_44_port, 
      negative_inputs_13_43_port, negative_inputs_13_42_port, 
      negative_inputs_13_41_port, negative_inputs_13_40_port, 
      negative_inputs_13_39_port, negative_inputs_13_38_port, 
      negative_inputs_13_37_port, negative_inputs_13_36_port, 
      negative_inputs_13_35_port, negative_inputs_13_34_port, 
      negative_inputs_13_33_port, negative_inputs_13_32_port, 
      negative_inputs_13_31_port, negative_inputs_13_30_port, 
      negative_inputs_13_29_port, negative_inputs_13_28_port, 
      negative_inputs_13_27_port, negative_inputs_13_26_port, 
      negative_inputs_13_25_port, negative_inputs_13_24_port, 
      negative_inputs_13_23_port, negative_inputs_13_22_port, 
      negative_inputs_13_21_port, negative_inputs_13_20_port, 
      negative_inputs_13_19_port, negative_inputs_13_18_port, 
      negative_inputs_13_17_port, negative_inputs_13_16_port, 
      negative_inputs_13_15_port, negative_inputs_13_14_port, 
      negative_inputs_13_13_port, negative_inputs_13_12_port, 
      negative_inputs_13_11_port, negative_inputs_13_10_port, 
      negative_inputs_13_9_port, negative_inputs_13_8_port, 
      negative_inputs_13_7_port, negative_inputs_13_6_port, 
      negative_inputs_13_5_port, negative_inputs_13_4_port, 
      negative_inputs_13_3_port, negative_inputs_13_2_port, 
      negative_inputs_13_1_port, negative_inputs_12_63_port, 
      negative_inputs_12_62_port, negative_inputs_12_61_port, 
      negative_inputs_12_60_port, negative_inputs_12_59_port, 
      negative_inputs_12_58_port, negative_inputs_12_57_port, 
      negative_inputs_12_56_port, negative_inputs_12_55_port, 
      negative_inputs_12_54_port, negative_inputs_12_53_port, 
      negative_inputs_12_52_port, negative_inputs_12_51_port, 
      negative_inputs_12_50_port, negative_inputs_12_49_port, 
      negative_inputs_12_48_port, negative_inputs_12_47_port, 
      negative_inputs_12_46_port, negative_inputs_12_45_port, 
      negative_inputs_12_44_port, negative_inputs_12_43_port, 
      negative_inputs_12_42_port, negative_inputs_12_41_port, 
      negative_inputs_12_40_port, negative_inputs_12_39_port, 
      negative_inputs_12_38_port, negative_inputs_12_37_port, 
      negative_inputs_12_36_port, negative_inputs_12_35_port, 
      negative_inputs_12_34_port, negative_inputs_12_33_port, 
      negative_inputs_12_32_port, negative_inputs_12_31_port, 
      negative_inputs_12_30_port, negative_inputs_12_29_port, 
      negative_inputs_12_28_port, negative_inputs_12_27_port, 
      negative_inputs_12_26_port, negative_inputs_12_25_port, 
      negative_inputs_12_24_port, negative_inputs_12_23_port, 
      negative_inputs_12_22_port, negative_inputs_12_21_port, 
      negative_inputs_12_20_port, negative_inputs_12_19_port, 
      negative_inputs_12_18_port, negative_inputs_12_17_port, 
      negative_inputs_12_16_port, negative_inputs_12_15_port, 
      negative_inputs_12_14_port, negative_inputs_12_13_port, 
      negative_inputs_12_12_port, negative_inputs_12_11_port, 
      negative_inputs_12_10_port, negative_inputs_12_9_port, 
      negative_inputs_12_8_port, negative_inputs_12_7_port, 
      negative_inputs_12_6_port, negative_inputs_12_5_port, 
      negative_inputs_12_4_port, negative_inputs_12_3_port, 
      negative_inputs_12_2_port, negative_inputs_12_1_port, 
      negative_inputs_11_63_port, negative_inputs_11_62_port, 
      negative_inputs_11_61_port, negative_inputs_11_60_port, 
      negative_inputs_11_59_port, negative_inputs_11_58_port, 
      negative_inputs_11_57_port, negative_inputs_11_56_port, 
      negative_inputs_11_55_port, negative_inputs_11_54_port, 
      negative_inputs_11_53_port, negative_inputs_11_52_port, 
      negative_inputs_11_51_port, negative_inputs_11_50_port, 
      negative_inputs_11_49_port, negative_inputs_11_48_port, 
      negative_inputs_11_47_port, negative_inputs_11_46_port, 
      negative_inputs_11_45_port, negative_inputs_11_44_port, 
      negative_inputs_11_43_port, negative_inputs_11_42_port, 
      negative_inputs_11_41_port, negative_inputs_11_40_port, 
      negative_inputs_11_39_port, negative_inputs_11_38_port, 
      negative_inputs_11_37_port, negative_inputs_11_36_port, 
      negative_inputs_11_35_port, negative_inputs_11_34_port, 
      negative_inputs_11_33_port, negative_inputs_11_32_port, 
      negative_inputs_11_31_port, negative_inputs_11_30_port, 
      negative_inputs_11_29_port, negative_inputs_11_28_port, 
      negative_inputs_11_27_port, negative_inputs_11_26_port, 
      negative_inputs_11_25_port, negative_inputs_11_24_port, 
      negative_inputs_11_23_port, negative_inputs_11_22_port, 
      negative_inputs_11_21_port, negative_inputs_11_20_port, 
      negative_inputs_11_19_port, negative_inputs_11_18_port, 
      negative_inputs_11_17_port, negative_inputs_11_16_port, 
      negative_inputs_11_15_port, negative_inputs_11_14_port, 
      negative_inputs_11_13_port, negative_inputs_11_12_port, 
      negative_inputs_11_11_port, negative_inputs_11_10_port, 
      negative_inputs_11_9_port, negative_inputs_11_8_port, 
      negative_inputs_11_7_port, negative_inputs_11_6_port, 
      negative_inputs_11_5_port, negative_inputs_11_4_port, 
      negative_inputs_11_3_port, negative_inputs_11_2_port, 
      negative_inputs_11_1_port, negative_inputs_10_63_port, 
      negative_inputs_10_62_port, negative_inputs_10_61_port, 
      negative_inputs_10_60_port, negative_inputs_10_59_port, 
      negative_inputs_10_58_port, negative_inputs_10_57_port, 
      negative_inputs_10_56_port, negative_inputs_10_55_port, 
      negative_inputs_10_54_port, negative_inputs_10_53_port, 
      negative_inputs_10_52_port, negative_inputs_10_51_port, 
      negative_inputs_10_50_port, negative_inputs_10_49_port, 
      negative_inputs_10_48_port, negative_inputs_10_47_port, 
      negative_inputs_10_46_port, negative_inputs_10_45_port, 
      negative_inputs_10_44_port, negative_inputs_10_43_port, 
      negative_inputs_10_42_port, negative_inputs_10_41_port, 
      negative_inputs_10_40_port, negative_inputs_10_39_port, 
      negative_inputs_10_38_port, negative_inputs_10_37_port, 
      negative_inputs_10_36_port, negative_inputs_10_35_port, 
      negative_inputs_10_34_port, negative_inputs_10_33_port, 
      negative_inputs_10_32_port, negative_inputs_10_31_port, 
      negative_inputs_10_30_port, negative_inputs_10_29_port, 
      negative_inputs_10_28_port, negative_inputs_10_27_port, 
      negative_inputs_10_26_port, negative_inputs_10_25_port, 
      negative_inputs_10_24_port, negative_inputs_10_23_port, 
      negative_inputs_10_22_port, negative_inputs_10_21_port, 
      negative_inputs_10_20_port, negative_inputs_10_19_port, 
      negative_inputs_10_18_port, negative_inputs_10_17_port, 
      negative_inputs_10_16_port, negative_inputs_10_15_port, 
      negative_inputs_10_14_port, negative_inputs_10_13_port, 
      negative_inputs_10_12_port, negative_inputs_10_11_port, 
      negative_inputs_10_10_port, negative_inputs_10_9_port, 
      negative_inputs_10_8_port, negative_inputs_10_7_port, 
      negative_inputs_10_6_port, negative_inputs_10_5_port, 
      negative_inputs_10_4_port, negative_inputs_10_3_port, 
      negative_inputs_10_2_port, negative_inputs_10_1_port, 
      negative_inputs_9_63_port, negative_inputs_9_62_port, 
      negative_inputs_9_61_port, negative_inputs_9_60_port, 
      negative_inputs_9_59_port, negative_inputs_9_58_port, 
      negative_inputs_9_57_port, negative_inputs_9_56_port, 
      negative_inputs_9_55_port, negative_inputs_9_54_port, 
      negative_inputs_9_53_port, negative_inputs_9_52_port, 
      negative_inputs_9_51_port, negative_inputs_9_50_port, 
      negative_inputs_9_49_port, negative_inputs_9_48_port, 
      negative_inputs_9_47_port, negative_inputs_9_46_port, 
      negative_inputs_9_45_port, negative_inputs_9_44_port, 
      negative_inputs_9_43_port, negative_inputs_9_42_port, 
      negative_inputs_9_41_port, negative_inputs_9_40_port, 
      negative_inputs_9_39_port, negative_inputs_9_38_port, 
      negative_inputs_9_37_port, negative_inputs_9_36_port, 
      negative_inputs_9_35_port, negative_inputs_9_34_port, 
      negative_inputs_9_33_port, negative_inputs_9_32_port, 
      negative_inputs_9_31_port, negative_inputs_9_30_port, 
      negative_inputs_9_29_port, negative_inputs_9_28_port, 
      negative_inputs_9_27_port, negative_inputs_9_26_port, 
      negative_inputs_9_25_port, negative_inputs_9_24_port, 
      negative_inputs_9_23_port, negative_inputs_9_22_port, 
      negative_inputs_9_21_port, negative_inputs_9_20_port, 
      negative_inputs_9_19_port, negative_inputs_9_18_port, 
      negative_inputs_9_17_port, negative_inputs_9_16_port, 
      negative_inputs_9_15_port, negative_inputs_9_14_port, 
      negative_inputs_9_13_port, negative_inputs_9_12_port, 
      negative_inputs_9_11_port, negative_inputs_9_10_port, 
      negative_inputs_9_9_port, negative_inputs_9_8_port, 
      negative_inputs_9_7_port, negative_inputs_9_6_port, 
      negative_inputs_9_5_port, negative_inputs_9_4_port, 
      negative_inputs_9_3_port, negative_inputs_9_2_port, 
      negative_inputs_9_1_port, negative_inputs_24_63_port, 
      negative_inputs_24_62_port, negative_inputs_24_61_port, 
      negative_inputs_24_60_port, negative_inputs_24_59_port, 
      negative_inputs_24_58_port, negative_inputs_24_57_port, 
      negative_inputs_24_56_port, negative_inputs_24_55_port, 
      negative_inputs_24_54_port, negative_inputs_24_53_port, 
      negative_inputs_24_52_port, negative_inputs_24_51_port, 
      negative_inputs_24_50_port, negative_inputs_24_49_port, 
      negative_inputs_24_48_port, negative_inputs_24_47_port, 
      negative_inputs_24_46_port, negative_inputs_24_45_port, 
      negative_inputs_24_44_port, negative_inputs_24_43_port, 
      negative_inputs_24_42_port, negative_inputs_24_41_port, 
      negative_inputs_24_40_port, negative_inputs_24_39_port, 
      negative_inputs_24_38_port, negative_inputs_24_37_port, 
      negative_inputs_24_36_port, negative_inputs_24_35_port, 
      negative_inputs_24_34_port, negative_inputs_24_33_port, 
      negative_inputs_24_32_port, negative_inputs_24_31_port, 
      negative_inputs_24_30_port, negative_inputs_24_29_port, 
      negative_inputs_24_28_port, negative_inputs_24_27_port, 
      negative_inputs_24_26_port, negative_inputs_24_25_port, 
      negative_inputs_24_24_port, negative_inputs_24_23_port, 
      negative_inputs_24_22_port, negative_inputs_24_21_port, 
      negative_inputs_24_20_port, negative_inputs_24_19_port, 
      negative_inputs_24_18_port, negative_inputs_24_17_port, 
      negative_inputs_24_16_port, negative_inputs_24_15_port, 
      negative_inputs_24_14_port, negative_inputs_24_13_port, 
      negative_inputs_24_12_port, negative_inputs_24_11_port, 
      negative_inputs_24_10_port, negative_inputs_24_9_port, 
      negative_inputs_24_8_port, negative_inputs_24_7_port, 
      negative_inputs_24_6_port, negative_inputs_24_5_port, 
      negative_inputs_24_4_port, negative_inputs_24_3_port, 
      negative_inputs_24_2_port, negative_inputs_24_1_port, 
      negative_inputs_23_63_port, negative_inputs_23_62_port, 
      negative_inputs_23_61_port, negative_inputs_23_60_port, 
      negative_inputs_23_59_port, negative_inputs_23_58_port, 
      negative_inputs_23_57_port, negative_inputs_23_56_port, 
      negative_inputs_23_55_port, negative_inputs_23_54_port, 
      negative_inputs_23_53_port, negative_inputs_23_52_port, 
      negative_inputs_23_51_port, negative_inputs_23_50_port, 
      negative_inputs_23_49_port, negative_inputs_23_48_port, 
      negative_inputs_23_47_port, negative_inputs_23_46_port, 
      negative_inputs_23_45_port, negative_inputs_23_44_port, 
      negative_inputs_23_43_port, negative_inputs_23_42_port, 
      negative_inputs_23_41_port, negative_inputs_23_40_port, 
      negative_inputs_23_39_port, negative_inputs_23_38_port, 
      negative_inputs_23_37_port, negative_inputs_23_36_port, 
      negative_inputs_23_35_port, negative_inputs_23_34_port, 
      negative_inputs_23_33_port, negative_inputs_23_32_port, 
      negative_inputs_23_31_port, negative_inputs_23_30_port, 
      negative_inputs_23_29_port, negative_inputs_23_28_port, 
      negative_inputs_23_27_port, negative_inputs_23_26_port, 
      negative_inputs_23_25_port, negative_inputs_23_24_port, 
      negative_inputs_23_23_port, negative_inputs_23_22_port, 
      negative_inputs_23_21_port, negative_inputs_23_20_port, 
      negative_inputs_23_19_port, negative_inputs_23_18_port, 
      negative_inputs_23_17_port, negative_inputs_23_16_port, 
      negative_inputs_23_15_port, negative_inputs_23_14_port, 
      negative_inputs_23_13_port, negative_inputs_23_12_port, 
      negative_inputs_23_11_port, negative_inputs_23_10_port, 
      negative_inputs_23_9_port, negative_inputs_23_8_port, 
      negative_inputs_23_7_port, negative_inputs_23_6_port, 
      negative_inputs_23_5_port, negative_inputs_23_4_port, 
      negative_inputs_23_3_port, negative_inputs_23_2_port, 
      negative_inputs_23_1_port, negative_inputs_22_63_port, 
      negative_inputs_22_62_port, negative_inputs_22_61_port, 
      negative_inputs_22_60_port, negative_inputs_22_59_port, 
      negative_inputs_22_58_port, negative_inputs_22_57_port, 
      negative_inputs_22_56_port, negative_inputs_22_55_port, 
      negative_inputs_22_54_port, negative_inputs_22_53_port, 
      negative_inputs_22_52_port, negative_inputs_22_51_port, 
      negative_inputs_22_50_port, negative_inputs_22_49_port, 
      negative_inputs_22_48_port, negative_inputs_22_47_port, 
      negative_inputs_22_46_port, negative_inputs_22_45_port, 
      negative_inputs_22_44_port, negative_inputs_22_43_port, 
      negative_inputs_22_42_port, negative_inputs_22_41_port, 
      negative_inputs_22_40_port, negative_inputs_22_39_port, 
      negative_inputs_22_38_port, negative_inputs_22_37_port, 
      negative_inputs_22_36_port, negative_inputs_22_35_port, 
      negative_inputs_22_34_port, negative_inputs_22_33_port, 
      negative_inputs_22_32_port, negative_inputs_22_31_port, 
      negative_inputs_22_30_port, negative_inputs_22_29_port, 
      negative_inputs_22_28_port, negative_inputs_22_27_port, 
      negative_inputs_22_26_port, negative_inputs_22_25_port, 
      negative_inputs_22_24_port, negative_inputs_22_23_port, 
      negative_inputs_22_22_port, negative_inputs_22_21_port, 
      negative_inputs_22_20_port, negative_inputs_22_19_port, 
      negative_inputs_22_18_port, negative_inputs_22_17_port, 
      negative_inputs_22_16_port, negative_inputs_22_15_port, 
      negative_inputs_22_14_port, negative_inputs_22_13_port, 
      negative_inputs_22_12_port, negative_inputs_22_11_port, 
      negative_inputs_22_10_port, negative_inputs_22_9_port, 
      negative_inputs_22_8_port, negative_inputs_22_7_port, 
      negative_inputs_22_6_port, negative_inputs_22_5_port, 
      negative_inputs_22_4_port, negative_inputs_22_3_port, 
      negative_inputs_22_2_port, negative_inputs_22_1_port, 
      negative_inputs_21_63_port, negative_inputs_21_62_port, 
      negative_inputs_21_61_port, negative_inputs_21_60_port, 
      negative_inputs_21_59_port, negative_inputs_21_58_port, 
      negative_inputs_21_57_port, negative_inputs_21_56_port, 
      negative_inputs_21_55_port, negative_inputs_21_54_port, 
      negative_inputs_21_53_port, negative_inputs_21_52_port, 
      negative_inputs_21_51_port, negative_inputs_21_50_port, 
      negative_inputs_21_49_port, negative_inputs_21_48_port, 
      negative_inputs_21_47_port, negative_inputs_21_46_port, 
      negative_inputs_21_45_port, negative_inputs_21_44_port, 
      negative_inputs_21_43_port, negative_inputs_21_42_port, 
      negative_inputs_21_41_port, negative_inputs_21_40_port, 
      negative_inputs_21_39_port, negative_inputs_21_38_port, 
      negative_inputs_21_37_port, negative_inputs_21_36_port, 
      negative_inputs_21_35_port, negative_inputs_21_34_port, 
      negative_inputs_21_33_port, negative_inputs_21_32_port, 
      negative_inputs_21_31_port, negative_inputs_21_30_port, 
      negative_inputs_21_29_port, negative_inputs_21_28_port, 
      negative_inputs_21_27_port, negative_inputs_21_26_port, 
      negative_inputs_21_25_port, negative_inputs_21_24_port, 
      negative_inputs_21_23_port, negative_inputs_21_22_port, 
      negative_inputs_21_21_port, negative_inputs_21_20_port, 
      negative_inputs_21_19_port, negative_inputs_21_18_port, 
      negative_inputs_21_17_port, negative_inputs_21_16_port, 
      negative_inputs_21_15_port, negative_inputs_21_14_port, 
      negative_inputs_21_13_port, negative_inputs_21_12_port, 
      negative_inputs_21_11_port, negative_inputs_21_10_port, 
      negative_inputs_21_9_port, negative_inputs_21_8_port, 
      negative_inputs_21_7_port, negative_inputs_21_6_port, 
      negative_inputs_21_5_port, negative_inputs_21_4_port, 
      negative_inputs_21_3_port, negative_inputs_21_2_port, 
      negative_inputs_21_1_port, negative_inputs_20_63_port, 
      negative_inputs_20_62_port, negative_inputs_20_61_port, 
      negative_inputs_20_60_port, negative_inputs_20_59_port, 
      negative_inputs_20_58_port, negative_inputs_20_57_port, 
      negative_inputs_20_56_port, negative_inputs_20_55_port, 
      negative_inputs_20_54_port, negative_inputs_20_53_port, 
      negative_inputs_20_52_port, negative_inputs_20_51_port, 
      negative_inputs_20_50_port, negative_inputs_20_49_port, 
      negative_inputs_20_48_port, negative_inputs_20_47_port, 
      negative_inputs_20_46_port, negative_inputs_20_45_port, 
      negative_inputs_20_44_port, negative_inputs_20_43_port, 
      negative_inputs_20_42_port, negative_inputs_20_41_port, 
      negative_inputs_20_40_port, negative_inputs_20_39_port, 
      negative_inputs_20_38_port, negative_inputs_20_37_port, 
      negative_inputs_20_36_port, negative_inputs_20_35_port, 
      negative_inputs_20_34_port, negative_inputs_20_33_port, 
      negative_inputs_20_32_port, negative_inputs_20_31_port, 
      negative_inputs_20_30_port, negative_inputs_20_29_port, 
      negative_inputs_20_28_port, negative_inputs_20_27_port, 
      negative_inputs_20_26_port, negative_inputs_20_25_port, 
      negative_inputs_20_24_port, negative_inputs_20_23_port, 
      negative_inputs_20_22_port, negative_inputs_20_21_port, 
      negative_inputs_20_20_port, negative_inputs_20_19_port, 
      negative_inputs_20_18_port, negative_inputs_20_17_port, 
      negative_inputs_20_16_port, negative_inputs_20_15_port, 
      negative_inputs_20_14_port, negative_inputs_20_13_port, 
      negative_inputs_20_12_port, negative_inputs_20_11_port, 
      negative_inputs_20_10_port, negative_inputs_20_9_port, 
      negative_inputs_20_8_port, negative_inputs_20_7_port, 
      negative_inputs_20_6_port, negative_inputs_20_5_port, 
      negative_inputs_20_4_port, negative_inputs_20_3_port, 
      negative_inputs_20_2_port, negative_inputs_20_1_port, 
      negative_inputs_19_63_port, negative_inputs_19_62_port, 
      negative_inputs_19_61_port, negative_inputs_19_60_port, 
      negative_inputs_19_59_port, negative_inputs_19_58_port, 
      negative_inputs_19_57_port, negative_inputs_19_56_port, 
      negative_inputs_19_55_port, negative_inputs_19_54_port, 
      negative_inputs_19_53_port, negative_inputs_19_52_port, 
      negative_inputs_19_51_port, negative_inputs_19_50_port, 
      negative_inputs_19_49_port, negative_inputs_19_48_port, 
      negative_inputs_19_47_port, negative_inputs_19_46_port, 
      negative_inputs_19_45_port, negative_inputs_19_44_port, 
      negative_inputs_19_43_port, negative_inputs_19_42_port, 
      negative_inputs_19_41_port, negative_inputs_19_40_port, 
      negative_inputs_19_39_port, negative_inputs_19_38_port, 
      negative_inputs_19_37_port, negative_inputs_19_36_port, 
      negative_inputs_19_35_port, negative_inputs_19_34_port, 
      negative_inputs_19_33_port, negative_inputs_19_32_port, 
      negative_inputs_19_31_port, negative_inputs_19_30_port, 
      negative_inputs_19_29_port, negative_inputs_19_28_port, 
      negative_inputs_19_27_port, negative_inputs_19_26_port, 
      negative_inputs_19_25_port, negative_inputs_19_24_port, 
      negative_inputs_19_23_port, negative_inputs_19_22_port, 
      negative_inputs_19_21_port, negative_inputs_19_20_port, 
      negative_inputs_19_19_port, negative_inputs_19_18_port, 
      negative_inputs_19_17_port, negative_inputs_19_16_port, 
      negative_inputs_19_15_port, negative_inputs_19_14_port, 
      negative_inputs_19_13_port, negative_inputs_19_12_port, 
      negative_inputs_19_11_port, negative_inputs_19_10_port, 
      negative_inputs_19_9_port, negative_inputs_19_8_port, 
      negative_inputs_19_7_port, negative_inputs_19_6_port, 
      negative_inputs_19_5_port, negative_inputs_19_4_port, 
      negative_inputs_19_3_port, negative_inputs_19_2_port, 
      negative_inputs_19_1_port, negative_inputs_18_63_port, 
      negative_inputs_18_62_port, negative_inputs_18_61_port, 
      negative_inputs_18_60_port, negative_inputs_18_59_port, 
      negative_inputs_18_58_port, negative_inputs_18_57_port, 
      negative_inputs_18_56_port, negative_inputs_18_55_port, 
      negative_inputs_18_54_port, negative_inputs_18_53_port, 
      negative_inputs_18_52_port, negative_inputs_18_51_port, 
      negative_inputs_18_50_port, negative_inputs_18_49_port, 
      negative_inputs_18_48_port, negative_inputs_18_47_port, 
      negative_inputs_18_46_port, negative_inputs_18_45_port, 
      negative_inputs_18_44_port, negative_inputs_18_43_port, 
      negative_inputs_18_42_port, negative_inputs_18_41_port, 
      negative_inputs_18_40_port, negative_inputs_18_39_port, 
      negative_inputs_18_38_port, negative_inputs_18_37_port, 
      negative_inputs_18_36_port, negative_inputs_18_35_port, 
      negative_inputs_18_34_port, negative_inputs_18_33_port, 
      negative_inputs_18_32_port, negative_inputs_18_31_port, 
      negative_inputs_18_30_port, negative_inputs_18_29_port, 
      negative_inputs_18_28_port, negative_inputs_18_27_port, 
      negative_inputs_18_26_port, negative_inputs_18_25_port, 
      negative_inputs_18_24_port, negative_inputs_18_23_port, 
      negative_inputs_18_22_port, negative_inputs_18_21_port, 
      negative_inputs_18_20_port, negative_inputs_18_19_port, 
      negative_inputs_18_18_port, negative_inputs_18_17_port, 
      negative_inputs_18_16_port, negative_inputs_18_15_port, 
      negative_inputs_18_14_port, negative_inputs_18_13_port, 
      negative_inputs_18_12_port, negative_inputs_18_11_port, 
      negative_inputs_18_10_port, negative_inputs_18_9_port, 
      negative_inputs_18_8_port, negative_inputs_18_7_port, 
      negative_inputs_18_6_port, negative_inputs_18_5_port, 
      negative_inputs_18_4_port, negative_inputs_18_3_port, 
      negative_inputs_18_2_port, negative_inputs_18_1_port, 
      negative_inputs_17_63_port, negative_inputs_17_62_port, 
      negative_inputs_17_61_port, negative_inputs_17_60_port, 
      negative_inputs_17_59_port, negative_inputs_17_58_port, 
      negative_inputs_17_57_port, negative_inputs_17_56_port, 
      negative_inputs_17_55_port, negative_inputs_17_54_port, 
      negative_inputs_17_53_port, negative_inputs_17_52_port, 
      negative_inputs_17_51_port, negative_inputs_17_50_port, 
      negative_inputs_17_49_port, negative_inputs_17_48_port, 
      negative_inputs_17_47_port, negative_inputs_17_46_port, 
      negative_inputs_17_45_port, negative_inputs_17_44_port, 
      negative_inputs_17_43_port, negative_inputs_17_42_port, 
      negative_inputs_17_41_port, negative_inputs_17_40_port, 
      negative_inputs_17_39_port, negative_inputs_17_38_port, 
      negative_inputs_17_37_port, negative_inputs_17_36_port, 
      negative_inputs_17_35_port, negative_inputs_17_34_port, 
      negative_inputs_17_33_port, negative_inputs_17_32_port, 
      negative_inputs_17_31_port, negative_inputs_17_30_port, 
      negative_inputs_17_29_port, negative_inputs_17_28_port, 
      negative_inputs_17_27_port, negative_inputs_17_26_port, 
      negative_inputs_17_25_port, negative_inputs_17_24_port, 
      negative_inputs_17_23_port, negative_inputs_17_22_port, 
      negative_inputs_17_21_port, negative_inputs_17_20_port, 
      negative_inputs_17_19_port, negative_inputs_17_18_port, 
      negative_inputs_17_17_port, negative_inputs_17_16_port, 
      negative_inputs_17_15_port, negative_inputs_17_14_port, 
      negative_inputs_17_13_port, negative_inputs_17_12_port, 
      negative_inputs_17_11_port, negative_inputs_17_10_port, 
      negative_inputs_17_9_port, negative_inputs_17_8_port, 
      negative_inputs_17_7_port, negative_inputs_17_6_port, 
      negative_inputs_17_5_port, negative_inputs_17_4_port, 
      negative_inputs_17_3_port, negative_inputs_17_2_port, 
      negative_inputs_17_1_port, negative_inputs_31_63_port, 
      negative_inputs_31_62_port, negative_inputs_31_61_port, 
      negative_inputs_31_60_port, negative_inputs_31_59_port, 
      negative_inputs_31_58_port, negative_inputs_31_57_port, 
      negative_inputs_31_56_port, negative_inputs_31_55_port, 
      negative_inputs_31_54_port, negative_inputs_31_53_port, 
      negative_inputs_31_52_port, negative_inputs_31_51_port, 
      negative_inputs_31_50_port, negative_inputs_31_49_port, 
      negative_inputs_31_48_port, negative_inputs_31_47_port, 
      negative_inputs_31_46_port, negative_inputs_31_45_port, 
      negative_inputs_31_44_port, negative_inputs_31_43_port, 
      negative_inputs_31_42_port, negative_inputs_31_41_port, 
      negative_inputs_31_40_port, negative_inputs_31_39_port, 
      negative_inputs_31_38_port, negative_inputs_31_37_port, 
      negative_inputs_31_36_port, negative_inputs_31_35_port, 
      negative_inputs_31_34_port, negative_inputs_31_33_port, 
      negative_inputs_31_32_port, negative_inputs_31_31_port, 
      negative_inputs_31_30_port, negative_inputs_31_29_port, 
      negative_inputs_31_28_port, negative_inputs_31_27_port, 
      negative_inputs_31_26_port, negative_inputs_31_25_port, 
      negative_inputs_31_24_port, negative_inputs_31_23_port, 
      negative_inputs_31_22_port, negative_inputs_31_21_port, 
      negative_inputs_31_20_port, negative_inputs_31_19_port, 
      negative_inputs_31_18_port, negative_inputs_31_17_port, 
      negative_inputs_31_16_port, negative_inputs_31_15_port, 
      negative_inputs_31_14_port, negative_inputs_31_13_port, 
      negative_inputs_31_12_port, negative_inputs_31_11_port, 
      negative_inputs_31_10_port, negative_inputs_31_9_port, 
      negative_inputs_31_8_port, negative_inputs_31_7_port, 
      negative_inputs_31_6_port, negative_inputs_31_5_port, 
      negative_inputs_31_4_port, negative_inputs_31_3_port, 
      negative_inputs_31_2_port, negative_inputs_31_1_port, 
      negative_inputs_30_63_port, negative_inputs_30_62_port, 
      negative_inputs_30_61_port, negative_inputs_30_60_port, 
      negative_inputs_30_59_port, negative_inputs_30_58_port, 
      negative_inputs_30_57_port, negative_inputs_30_56_port, 
      negative_inputs_30_55_port, negative_inputs_30_54_port, 
      negative_inputs_30_53_port, negative_inputs_30_52_port, 
      negative_inputs_30_51_port, negative_inputs_30_50_port, 
      negative_inputs_30_49_port, negative_inputs_30_48_port, 
      negative_inputs_30_47_port, negative_inputs_30_46_port, 
      negative_inputs_30_45_port, negative_inputs_30_44_port, 
      negative_inputs_30_43_port, negative_inputs_30_42_port, 
      negative_inputs_30_41_port, negative_inputs_30_40_port, 
      negative_inputs_30_39_port, negative_inputs_30_38_port, 
      negative_inputs_30_37_port, negative_inputs_30_36_port, 
      negative_inputs_30_35_port, negative_inputs_30_34_port, 
      negative_inputs_30_33_port, negative_inputs_30_32_port, 
      negative_inputs_30_31_port, negative_inputs_30_30_port, 
      negative_inputs_30_29_port, negative_inputs_30_28_port, 
      negative_inputs_30_27_port, negative_inputs_30_26_port, 
      negative_inputs_30_25_port, negative_inputs_30_24_port, 
      negative_inputs_30_23_port, negative_inputs_30_22_port, 
      negative_inputs_30_21_port, negative_inputs_30_20_port, 
      negative_inputs_30_19_port, negative_inputs_30_18_port, 
      negative_inputs_30_17_port, negative_inputs_30_16_port, 
      negative_inputs_30_15_port, negative_inputs_30_14_port, 
      negative_inputs_30_13_port, negative_inputs_30_12_port, 
      negative_inputs_30_11_port, negative_inputs_30_10_port, 
      negative_inputs_30_9_port, negative_inputs_30_8_port, 
      negative_inputs_30_7_port, negative_inputs_30_6_port, 
      negative_inputs_30_5_port, negative_inputs_30_4_port, 
      negative_inputs_30_3_port, negative_inputs_30_2_port, 
      negative_inputs_30_1_port, negative_inputs_29_63_port, 
      negative_inputs_29_62_port, negative_inputs_29_61_port, 
      negative_inputs_29_60_port, negative_inputs_29_59_port, 
      negative_inputs_29_58_port, negative_inputs_29_57_port, 
      negative_inputs_29_56_port, negative_inputs_29_55_port, 
      negative_inputs_29_54_port, negative_inputs_29_53_port, 
      negative_inputs_29_52_port, negative_inputs_29_51_port, 
      negative_inputs_29_50_port, negative_inputs_29_49_port, 
      negative_inputs_29_48_port, negative_inputs_29_47_port, 
      negative_inputs_29_46_port, negative_inputs_29_45_port, 
      negative_inputs_29_44_port, negative_inputs_29_43_port, 
      negative_inputs_29_42_port, negative_inputs_29_41_port, 
      negative_inputs_29_40_port, negative_inputs_29_39_port, 
      negative_inputs_29_38_port, negative_inputs_29_37_port, 
      negative_inputs_29_36_port, negative_inputs_29_35_port, 
      negative_inputs_29_34_port, negative_inputs_29_33_port, 
      negative_inputs_29_32_port, negative_inputs_29_31_port, 
      negative_inputs_29_30_port, negative_inputs_29_29_port, 
      negative_inputs_29_28_port, negative_inputs_29_27_port, 
      negative_inputs_29_26_port, negative_inputs_29_25_port, 
      negative_inputs_29_24_port, negative_inputs_29_23_port, 
      negative_inputs_29_22_port, negative_inputs_29_21_port, 
      negative_inputs_29_20_port, negative_inputs_29_19_port, 
      negative_inputs_29_18_port, negative_inputs_29_17_port, 
      negative_inputs_29_16_port, negative_inputs_29_15_port, 
      negative_inputs_29_14_port, negative_inputs_29_13_port, 
      negative_inputs_29_12_port, negative_inputs_29_11_port, 
      negative_inputs_29_10_port, negative_inputs_29_9_port, 
      negative_inputs_29_8_port, negative_inputs_29_7_port, 
      negative_inputs_29_6_port, negative_inputs_29_5_port, 
      negative_inputs_29_4_port, negative_inputs_29_3_port, 
      negative_inputs_29_2_port, negative_inputs_29_1_port, 
      negative_inputs_28_63_port, negative_inputs_28_62_port, 
      negative_inputs_28_61_port, negative_inputs_28_60_port, 
      negative_inputs_28_59_port, negative_inputs_28_58_port, 
      negative_inputs_28_57_port, negative_inputs_28_56_port, 
      negative_inputs_28_55_port, negative_inputs_28_54_port, 
      negative_inputs_28_53_port, negative_inputs_28_52_port, 
      negative_inputs_28_51_port, negative_inputs_28_50_port, 
      negative_inputs_28_49_port, negative_inputs_28_48_port, 
      negative_inputs_28_47_port, negative_inputs_28_46_port, 
      negative_inputs_28_45_port, negative_inputs_28_44_port, 
      negative_inputs_28_43_port, negative_inputs_28_42_port, 
      negative_inputs_28_41_port, negative_inputs_28_40_port, 
      negative_inputs_28_39_port, negative_inputs_28_38_port, 
      negative_inputs_28_37_port, negative_inputs_28_36_port, 
      negative_inputs_28_35_port, negative_inputs_28_34_port, 
      negative_inputs_28_33_port, negative_inputs_28_32_port, 
      negative_inputs_28_31_port, negative_inputs_28_30_port, 
      negative_inputs_28_29_port, negative_inputs_28_28_port, 
      negative_inputs_28_27_port, negative_inputs_28_26_port, 
      negative_inputs_28_25_port, negative_inputs_28_24_port, 
      negative_inputs_28_23_port, negative_inputs_28_22_port, 
      negative_inputs_28_21_port, negative_inputs_28_20_port, 
      negative_inputs_28_19_port, negative_inputs_28_18_port, 
      negative_inputs_28_17_port, negative_inputs_28_16_port, 
      negative_inputs_28_15_port, negative_inputs_28_14_port, 
      negative_inputs_28_13_port, negative_inputs_28_12_port, 
      negative_inputs_28_11_port, negative_inputs_28_10_port, 
      negative_inputs_28_9_port, negative_inputs_28_8_port, 
      negative_inputs_28_7_port, negative_inputs_28_6_port, 
      negative_inputs_28_5_port, negative_inputs_28_4_port, 
      negative_inputs_28_3_port, negative_inputs_28_2_port, 
      negative_inputs_28_1_port, negative_inputs_27_63_port, 
      negative_inputs_27_62_port, negative_inputs_27_61_port, 
      negative_inputs_27_60_port, negative_inputs_27_59_port, 
      negative_inputs_27_58_port, negative_inputs_27_57_port, 
      negative_inputs_27_56_port, negative_inputs_27_55_port, 
      negative_inputs_27_54_port, negative_inputs_27_53_port, 
      negative_inputs_27_52_port, negative_inputs_27_51_port, 
      negative_inputs_27_50_port, negative_inputs_27_49_port, 
      negative_inputs_27_48_port, negative_inputs_27_47_port, 
      negative_inputs_27_46_port, negative_inputs_27_45_port, 
      negative_inputs_27_44_port, negative_inputs_27_43_port, 
      negative_inputs_27_42_port, negative_inputs_27_41_port, 
      negative_inputs_27_40_port, negative_inputs_27_39_port, 
      negative_inputs_27_38_port, negative_inputs_27_37_port, 
      negative_inputs_27_36_port, negative_inputs_27_35_port, 
      negative_inputs_27_34_port, negative_inputs_27_33_port, 
      negative_inputs_27_32_port, negative_inputs_27_31_port, 
      negative_inputs_27_30_port, negative_inputs_27_29_port, 
      negative_inputs_27_28_port, negative_inputs_27_27_port, 
      negative_inputs_27_26_port, negative_inputs_27_25_port, 
      negative_inputs_27_24_port, negative_inputs_27_23_port, 
      negative_inputs_27_22_port, negative_inputs_27_21_port, 
      negative_inputs_27_20_port, negative_inputs_27_19_port, 
      negative_inputs_27_18_port, negative_inputs_27_17_port, 
      negative_inputs_27_16_port, negative_inputs_27_15_port, 
      negative_inputs_27_14_port, negative_inputs_27_13_port, 
      negative_inputs_27_12_port, negative_inputs_27_11_port, 
      negative_inputs_27_10_port, negative_inputs_27_9_port, 
      negative_inputs_27_8_port, negative_inputs_27_7_port, 
      negative_inputs_27_6_port, negative_inputs_27_5_port, 
      negative_inputs_27_4_port, negative_inputs_27_3_port, 
      negative_inputs_27_2_port, negative_inputs_27_1_port, 
      negative_inputs_26_63_port, negative_inputs_26_62_port, 
      negative_inputs_26_61_port, negative_inputs_26_60_port, 
      negative_inputs_26_59_port, negative_inputs_26_58_port, 
      negative_inputs_26_57_port, negative_inputs_26_56_port, 
      negative_inputs_26_55_port, negative_inputs_26_54_port, 
      negative_inputs_26_53_port, negative_inputs_26_52_port, 
      negative_inputs_26_51_port, negative_inputs_26_50_port, 
      negative_inputs_26_49_port, negative_inputs_26_48_port, 
      negative_inputs_26_47_port, negative_inputs_26_46_port, 
      negative_inputs_26_45_port, negative_inputs_26_44_port, 
      negative_inputs_26_43_port, negative_inputs_26_42_port, 
      negative_inputs_26_41_port, negative_inputs_26_40_port, 
      negative_inputs_26_39_port, negative_inputs_26_38_port, 
      negative_inputs_26_37_port, negative_inputs_26_36_port, 
      negative_inputs_26_35_port, negative_inputs_26_34_port, 
      negative_inputs_26_33_port, negative_inputs_26_32_port, 
      negative_inputs_26_31_port, negative_inputs_26_30_port, 
      negative_inputs_26_29_port, negative_inputs_26_28_port, 
      negative_inputs_26_27_port, negative_inputs_26_26_port, 
      negative_inputs_26_25_port, negative_inputs_26_24_port, 
      negative_inputs_26_23_port, negative_inputs_26_22_port, 
      negative_inputs_26_21_port, negative_inputs_26_20_port, 
      negative_inputs_26_19_port, negative_inputs_26_18_port, 
      negative_inputs_26_17_port, negative_inputs_26_16_port, 
      negative_inputs_26_15_port, negative_inputs_26_14_port, 
      negative_inputs_26_13_port, negative_inputs_26_12_port, 
      negative_inputs_26_11_port, negative_inputs_26_10_port, 
      negative_inputs_26_9_port, negative_inputs_26_8_port, 
      negative_inputs_26_7_port, negative_inputs_26_6_port, 
      negative_inputs_26_5_port, negative_inputs_26_4_port, 
      negative_inputs_26_3_port, negative_inputs_26_2_port, 
      negative_inputs_26_1_port, negative_inputs_25_63_port, 
      negative_inputs_25_62_port, negative_inputs_25_61_port, 
      negative_inputs_25_60_port, negative_inputs_25_59_port, 
      negative_inputs_25_58_port, negative_inputs_25_57_port, 
      negative_inputs_25_56_port, negative_inputs_25_55_port, 
      negative_inputs_25_54_port, negative_inputs_25_53_port, 
      negative_inputs_25_52_port, negative_inputs_25_51_port, 
      negative_inputs_25_50_port, negative_inputs_25_49_port, 
      negative_inputs_25_48_port, negative_inputs_25_47_port, 
      negative_inputs_25_46_port, negative_inputs_25_45_port, 
      negative_inputs_25_44_port, negative_inputs_25_43_port, 
      negative_inputs_25_42_port, negative_inputs_25_41_port, 
      negative_inputs_25_40_port, negative_inputs_25_39_port, 
      negative_inputs_25_38_port, negative_inputs_25_37_port, 
      negative_inputs_25_36_port, negative_inputs_25_35_port, 
      negative_inputs_25_34_port, negative_inputs_25_33_port, 
      negative_inputs_25_32_port, negative_inputs_25_31_port, 
      negative_inputs_25_30_port, negative_inputs_25_29_port, 
      negative_inputs_25_28_port, negative_inputs_25_27_port, 
      negative_inputs_25_26_port, negative_inputs_25_25_port, 
      negative_inputs_25_24_port, negative_inputs_25_23_port, 
      negative_inputs_25_22_port, negative_inputs_25_21_port, 
      negative_inputs_25_20_port, negative_inputs_25_19_port, 
      negative_inputs_25_18_port, negative_inputs_25_17_port, 
      negative_inputs_25_16_port, negative_inputs_25_15_port, 
      negative_inputs_25_14_port, negative_inputs_25_13_port, 
      negative_inputs_25_12_port, negative_inputs_25_11_port, 
      negative_inputs_25_10_port, negative_inputs_25_9_port, 
      negative_inputs_25_8_port, negative_inputs_25_7_port, 
      negative_inputs_25_6_port, negative_inputs_25_5_port, 
      negative_inputs_25_4_port, negative_inputs_25_3_port, 
      negative_inputs_25_2_port, negative_inputs_25_1_port, sel_15_2_port, 
      sel_15_1_port, sel_15_0_port, sel_14_2_port, sel_14_1_port, sel_14_0_port
      , sel_13_2_port, sel_13_1_port, sel_13_0_port, sel_12_2_port, 
      sel_12_1_port, sel_12_0_port, sel_11_2_port, sel_11_1_port, sel_11_0_port
      , sel_10_2_port, sel_10_1_port, sel_10_0_port, sel_9_2_port, sel_9_1_port
      , sel_9_0_port, sel_8_2_port, sel_8_1_port, sel_8_0_port, sel_7_2_port, 
      sel_7_1_port, sel_7_0_port, sel_6_2_port, sel_6_1_port, sel_6_0_port, 
      sel_5_2_port, sel_5_1_port, sel_5_0_port, sel_4_2_port, sel_4_1_port, 
      sel_4_0_port, sel_3_2_port, sel_3_1_port, sel_3_0_port, sel_2_2_port, 
      sel_2_1_port, sel_2_0_port, sel_1_2_port, sel_1_1_port, sel_1_0_port, 
      sel_0_2_port, sel_0_1_port, sel_0_0_port, MuxOutputs_7_63_port, 
      MuxOutputs_7_62_port, MuxOutputs_7_61_port, MuxOutputs_7_60_port, 
      MuxOutputs_7_59_port, MuxOutputs_7_58_port, MuxOutputs_7_57_port, 
      MuxOutputs_7_56_port, MuxOutputs_7_55_port, MuxOutputs_7_54_port, 
      MuxOutputs_7_53_port, MuxOutputs_7_52_port, MuxOutputs_7_51_port, 
      MuxOutputs_7_50_port, MuxOutputs_7_49_port, MuxOutputs_7_48_port, 
      MuxOutputs_7_47_port, MuxOutputs_7_46_port, MuxOutputs_7_45_port, 
      MuxOutputs_7_44_port, MuxOutputs_7_43_port, MuxOutputs_7_42_port, 
      MuxOutputs_7_41_port, MuxOutputs_7_40_port, MuxOutputs_7_39_port, 
      MuxOutputs_7_38_port, MuxOutputs_7_37_port, MuxOutputs_7_36_port, 
      MuxOutputs_7_35_port, MuxOutputs_7_34_port, MuxOutputs_7_33_port, 
      MuxOutputs_7_32_port, MuxOutputs_7_31_port, MuxOutputs_7_30_port, 
      MuxOutputs_7_29_port, MuxOutputs_7_28_port, MuxOutputs_7_27_port, 
      MuxOutputs_7_26_port, MuxOutputs_7_25_port, MuxOutputs_7_24_port, 
      MuxOutputs_7_23_port, MuxOutputs_7_22_port, MuxOutputs_7_21_port, 
      MuxOutputs_7_20_port, MuxOutputs_7_19_port, MuxOutputs_7_18_port, 
      MuxOutputs_7_17_port, MuxOutputs_7_16_port, MuxOutputs_7_15_port, 
      MuxOutputs_7_14_port, MuxOutputs_7_13_port, MuxOutputs_7_12_port, 
      MuxOutputs_7_11_port, MuxOutputs_7_10_port, MuxOutputs_7_9_port, 
      MuxOutputs_7_8_port, MuxOutputs_7_7_port, MuxOutputs_7_6_port, 
      MuxOutputs_7_5_port, MuxOutputs_7_4_port, MuxOutputs_7_3_port, 
      MuxOutputs_7_2_port, MuxOutputs_7_1_port, MuxOutputs_7_0_port, 
      MuxOutputs_6_63_port, MuxOutputs_6_62_port, MuxOutputs_6_61_port, 
      MuxOutputs_6_60_port, MuxOutputs_6_59_port, MuxOutputs_6_58_port, 
      MuxOutputs_6_57_port, MuxOutputs_6_56_port, MuxOutputs_6_55_port, 
      MuxOutputs_6_54_port, MuxOutputs_6_53_port, MuxOutputs_6_52_port, 
      MuxOutputs_6_51_port, MuxOutputs_6_50_port, MuxOutputs_6_49_port, 
      MuxOutputs_6_48_port, MuxOutputs_6_47_port, MuxOutputs_6_46_port, 
      MuxOutputs_6_45_port, MuxOutputs_6_44_port, MuxOutputs_6_43_port, 
      MuxOutputs_6_42_port, MuxOutputs_6_41_port, MuxOutputs_6_40_port, 
      MuxOutputs_6_39_port, MuxOutputs_6_38_port, MuxOutputs_6_37_port, 
      MuxOutputs_6_36_port, MuxOutputs_6_35_port, MuxOutputs_6_34_port, 
      MuxOutputs_6_33_port, MuxOutputs_6_32_port, MuxOutputs_6_31_port, 
      MuxOutputs_6_30_port, MuxOutputs_6_29_port, MuxOutputs_6_28_port, 
      MuxOutputs_6_27_port, MuxOutputs_6_26_port, MuxOutputs_6_25_port, 
      MuxOutputs_6_24_port, MuxOutputs_6_23_port, MuxOutputs_6_22_port, 
      MuxOutputs_6_21_port, MuxOutputs_6_20_port, MuxOutputs_6_19_port, 
      MuxOutputs_6_18_port, MuxOutputs_6_17_port, MuxOutputs_6_16_port, 
      MuxOutputs_6_15_port, MuxOutputs_6_14_port, MuxOutputs_6_13_port, 
      MuxOutputs_6_12_port, MuxOutputs_6_11_port, MuxOutputs_6_10_port, 
      MuxOutputs_6_9_port, MuxOutputs_6_8_port, MuxOutputs_6_7_port, 
      MuxOutputs_6_6_port, MuxOutputs_6_5_port, MuxOutputs_6_4_port, 
      MuxOutputs_6_3_port, MuxOutputs_6_2_port, MuxOutputs_6_1_port, 
      MuxOutputs_6_0_port, MuxOutputs_5_63_port, MuxOutputs_5_62_port, 
      MuxOutputs_5_61_port, MuxOutputs_5_60_port, MuxOutputs_5_59_port, 
      MuxOutputs_5_58_port, MuxOutputs_5_57_port, MuxOutputs_5_56_port, 
      MuxOutputs_5_55_port, MuxOutputs_5_54_port, MuxOutputs_5_53_port, 
      MuxOutputs_5_52_port, MuxOutputs_5_51_port, MuxOutputs_5_50_port, 
      MuxOutputs_5_49_port, MuxOutputs_5_48_port, MuxOutputs_5_47_port, 
      MuxOutputs_5_46_port, MuxOutputs_5_45_port, MuxOutputs_5_44_port, 
      MuxOutputs_5_43_port, MuxOutputs_5_42_port, MuxOutputs_5_41_port, 
      MuxOutputs_5_40_port, MuxOutputs_5_39_port, MuxOutputs_5_38_port, 
      MuxOutputs_5_37_port, MuxOutputs_5_36_port, MuxOutputs_5_35_port, 
      MuxOutputs_5_34_port, MuxOutputs_5_33_port, MuxOutputs_5_32_port, 
      MuxOutputs_5_31_port, MuxOutputs_5_30_port, MuxOutputs_5_29_port, 
      MuxOutputs_5_28_port, MuxOutputs_5_27_port, MuxOutputs_5_26_port, 
      MuxOutputs_5_25_port, MuxOutputs_5_24_port, MuxOutputs_5_23_port, 
      MuxOutputs_5_22_port, MuxOutputs_5_21_port, MuxOutputs_5_20_port, 
      MuxOutputs_5_19_port, MuxOutputs_5_18_port, MuxOutputs_5_17_port, 
      MuxOutputs_5_16_port, MuxOutputs_5_15_port, MuxOutputs_5_14_port, 
      MuxOutputs_5_13_port, MuxOutputs_5_12_port, MuxOutputs_5_11_port, 
      MuxOutputs_5_10_port, MuxOutputs_5_9_port, MuxOutputs_5_8_port, 
      MuxOutputs_5_7_port, MuxOutputs_5_6_port, MuxOutputs_5_5_port, 
      MuxOutputs_5_4_port, MuxOutputs_5_3_port, MuxOutputs_5_2_port, 
      MuxOutputs_5_1_port, MuxOutputs_5_0_port, MuxOutputs_4_63_port, 
      MuxOutputs_4_62_port, MuxOutputs_4_61_port, MuxOutputs_4_60_port, 
      MuxOutputs_4_59_port, MuxOutputs_4_58_port, MuxOutputs_4_57_port, 
      MuxOutputs_4_56_port, MuxOutputs_4_55_port, MuxOutputs_4_54_port, 
      MuxOutputs_4_53_port, MuxOutputs_4_52_port, MuxOutputs_4_51_port, 
      MuxOutputs_4_50_port, MuxOutputs_4_49_port, MuxOutputs_4_48_port, 
      MuxOutputs_4_47_port, MuxOutputs_4_46_port, MuxOutputs_4_45_port, 
      MuxOutputs_4_44_port, MuxOutputs_4_43_port, MuxOutputs_4_42_port, 
      MuxOutputs_4_41_port, MuxOutputs_4_40_port, MuxOutputs_4_39_port, 
      MuxOutputs_4_38_port, MuxOutputs_4_37_port, MuxOutputs_4_36_port, 
      MuxOutputs_4_35_port, MuxOutputs_4_34_port, MuxOutputs_4_33_port, 
      MuxOutputs_4_32_port, MuxOutputs_4_31_port, MuxOutputs_4_30_port, 
      MuxOutputs_4_29_port, MuxOutputs_4_28_port, MuxOutputs_4_27_port, 
      MuxOutputs_4_26_port, MuxOutputs_4_25_port, MuxOutputs_4_24_port, 
      MuxOutputs_4_23_port, MuxOutputs_4_22_port, MuxOutputs_4_21_port, 
      MuxOutputs_4_20_port, MuxOutputs_4_19_port, MuxOutputs_4_18_port, 
      MuxOutputs_4_17_port, MuxOutputs_4_16_port, MuxOutputs_4_15_port, 
      MuxOutputs_4_14_port, MuxOutputs_4_13_port, MuxOutputs_4_12_port, 
      MuxOutputs_4_11_port, MuxOutputs_4_10_port, MuxOutputs_4_9_port, 
      MuxOutputs_4_8_port, MuxOutputs_4_7_port, MuxOutputs_4_6_port, 
      MuxOutputs_4_5_port, MuxOutputs_4_4_port, MuxOutputs_4_3_port, 
      MuxOutputs_4_2_port, MuxOutputs_4_1_port, MuxOutputs_4_0_port, 
      MuxOutputs_3_63_port, MuxOutputs_3_62_port, MuxOutputs_3_61_port, 
      MuxOutputs_3_60_port, MuxOutputs_3_59_port, MuxOutputs_3_58_port, 
      MuxOutputs_3_57_port, MuxOutputs_3_56_port, MuxOutputs_3_55_port, 
      MuxOutputs_3_54_port, MuxOutputs_3_53_port, MuxOutputs_3_52_port, 
      MuxOutputs_3_51_port, MuxOutputs_3_50_port, MuxOutputs_3_49_port, 
      MuxOutputs_3_48_port, MuxOutputs_3_47_port, MuxOutputs_3_46_port, 
      MuxOutputs_3_45_port, MuxOutputs_3_44_port, MuxOutputs_3_43_port, 
      MuxOutputs_3_42_port, MuxOutputs_3_41_port, MuxOutputs_3_40_port, 
      MuxOutputs_3_39_port, MuxOutputs_3_38_port, MuxOutputs_3_37_port, 
      MuxOutputs_3_36_port, MuxOutputs_3_35_port, MuxOutputs_3_34_port, 
      MuxOutputs_3_33_port, MuxOutputs_3_32_port, MuxOutputs_3_31_port, 
      MuxOutputs_3_30_port, MuxOutputs_3_29_port, MuxOutputs_3_28_port, 
      MuxOutputs_3_27_port, MuxOutputs_3_26_port, MuxOutputs_3_25_port, 
      MuxOutputs_3_24_port, MuxOutputs_3_23_port, MuxOutputs_3_22_port, 
      MuxOutputs_3_21_port, MuxOutputs_3_20_port, MuxOutputs_3_19_port, 
      MuxOutputs_3_18_port, MuxOutputs_3_17_port, MuxOutputs_3_16_port, 
      MuxOutputs_3_15_port, MuxOutputs_3_14_port, MuxOutputs_3_13_port, 
      MuxOutputs_3_12_port, MuxOutputs_3_11_port, MuxOutputs_3_10_port, 
      MuxOutputs_3_9_port, MuxOutputs_3_8_port, MuxOutputs_3_7_port, 
      MuxOutputs_3_6_port, MuxOutputs_3_5_port, MuxOutputs_3_4_port, 
      MuxOutputs_3_3_port, MuxOutputs_3_2_port, MuxOutputs_3_1_port, 
      MuxOutputs_3_0_port, MuxOutputs_2_63_port, MuxOutputs_2_62_port, 
      MuxOutputs_2_61_port, MuxOutputs_2_60_port, MuxOutputs_2_59_port, 
      MuxOutputs_2_58_port, MuxOutputs_2_57_port, MuxOutputs_2_56_port, 
      MuxOutputs_2_55_port, MuxOutputs_2_54_port, MuxOutputs_2_53_port, 
      MuxOutputs_2_52_port, MuxOutputs_2_51_port, MuxOutputs_2_50_port, 
      MuxOutputs_2_49_port, MuxOutputs_2_48_port, MuxOutputs_2_47_port, 
      MuxOutputs_2_46_port, MuxOutputs_2_45_port, MuxOutputs_2_44_port, 
      MuxOutputs_2_43_port, MuxOutputs_2_42_port, MuxOutputs_2_41_port, 
      MuxOutputs_2_40_port, MuxOutputs_2_39_port, MuxOutputs_2_38_port, 
      MuxOutputs_2_37_port, MuxOutputs_2_36_port, MuxOutputs_2_35_port, 
      MuxOutputs_2_34_port, MuxOutputs_2_33_port, MuxOutputs_2_32_port, 
      MuxOutputs_2_31_port, MuxOutputs_2_30_port, MuxOutputs_2_29_port, 
      MuxOutputs_2_28_port, MuxOutputs_2_27_port, MuxOutputs_2_26_port, 
      MuxOutputs_2_25_port, MuxOutputs_2_24_port, MuxOutputs_2_23_port, 
      MuxOutputs_2_22_port, MuxOutputs_2_21_port, MuxOutputs_2_20_port, 
      MuxOutputs_2_19_port, MuxOutputs_2_18_port, MuxOutputs_2_17_port, 
      MuxOutputs_2_16_port, MuxOutputs_2_15_port, MuxOutputs_2_14_port, 
      MuxOutputs_2_13_port, MuxOutputs_2_12_port, MuxOutputs_2_11_port, 
      MuxOutputs_2_10_port, MuxOutputs_2_9_port, MuxOutputs_2_8_port, 
      MuxOutputs_2_7_port, MuxOutputs_2_6_port, MuxOutputs_2_5_port, 
      MuxOutputs_2_4_port, MuxOutputs_2_3_port, MuxOutputs_2_2_port, 
      MuxOutputs_2_1_port, MuxOutputs_2_0_port, MuxOutputs_1_63_port, 
      MuxOutputs_1_62_port, MuxOutputs_1_61_port, MuxOutputs_1_60_port, 
      MuxOutputs_1_59_port, MuxOutputs_1_58_port, MuxOutputs_1_57_port, 
      MuxOutputs_1_56_port, MuxOutputs_1_55_port, MuxOutputs_1_54_port, 
      MuxOutputs_1_53_port, MuxOutputs_1_52_port, MuxOutputs_1_51_port, 
      MuxOutputs_1_50_port, MuxOutputs_1_49_port, MuxOutputs_1_48_port, 
      MuxOutputs_1_47_port, MuxOutputs_1_46_port, MuxOutputs_1_45_port, 
      MuxOutputs_1_44_port, MuxOutputs_1_43_port, MuxOutputs_1_42_port, 
      MuxOutputs_1_41_port, MuxOutputs_1_40_port, MuxOutputs_1_39_port, 
      MuxOutputs_1_38_port, MuxOutputs_1_37_port, MuxOutputs_1_36_port, 
      MuxOutputs_1_35_port, MuxOutputs_1_34_port, MuxOutputs_1_33_port, 
      MuxOutputs_1_32_port, MuxOutputs_1_31_port, MuxOutputs_1_30_port, 
      MuxOutputs_1_29_port, MuxOutputs_1_28_port, MuxOutputs_1_27_port, 
      MuxOutputs_1_26_port, MuxOutputs_1_25_port, MuxOutputs_1_24_port, 
      MuxOutputs_1_23_port, MuxOutputs_1_22_port, MuxOutputs_1_21_port, 
      MuxOutputs_1_20_port, MuxOutputs_1_19_port, MuxOutputs_1_18_port, 
      MuxOutputs_1_17_port, MuxOutputs_1_16_port, MuxOutputs_1_15_port, 
      MuxOutputs_1_14_port, MuxOutputs_1_13_port, MuxOutputs_1_12_port, 
      MuxOutputs_1_11_port, MuxOutputs_1_10_port, MuxOutputs_1_9_port, 
      MuxOutputs_1_8_port, MuxOutputs_1_7_port, MuxOutputs_1_6_port, 
      MuxOutputs_1_5_port, MuxOutputs_1_4_port, MuxOutputs_1_3_port, 
      MuxOutputs_1_2_port, MuxOutputs_1_1_port, MuxOutputs_1_0_port, 
      MuxOutputs_0_63_port, MuxOutputs_0_62_port, MuxOutputs_0_61_port, 
      MuxOutputs_0_60_port, MuxOutputs_0_59_port, MuxOutputs_0_58_port, 
      MuxOutputs_0_57_port, MuxOutputs_0_56_port, MuxOutputs_0_55_port, 
      MuxOutputs_0_54_port, MuxOutputs_0_53_port, MuxOutputs_0_52_port, 
      MuxOutputs_0_51_port, MuxOutputs_0_50_port, MuxOutputs_0_49_port, 
      MuxOutputs_0_48_port, MuxOutputs_0_47_port, MuxOutputs_0_46_port, 
      MuxOutputs_0_45_port, MuxOutputs_0_44_port, MuxOutputs_0_43_port, 
      MuxOutputs_0_42_port, MuxOutputs_0_41_port, MuxOutputs_0_40_port, 
      MuxOutputs_0_39_port, MuxOutputs_0_38_port, MuxOutputs_0_37_port, 
      MuxOutputs_0_36_port, MuxOutputs_0_35_port, MuxOutputs_0_34_port, 
      MuxOutputs_0_33_port, MuxOutputs_0_32_port, MuxOutputs_0_31_port, 
      MuxOutputs_0_30_port, MuxOutputs_0_29_port, MuxOutputs_0_28_port, 
      MuxOutputs_0_27_port, MuxOutputs_0_26_port, MuxOutputs_0_25_port, 
      MuxOutputs_0_24_port, MuxOutputs_0_23_port, MuxOutputs_0_22_port, 
      MuxOutputs_0_21_port, MuxOutputs_0_20_port, MuxOutputs_0_19_port, 
      MuxOutputs_0_18_port, MuxOutputs_0_17_port, MuxOutputs_0_16_port, 
      MuxOutputs_0_15_port, MuxOutputs_0_14_port, MuxOutputs_0_13_port, 
      MuxOutputs_0_12_port, MuxOutputs_0_11_port, MuxOutputs_0_10_port, 
      MuxOutputs_0_9_port, MuxOutputs_0_8_port, MuxOutputs_0_7_port, 
      MuxOutputs_0_6_port, MuxOutputs_0_5_port, MuxOutputs_0_4_port, 
      MuxOutputs_0_3_port, MuxOutputs_0_2_port, MuxOutputs_0_1_port, 
      MuxOutputs_0_0_port, MuxOutputs_15_63_port, MuxOutputs_15_62_port, 
      MuxOutputs_15_61_port, MuxOutputs_15_60_port, MuxOutputs_15_59_port, 
      MuxOutputs_15_58_port, MuxOutputs_15_57_port, MuxOutputs_15_56_port, 
      MuxOutputs_15_55_port, MuxOutputs_15_54_port, MuxOutputs_15_53_port, 
      MuxOutputs_15_52_port, MuxOutputs_15_51_port, MuxOutputs_15_50_port, 
      MuxOutputs_15_49_port, MuxOutputs_15_48_port, MuxOutputs_15_47_port, 
      MuxOutputs_15_46_port, MuxOutputs_15_45_port, MuxOutputs_15_44_port, 
      MuxOutputs_15_43_port, MuxOutputs_15_42_port, MuxOutputs_15_41_port, 
      MuxOutputs_15_40_port, MuxOutputs_15_39_port, MuxOutputs_15_38_port, 
      MuxOutputs_15_37_port, MuxOutputs_15_36_port, MuxOutputs_15_35_port, 
      MuxOutputs_15_34_port, MuxOutputs_15_33_port, MuxOutputs_15_32_port, 
      MuxOutputs_15_31_port, MuxOutputs_15_30_port, MuxOutputs_15_29_port, 
      MuxOutputs_15_28_port, MuxOutputs_15_27_port, MuxOutputs_15_26_port, 
      MuxOutputs_15_25_port, MuxOutputs_15_24_port, MuxOutputs_15_23_port, 
      MuxOutputs_15_22_port, MuxOutputs_15_21_port, MuxOutputs_15_20_port, 
      MuxOutputs_15_19_port, MuxOutputs_15_18_port, MuxOutputs_15_17_port, 
      MuxOutputs_15_16_port, MuxOutputs_15_15_port, MuxOutputs_15_14_port, 
      MuxOutputs_15_13_port, MuxOutputs_15_12_port, MuxOutputs_15_11_port, 
      MuxOutputs_15_10_port, MuxOutputs_15_9_port, MuxOutputs_15_8_port, 
      MuxOutputs_15_7_port, MuxOutputs_15_6_port, MuxOutputs_15_5_port, 
      MuxOutputs_15_4_port, MuxOutputs_15_3_port, MuxOutputs_15_2_port, 
      MuxOutputs_15_1_port, MuxOutputs_15_0_port, MuxOutputs_14_63_port, 
      MuxOutputs_14_62_port, MuxOutputs_14_61_port, MuxOutputs_14_60_port, 
      MuxOutputs_14_59_port, MuxOutputs_14_58_port, MuxOutputs_14_57_port, 
      MuxOutputs_14_56_port, MuxOutputs_14_55_port, MuxOutputs_14_54_port, 
      MuxOutputs_14_53_port, MuxOutputs_14_52_port, MuxOutputs_14_51_port, 
      MuxOutputs_14_50_port, MuxOutputs_14_49_port, MuxOutputs_14_48_port, 
      MuxOutputs_14_47_port, MuxOutputs_14_46_port, MuxOutputs_14_45_port, 
      MuxOutputs_14_44_port, MuxOutputs_14_43_port, MuxOutputs_14_42_port, 
      MuxOutputs_14_41_port, MuxOutputs_14_40_port, MuxOutputs_14_39_port, 
      MuxOutputs_14_38_port, MuxOutputs_14_37_port, MuxOutputs_14_36_port, 
      MuxOutputs_14_35_port, MuxOutputs_14_34_port, MuxOutputs_14_33_port, 
      MuxOutputs_14_32_port, MuxOutputs_14_31_port, MuxOutputs_14_30_port, 
      MuxOutputs_14_29_port, MuxOutputs_14_28_port, MuxOutputs_14_27_port, 
      MuxOutputs_14_26_port, MuxOutputs_14_25_port, MuxOutputs_14_24_port, 
      MuxOutputs_14_23_port, MuxOutputs_14_22_port, MuxOutputs_14_21_port, 
      MuxOutputs_14_20_port, MuxOutputs_14_19_port, MuxOutputs_14_18_port, 
      MuxOutputs_14_17_port, MuxOutputs_14_16_port, MuxOutputs_14_15_port, 
      MuxOutputs_14_14_port, MuxOutputs_14_13_port, MuxOutputs_14_12_port, 
      MuxOutputs_14_11_port, MuxOutputs_14_10_port, MuxOutputs_14_9_port, 
      MuxOutputs_14_8_port, MuxOutputs_14_7_port, MuxOutputs_14_6_port, 
      MuxOutputs_14_5_port, MuxOutputs_14_4_port, MuxOutputs_14_3_port, 
      MuxOutputs_14_2_port, MuxOutputs_14_1_port, MuxOutputs_14_0_port, 
      MuxOutputs_13_63_port, MuxOutputs_13_62_port, MuxOutputs_13_61_port, 
      MuxOutputs_13_60_port, MuxOutputs_13_59_port, MuxOutputs_13_58_port, 
      MuxOutputs_13_57_port, MuxOutputs_13_56_port, MuxOutputs_13_55_port, 
      MuxOutputs_13_54_port, MuxOutputs_13_53_port, MuxOutputs_13_52_port, 
      MuxOutputs_13_51_port, MuxOutputs_13_50_port, MuxOutputs_13_49_port, 
      MuxOutputs_13_48_port, MuxOutputs_13_47_port, MuxOutputs_13_46_port, 
      MuxOutputs_13_45_port, MuxOutputs_13_44_port, MuxOutputs_13_43_port, 
      MuxOutputs_13_42_port, MuxOutputs_13_41_port, MuxOutputs_13_40_port, 
      MuxOutputs_13_39_port, MuxOutputs_13_38_port, MuxOutputs_13_37_port, 
      MuxOutputs_13_36_port, MuxOutputs_13_35_port, MuxOutputs_13_34_port, 
      MuxOutputs_13_33_port, MuxOutputs_13_32_port, MuxOutputs_13_31_port, 
      MuxOutputs_13_30_port, MuxOutputs_13_29_port, MuxOutputs_13_28_port, 
      MuxOutputs_13_27_port, MuxOutputs_13_26_port, MuxOutputs_13_25_port, 
      MuxOutputs_13_24_port, MuxOutputs_13_23_port, MuxOutputs_13_22_port, 
      MuxOutputs_13_21_port, MuxOutputs_13_20_port, MuxOutputs_13_19_port, 
      MuxOutputs_13_18_port, MuxOutputs_13_17_port, MuxOutputs_13_16_port, 
      MuxOutputs_13_15_port, MuxOutputs_13_14_port, MuxOutputs_13_13_port, 
      MuxOutputs_13_12_port, MuxOutputs_13_11_port, MuxOutputs_13_10_port, 
      MuxOutputs_13_9_port, MuxOutputs_13_8_port, MuxOutputs_13_7_port, 
      MuxOutputs_13_6_port, MuxOutputs_13_5_port, MuxOutputs_13_4_port, 
      MuxOutputs_13_3_port, MuxOutputs_13_2_port, MuxOutputs_13_1_port, 
      MuxOutputs_13_0_port, MuxOutputs_12_63_port, MuxOutputs_12_62_port, 
      MuxOutputs_12_61_port, MuxOutputs_12_60_port, MuxOutputs_12_59_port, 
      MuxOutputs_12_58_port, MuxOutputs_12_57_port, MuxOutputs_12_56_port, 
      MuxOutputs_12_55_port, MuxOutputs_12_54_port, MuxOutputs_12_53_port, 
      MuxOutputs_12_52_port, MuxOutputs_12_51_port, MuxOutputs_12_50_port, 
      MuxOutputs_12_49_port, MuxOutputs_12_48_port, MuxOutputs_12_47_port, 
      MuxOutputs_12_46_port, MuxOutputs_12_45_port, MuxOutputs_12_44_port, 
      MuxOutputs_12_43_port, MuxOutputs_12_42_port, MuxOutputs_12_41_port, 
      MuxOutputs_12_40_port, MuxOutputs_12_39_port, MuxOutputs_12_38_port, 
      MuxOutputs_12_37_port, MuxOutputs_12_36_port, MuxOutputs_12_35_port, 
      MuxOutputs_12_34_port, MuxOutputs_12_33_port, MuxOutputs_12_32_port, 
      MuxOutputs_12_31_port, MuxOutputs_12_30_port, MuxOutputs_12_29_port, 
      MuxOutputs_12_28_port, MuxOutputs_12_27_port, MuxOutputs_12_26_port, 
      MuxOutputs_12_25_port, MuxOutputs_12_24_port, MuxOutputs_12_23_port, 
      MuxOutputs_12_22_port, MuxOutputs_12_21_port, MuxOutputs_12_20_port, 
      MuxOutputs_12_19_port, MuxOutputs_12_18_port, MuxOutputs_12_17_port, 
      MuxOutputs_12_16_port, MuxOutputs_12_15_port, MuxOutputs_12_14_port, 
      MuxOutputs_12_13_port, MuxOutputs_12_12_port, MuxOutputs_12_11_port, 
      MuxOutputs_12_10_port, MuxOutputs_12_9_port, MuxOutputs_12_8_port, 
      MuxOutputs_12_7_port, MuxOutputs_12_6_port, MuxOutputs_12_5_port, 
      MuxOutputs_12_4_port, MuxOutputs_12_3_port, MuxOutputs_12_2_port, 
      MuxOutputs_12_1_port, MuxOutputs_12_0_port, MuxOutputs_11_63_port, 
      MuxOutputs_11_62_port, MuxOutputs_11_61_port, MuxOutputs_11_60_port, 
      MuxOutputs_11_59_port, MuxOutputs_11_58_port, MuxOutputs_11_57_port, 
      MuxOutputs_11_56_port, MuxOutputs_11_55_port, MuxOutputs_11_54_port, 
      MuxOutputs_11_53_port, MuxOutputs_11_52_port, MuxOutputs_11_51_port, 
      MuxOutputs_11_50_port, MuxOutputs_11_49_port, MuxOutputs_11_48_port, 
      MuxOutputs_11_47_port, MuxOutputs_11_46_port, MuxOutputs_11_45_port, 
      MuxOutputs_11_44_port, MuxOutputs_11_43_port, MuxOutputs_11_42_port, 
      MuxOutputs_11_41_port, MuxOutputs_11_40_port, MuxOutputs_11_39_port, 
      MuxOutputs_11_38_port, MuxOutputs_11_37_port, MuxOutputs_11_36_port, 
      MuxOutputs_11_35_port, MuxOutputs_11_34_port, MuxOutputs_11_33_port, 
      MuxOutputs_11_32_port, MuxOutputs_11_31_port, MuxOutputs_11_30_port, 
      MuxOutputs_11_29_port, MuxOutputs_11_28_port, MuxOutputs_11_27_port, 
      MuxOutputs_11_26_port, MuxOutputs_11_25_port, MuxOutputs_11_24_port, 
      MuxOutputs_11_23_port, MuxOutputs_11_22_port, MuxOutputs_11_21_port, 
      MuxOutputs_11_20_port, MuxOutputs_11_19_port, MuxOutputs_11_18_port, 
      MuxOutputs_11_17_port, MuxOutputs_11_16_port, MuxOutputs_11_15_port, 
      MuxOutputs_11_14_port, MuxOutputs_11_13_port, MuxOutputs_11_12_port, 
      MuxOutputs_11_11_port, MuxOutputs_11_10_port, MuxOutputs_11_9_port, 
      MuxOutputs_11_8_port, MuxOutputs_11_7_port, MuxOutputs_11_6_port, 
      MuxOutputs_11_5_port, MuxOutputs_11_4_port, MuxOutputs_11_3_port, 
      MuxOutputs_11_2_port, MuxOutputs_11_1_port, MuxOutputs_11_0_port, 
      MuxOutputs_10_63_port, MuxOutputs_10_62_port, MuxOutputs_10_61_port, 
      MuxOutputs_10_60_port, MuxOutputs_10_59_port, MuxOutputs_10_58_port, 
      MuxOutputs_10_57_port, MuxOutputs_10_56_port, MuxOutputs_10_55_port, 
      MuxOutputs_10_54_port, MuxOutputs_10_53_port, MuxOutputs_10_52_port, 
      MuxOutputs_10_51_port, MuxOutputs_10_50_port, MuxOutputs_10_49_port, 
      MuxOutputs_10_48_port, MuxOutputs_10_47_port, MuxOutputs_10_46_port, 
      MuxOutputs_10_45_port, MuxOutputs_10_44_port, MuxOutputs_10_43_port, 
      MuxOutputs_10_42_port, MuxOutputs_10_41_port, MuxOutputs_10_40_port, 
      MuxOutputs_10_39_port, MuxOutputs_10_38_port, MuxOutputs_10_37_port, 
      MuxOutputs_10_36_port, MuxOutputs_10_35_port, MuxOutputs_10_34_port, 
      MuxOutputs_10_33_port, MuxOutputs_10_32_port, MuxOutputs_10_31_port, 
      MuxOutputs_10_30_port, MuxOutputs_10_29_port, MuxOutputs_10_28_port, 
      MuxOutputs_10_27_port, MuxOutputs_10_26_port, MuxOutputs_10_25_port, 
      MuxOutputs_10_24_port, MuxOutputs_10_23_port, MuxOutputs_10_22_port, 
      MuxOutputs_10_21_port, MuxOutputs_10_20_port, MuxOutputs_10_19_port, 
      MuxOutputs_10_18_port, MuxOutputs_10_17_port, MuxOutputs_10_16_port, 
      MuxOutputs_10_15_port, MuxOutputs_10_14_port, MuxOutputs_10_13_port, 
      MuxOutputs_10_12_port, MuxOutputs_10_11_port, MuxOutputs_10_10_port, 
      MuxOutputs_10_9_port, MuxOutputs_10_8_port, MuxOutputs_10_7_port, 
      MuxOutputs_10_6_port, MuxOutputs_10_5_port, MuxOutputs_10_4_port, 
      MuxOutputs_10_3_port, MuxOutputs_10_2_port, MuxOutputs_10_1_port, 
      MuxOutputs_10_0_port, MuxOutputs_9_63_port, MuxOutputs_9_62_port, 
      MuxOutputs_9_61_port, MuxOutputs_9_60_port, MuxOutputs_9_59_port, 
      MuxOutputs_9_58_port, MuxOutputs_9_57_port, MuxOutputs_9_56_port, 
      MuxOutputs_9_55_port, MuxOutputs_9_54_port, MuxOutputs_9_53_port, 
      MuxOutputs_9_52_port, MuxOutputs_9_51_port, MuxOutputs_9_50_port, 
      MuxOutputs_9_49_port, MuxOutputs_9_48_port, MuxOutputs_9_47_port, 
      MuxOutputs_9_46_port, MuxOutputs_9_45_port, MuxOutputs_9_44_port, 
      MuxOutputs_9_43_port, MuxOutputs_9_42_port, MuxOutputs_9_41_port, 
      MuxOutputs_9_40_port, MuxOutputs_9_39_port, MuxOutputs_9_38_port, 
      MuxOutputs_9_37_port, MuxOutputs_9_36_port, MuxOutputs_9_35_port, 
      MuxOutputs_9_34_port, MuxOutputs_9_33_port, MuxOutputs_9_32_port, 
      MuxOutputs_9_31_port, MuxOutputs_9_30_port, MuxOutputs_9_29_port, 
      MuxOutputs_9_28_port, MuxOutputs_9_27_port, MuxOutputs_9_26_port, 
      MuxOutputs_9_25_port, MuxOutputs_9_24_port, MuxOutputs_9_23_port, 
      MuxOutputs_9_22_port, MuxOutputs_9_21_port, MuxOutputs_9_20_port, 
      MuxOutputs_9_19_port, MuxOutputs_9_18_port, MuxOutputs_9_17_port, 
      MuxOutputs_9_16_port, MuxOutputs_9_15_port, MuxOutputs_9_14_port, 
      MuxOutputs_9_13_port, MuxOutputs_9_12_port, MuxOutputs_9_11_port, 
      MuxOutputs_9_10_port, MuxOutputs_9_9_port, MuxOutputs_9_8_port, 
      MuxOutputs_9_7_port, MuxOutputs_9_6_port, MuxOutputs_9_5_port, 
      MuxOutputs_9_4_port, MuxOutputs_9_3_port, MuxOutputs_9_2_port, 
      MuxOutputs_9_1_port, MuxOutputs_9_0_port, MuxOutputs_8_63_port, 
      MuxOutputs_8_62_port, MuxOutputs_8_61_port, MuxOutputs_8_60_port, 
      MuxOutputs_8_59_port, MuxOutputs_8_58_port, MuxOutputs_8_57_port, 
      MuxOutputs_8_56_port, MuxOutputs_8_55_port, MuxOutputs_8_54_port, 
      MuxOutputs_8_53_port, MuxOutputs_8_52_port, MuxOutputs_8_51_port, 
      MuxOutputs_8_50_port, MuxOutputs_8_49_port, MuxOutputs_8_48_port, 
      MuxOutputs_8_47_port, MuxOutputs_8_46_port, MuxOutputs_8_45_port, 
      MuxOutputs_8_44_port, MuxOutputs_8_43_port, MuxOutputs_8_42_port, 
      MuxOutputs_8_41_port, MuxOutputs_8_40_port, MuxOutputs_8_39_port, 
      MuxOutputs_8_38_port, MuxOutputs_8_37_port, MuxOutputs_8_36_port, 
      MuxOutputs_8_35_port, MuxOutputs_8_34_port, MuxOutputs_8_33_port, 
      MuxOutputs_8_32_port, MuxOutputs_8_31_port, MuxOutputs_8_30_port, 
      MuxOutputs_8_29_port, MuxOutputs_8_28_port, MuxOutputs_8_27_port, 
      MuxOutputs_8_26_port, MuxOutputs_8_25_port, MuxOutputs_8_24_port, 
      MuxOutputs_8_23_port, MuxOutputs_8_22_port, MuxOutputs_8_21_port, 
      MuxOutputs_8_20_port, MuxOutputs_8_19_port, MuxOutputs_8_18_port, 
      MuxOutputs_8_17_port, MuxOutputs_8_16_port, MuxOutputs_8_15_port, 
      MuxOutputs_8_14_port, MuxOutputs_8_13_port, MuxOutputs_8_12_port, 
      MuxOutputs_8_11_port, MuxOutputs_8_10_port, MuxOutputs_8_9_port, 
      MuxOutputs_8_8_port, MuxOutputs_8_7_port, MuxOutputs_8_6_port, 
      MuxOutputs_8_5_port, MuxOutputs_8_4_port, MuxOutputs_8_3_port, 
      MuxOutputs_8_2_port, MuxOutputs_8_1_port, MuxOutputs_8_0_port, 
      SumOutputs_7_63_port, SumOutputs_7_62_port, SumOutputs_7_61_port, 
      SumOutputs_7_60_port, SumOutputs_7_59_port, SumOutputs_7_58_port, 
      SumOutputs_7_57_port, SumOutputs_7_56_port, SumOutputs_7_55_port, 
      SumOutputs_7_54_port, SumOutputs_7_53_port, SumOutputs_7_52_port, 
      SumOutputs_7_51_port, SumOutputs_7_50_port, SumOutputs_7_49_port, 
      SumOutputs_7_48_port, SumOutputs_7_47_port, SumOutputs_7_46_port, 
      SumOutputs_7_45_port, SumOutputs_7_44_port, SumOutputs_7_43_port, 
      SumOutputs_7_42_port, SumOutputs_7_41_port, SumOutputs_7_40_port, 
      SumOutputs_7_39_port, SumOutputs_7_38_port, SumOutputs_7_37_port, 
      SumOutputs_7_36_port, SumOutputs_7_35_port, SumOutputs_7_34_port, 
      SumOutputs_7_33_port, SumOutputs_7_32_port, SumOutputs_7_31_port, 
      SumOutputs_7_30_port, SumOutputs_7_29_port, SumOutputs_7_28_port, 
      SumOutputs_7_27_port, SumOutputs_7_26_port, SumOutputs_7_25_port, 
      SumOutputs_7_24_port, SumOutputs_7_23_port, SumOutputs_7_22_port, 
      SumOutputs_7_21_port, SumOutputs_7_20_port, SumOutputs_7_19_port, 
      SumOutputs_7_18_port, SumOutputs_7_17_port, SumOutputs_7_16_port, 
      SumOutputs_7_15_port, SumOutputs_7_14_port, SumOutputs_7_13_port, 
      SumOutputs_7_12_port, SumOutputs_7_11_port, SumOutputs_7_10_port, 
      SumOutputs_7_9_port, SumOutputs_7_8_port, SumOutputs_7_7_port, 
      SumOutputs_7_6_port, SumOutputs_7_5_port, SumOutputs_7_4_port, 
      SumOutputs_7_3_port, SumOutputs_7_2_port, SumOutputs_7_1_port, 
      SumOutputs_7_0_port, SumOutputs_6_63_port, SumOutputs_6_62_port, 
      SumOutputs_6_61_port, SumOutputs_6_60_port, SumOutputs_6_59_port, 
      SumOutputs_6_58_port, SumOutputs_6_57_port, SumOutputs_6_56_port, 
      SumOutputs_6_55_port, SumOutputs_6_54_port, SumOutputs_6_53_port, 
      SumOutputs_6_52_port, SumOutputs_6_51_port, SumOutputs_6_50_port, 
      SumOutputs_6_49_port, SumOutputs_6_48_port, SumOutputs_6_47_port, 
      SumOutputs_6_46_port, SumOutputs_6_45_port, SumOutputs_6_44_port, 
      SumOutputs_6_43_port, SumOutputs_6_42_port, SumOutputs_6_41_port, 
      SumOutputs_6_40_port, SumOutputs_6_39_port, SumOutputs_6_38_port, 
      SumOutputs_6_37_port, SumOutputs_6_36_port, SumOutputs_6_35_port, 
      SumOutputs_6_34_port, SumOutputs_6_33_port, SumOutputs_6_32_port, 
      SumOutputs_6_31_port, SumOutputs_6_30_port, SumOutputs_6_29_port, 
      SumOutputs_6_28_port, SumOutputs_6_27_port, SumOutputs_6_26_port, 
      SumOutputs_6_25_port, SumOutputs_6_24_port, SumOutputs_6_23_port, 
      SumOutputs_6_22_port, SumOutputs_6_21_port, SumOutputs_6_20_port, 
      SumOutputs_6_19_port, SumOutputs_6_18_port, SumOutputs_6_17_port, 
      SumOutputs_6_16_port, SumOutputs_6_15_port, SumOutputs_6_14_port, 
      SumOutputs_6_13_port, SumOutputs_6_12_port, SumOutputs_6_11_port, 
      SumOutputs_6_10_port, SumOutputs_6_9_port, SumOutputs_6_8_port, 
      SumOutputs_6_7_port, SumOutputs_6_6_port, SumOutputs_6_5_port, 
      SumOutputs_6_4_port, SumOutputs_6_3_port, SumOutputs_6_2_port, 
      SumOutputs_6_1_port, SumOutputs_6_0_port, SumOutputs_5_63_port, 
      SumOutputs_5_62_port, SumOutputs_5_61_port, SumOutputs_5_60_port, 
      SumOutputs_5_59_port, SumOutputs_5_58_port, SumOutputs_5_57_port, 
      SumOutputs_5_56_port, SumOutputs_5_55_port, SumOutputs_5_54_port, 
      SumOutputs_5_53_port, SumOutputs_5_52_port, SumOutputs_5_51_port, 
      SumOutputs_5_50_port, SumOutputs_5_49_port, SumOutputs_5_48_port, 
      SumOutputs_5_47_port, SumOutputs_5_46_port, SumOutputs_5_45_port, 
      SumOutputs_5_44_port, SumOutputs_5_43_port, SumOutputs_5_42_port, 
      SumOutputs_5_41_port, SumOutputs_5_40_port, SumOutputs_5_39_port, 
      SumOutputs_5_38_port, SumOutputs_5_37_port, SumOutputs_5_36_port, 
      SumOutputs_5_35_port, SumOutputs_5_34_port, SumOutputs_5_33_port, 
      SumOutputs_5_32_port, SumOutputs_5_31_port, SumOutputs_5_30_port, 
      SumOutputs_5_29_port, SumOutputs_5_28_port, SumOutputs_5_27_port, 
      SumOutputs_5_26_port, SumOutputs_5_25_port, SumOutputs_5_24_port, 
      SumOutputs_5_23_port, SumOutputs_5_22_port, SumOutputs_5_21_port, 
      SumOutputs_5_20_port, SumOutputs_5_19_port, SumOutputs_5_18_port, 
      SumOutputs_5_17_port, SumOutputs_5_16_port, SumOutputs_5_15_port, 
      SumOutputs_5_14_port, SumOutputs_5_13_port, SumOutputs_5_12_port, 
      SumOutputs_5_11_port, SumOutputs_5_10_port, SumOutputs_5_9_port, 
      SumOutputs_5_8_port, SumOutputs_5_7_port, SumOutputs_5_6_port, 
      SumOutputs_5_5_port, SumOutputs_5_4_port, SumOutputs_5_3_port, 
      SumOutputs_5_2_port, SumOutputs_5_1_port, SumOutputs_5_0_port, 
      SumOutputs_4_63_port, SumOutputs_4_62_port, SumOutputs_4_61_port, 
      SumOutputs_4_60_port, SumOutputs_4_59_port, SumOutputs_4_58_port, 
      SumOutputs_4_57_port, SumOutputs_4_56_port, SumOutputs_4_55_port, 
      SumOutputs_4_54_port, SumOutputs_4_53_port, SumOutputs_4_52_port, 
      SumOutputs_4_51_port, SumOutputs_4_50_port, SumOutputs_4_49_port, 
      SumOutputs_4_48_port, SumOutputs_4_47_port, SumOutputs_4_46_port, 
      SumOutputs_4_45_port, SumOutputs_4_44_port, SumOutputs_4_43_port, 
      SumOutputs_4_42_port, SumOutputs_4_41_port, SumOutputs_4_40_port, 
      SumOutputs_4_39_port, SumOutputs_4_38_port, SumOutputs_4_37_port, 
      SumOutputs_4_36_port, SumOutputs_4_35_port, SumOutputs_4_34_port, 
      SumOutputs_4_33_port, SumOutputs_4_32_port, SumOutputs_4_31_port, 
      SumOutputs_4_30_port, SumOutputs_4_29_port, SumOutputs_4_28_port, 
      SumOutputs_4_27_port, SumOutputs_4_26_port, SumOutputs_4_25_port, 
      SumOutputs_4_24_port, SumOutputs_4_23_port, SumOutputs_4_22_port, 
      SumOutputs_4_21_port, SumOutputs_4_20_port, SumOutputs_4_19_port, 
      SumOutputs_4_18_port, SumOutputs_4_17_port, SumOutputs_4_16_port, 
      SumOutputs_4_15_port, SumOutputs_4_14_port, SumOutputs_4_13_port, 
      SumOutputs_4_12_port, SumOutputs_4_11_port, SumOutputs_4_10_port, 
      SumOutputs_4_9_port, SumOutputs_4_8_port, SumOutputs_4_7_port, 
      SumOutputs_4_6_port, SumOutputs_4_5_port, SumOutputs_4_4_port, 
      SumOutputs_4_3_port, SumOutputs_4_2_port, SumOutputs_4_1_port, 
      SumOutputs_4_0_port, SumOutputs_3_63_port, SumOutputs_3_62_port, 
      SumOutputs_3_61_port, SumOutputs_3_60_port, SumOutputs_3_59_port, 
      SumOutputs_3_58_port, SumOutputs_3_57_port, SumOutputs_3_56_port, 
      SumOutputs_3_55_port, SumOutputs_3_54_port, SumOutputs_3_53_port, 
      SumOutputs_3_52_port, SumOutputs_3_51_port, SumOutputs_3_50_port, 
      SumOutputs_3_49_port, SumOutputs_3_48_port, SumOutputs_3_47_port, 
      SumOutputs_3_46_port, SumOutputs_3_45_port, SumOutputs_3_44_port, 
      SumOutputs_3_43_port, SumOutputs_3_42_port, SumOutputs_3_41_port, 
      SumOutputs_3_40_port, SumOutputs_3_39_port, SumOutputs_3_38_port, 
      SumOutputs_3_37_port, SumOutputs_3_36_port, SumOutputs_3_35_port, 
      SumOutputs_3_34_port, SumOutputs_3_33_port, SumOutputs_3_32_port, 
      SumOutputs_3_31_port, SumOutputs_3_30_port, SumOutputs_3_29_port, 
      SumOutputs_3_28_port, SumOutputs_3_27_port, SumOutputs_3_26_port, 
      SumOutputs_3_25_port, SumOutputs_3_24_port, SumOutputs_3_23_port, 
      SumOutputs_3_22_port, SumOutputs_3_21_port, SumOutputs_3_20_port, 
      SumOutputs_3_19_port, SumOutputs_3_18_port, SumOutputs_3_17_port, 
      SumOutputs_3_16_port, SumOutputs_3_15_port, SumOutputs_3_14_port, 
      SumOutputs_3_13_port, SumOutputs_3_12_port, SumOutputs_3_11_port, 
      SumOutputs_3_10_port, SumOutputs_3_9_port, SumOutputs_3_8_port, 
      SumOutputs_3_7_port, SumOutputs_3_6_port, SumOutputs_3_5_port, 
      SumOutputs_3_4_port, SumOutputs_3_3_port, SumOutputs_3_2_port, 
      SumOutputs_3_1_port, SumOutputs_3_0_port, SumOutputs_2_63_port, 
      SumOutputs_2_62_port, SumOutputs_2_61_port, SumOutputs_2_60_port, 
      SumOutputs_2_59_port, SumOutputs_2_58_port, SumOutputs_2_57_port, 
      SumOutputs_2_56_port, SumOutputs_2_55_port, SumOutputs_2_54_port, 
      SumOutputs_2_53_port, SumOutputs_2_52_port, SumOutputs_2_51_port, 
      SumOutputs_2_50_port, SumOutputs_2_49_port, SumOutputs_2_48_port, 
      SumOutputs_2_47_port, SumOutputs_2_46_port, SumOutputs_2_45_port, 
      SumOutputs_2_44_port, SumOutputs_2_43_port, SumOutputs_2_42_port, 
      SumOutputs_2_41_port, SumOutputs_2_40_port, SumOutputs_2_39_port, 
      SumOutputs_2_38_port, SumOutputs_2_37_port, SumOutputs_2_36_port, 
      SumOutputs_2_35_port, SumOutputs_2_34_port, SumOutputs_2_33_port, 
      SumOutputs_2_32_port, SumOutputs_2_31_port, SumOutputs_2_30_port, 
      SumOutputs_2_29_port, SumOutputs_2_28_port, SumOutputs_2_27_port, 
      SumOutputs_2_26_port, SumOutputs_2_25_port, SumOutputs_2_24_port, 
      SumOutputs_2_23_port, SumOutputs_2_22_port, SumOutputs_2_21_port, 
      SumOutputs_2_20_port, SumOutputs_2_19_port, SumOutputs_2_18_port, 
      SumOutputs_2_17_port, SumOutputs_2_16_port, SumOutputs_2_15_port, 
      SumOutputs_2_14_port, SumOutputs_2_13_port, SumOutputs_2_12_port, 
      SumOutputs_2_11_port, SumOutputs_2_10_port, SumOutputs_2_9_port, 
      SumOutputs_2_8_port, SumOutputs_2_7_port, SumOutputs_2_6_port, 
      SumOutputs_2_5_port, SumOutputs_2_4_port, SumOutputs_2_3_port, 
      SumOutputs_2_2_port, SumOutputs_2_1_port, SumOutputs_2_0_port, 
      SumOutputs_1_63_port, SumOutputs_1_62_port, SumOutputs_1_61_port, 
      SumOutputs_1_60_port, SumOutputs_1_59_port, SumOutputs_1_58_port, 
      SumOutputs_1_57_port, SumOutputs_1_56_port, SumOutputs_1_55_port, 
      SumOutputs_1_54_port, SumOutputs_1_53_port, SumOutputs_1_52_port, 
      SumOutputs_1_51_port, SumOutputs_1_50_port, SumOutputs_1_49_port, 
      SumOutputs_1_48_port, SumOutputs_1_47_port, SumOutputs_1_46_port, 
      SumOutputs_1_45_port, SumOutputs_1_44_port, SumOutputs_1_43_port, 
      SumOutputs_1_42_port, SumOutputs_1_41_port, SumOutputs_1_40_port, 
      SumOutputs_1_39_port, SumOutputs_1_38_port, SumOutputs_1_37_port, 
      SumOutputs_1_36_port, SumOutputs_1_35_port, SumOutputs_1_34_port, 
      SumOutputs_1_33_port, SumOutputs_1_32_port, SumOutputs_1_31_port, 
      SumOutputs_1_30_port, SumOutputs_1_29_port, SumOutputs_1_28_port, 
      SumOutputs_1_27_port, SumOutputs_1_26_port, SumOutputs_1_25_port, 
      SumOutputs_1_24_port, SumOutputs_1_23_port, SumOutputs_1_22_port, 
      SumOutputs_1_21_port, SumOutputs_1_20_port, SumOutputs_1_19_port, 
      SumOutputs_1_18_port, SumOutputs_1_17_port, SumOutputs_1_16_port, 
      SumOutputs_1_15_port, SumOutputs_1_14_port, SumOutputs_1_13_port, 
      SumOutputs_1_12_port, SumOutputs_1_11_port, SumOutputs_1_10_port, 
      SumOutputs_1_9_port, SumOutputs_1_8_port, SumOutputs_1_7_port, 
      SumOutputs_1_6_port, SumOutputs_1_5_port, SumOutputs_1_4_port, 
      SumOutputs_1_3_port, SumOutputs_1_2_port, SumOutputs_1_1_port, 
      SumOutputs_1_0_port, SumOutputs_0_63_port, SumOutputs_0_62_port, 
      SumOutputs_0_61_port, SumOutputs_0_60_port, SumOutputs_0_59_port, 
      SumOutputs_0_58_port, SumOutputs_0_57_port, SumOutputs_0_56_port, 
      SumOutputs_0_55_port, SumOutputs_0_54_port, SumOutputs_0_53_port, 
      SumOutputs_0_52_port, SumOutputs_0_51_port, SumOutputs_0_50_port, 
      SumOutputs_0_49_port, SumOutputs_0_48_port, SumOutputs_0_47_port, 
      SumOutputs_0_46_port, SumOutputs_0_45_port, SumOutputs_0_44_port, 
      SumOutputs_0_43_port, SumOutputs_0_42_port, SumOutputs_0_41_port, 
      SumOutputs_0_40_port, SumOutputs_0_39_port, SumOutputs_0_38_port, 
      SumOutputs_0_37_port, SumOutputs_0_36_port, SumOutputs_0_35_port, 
      SumOutputs_0_34_port, SumOutputs_0_33_port, SumOutputs_0_32_port, 
      SumOutputs_0_31_port, SumOutputs_0_30_port, SumOutputs_0_29_port, 
      SumOutputs_0_28_port, SumOutputs_0_27_port, SumOutputs_0_26_port, 
      SumOutputs_0_25_port, SumOutputs_0_24_port, SumOutputs_0_23_port, 
      SumOutputs_0_22_port, SumOutputs_0_21_port, SumOutputs_0_20_port, 
      SumOutputs_0_19_port, SumOutputs_0_18_port, SumOutputs_0_17_port, 
      SumOutputs_0_16_port, SumOutputs_0_15_port, SumOutputs_0_14_port, 
      SumOutputs_0_13_port, SumOutputs_0_12_port, SumOutputs_0_11_port, 
      SumOutputs_0_10_port, SumOutputs_0_9_port, SumOutputs_0_8_port, 
      SumOutputs_0_7_port, SumOutputs_0_6_port, SumOutputs_0_5_port, 
      SumOutputs_0_4_port, SumOutputs_0_3_port, SumOutputs_0_2_port, 
      SumOutputs_0_1_port, SumOutputs_0_0_port, SumOutputs_13_63_port, 
      SumOutputs_13_62_port, SumOutputs_13_61_port, SumOutputs_13_60_port, 
      SumOutputs_13_59_port, SumOutputs_13_58_port, SumOutputs_13_57_port, 
      SumOutputs_13_56_port, SumOutputs_13_55_port, SumOutputs_13_54_port, 
      SumOutputs_13_53_port, SumOutputs_13_52_port, SumOutputs_13_51_port, 
      SumOutputs_13_50_port, SumOutputs_13_49_port, SumOutputs_13_48_port, 
      SumOutputs_13_47_port, SumOutputs_13_46_port, SumOutputs_13_45_port, 
      SumOutputs_13_44_port, SumOutputs_13_43_port, SumOutputs_13_42_port, 
      SumOutputs_13_41_port, SumOutputs_13_40_port, SumOutputs_13_39_port, 
      SumOutputs_13_38_port, SumOutputs_13_37_port, SumOutputs_13_36_port, 
      SumOutputs_13_35_port, SumOutputs_13_34_port, SumOutputs_13_33_port, 
      SumOutputs_13_32_port, SumOutputs_13_31_port, SumOutputs_13_30_port, 
      SumOutputs_13_29_port, SumOutputs_13_28_port, SumOutputs_13_27_port, 
      SumOutputs_13_26_port, SumOutputs_13_25_port, SumOutputs_13_24_port, 
      SumOutputs_13_23_port, SumOutputs_13_22_port, SumOutputs_13_21_port, 
      SumOutputs_13_20_port, SumOutputs_13_19_port, SumOutputs_13_18_port, 
      SumOutputs_13_17_port, SumOutputs_13_16_port, SumOutputs_13_15_port, 
      SumOutputs_13_14_port, SumOutputs_13_13_port, SumOutputs_13_12_port, 
      SumOutputs_13_11_port, SumOutputs_13_10_port, SumOutputs_13_9_port, 
      SumOutputs_13_8_port, SumOutputs_13_7_port, SumOutputs_13_6_port, 
      SumOutputs_13_5_port, SumOutputs_13_4_port, SumOutputs_13_3_port, 
      SumOutputs_13_2_port, SumOutputs_13_1_port, SumOutputs_13_0_port, 
      SumOutputs_12_63_port, SumOutputs_12_62_port, SumOutputs_12_61_port, 
      SumOutputs_12_60_port, SumOutputs_12_59_port, SumOutputs_12_58_port, 
      SumOutputs_12_57_port, SumOutputs_12_56_port, SumOutputs_12_55_port, 
      SumOutputs_12_54_port, SumOutputs_12_53_port, SumOutputs_12_52_port, 
      SumOutputs_12_51_port, SumOutputs_12_50_port, SumOutputs_12_49_port, 
      SumOutputs_12_48_port, SumOutputs_12_47_port, SumOutputs_12_46_port, 
      SumOutputs_12_45_port, SumOutputs_12_44_port, SumOutputs_12_43_port, 
      SumOutputs_12_42_port, SumOutputs_12_41_port, SumOutputs_12_40_port, 
      SumOutputs_12_39_port, SumOutputs_12_38_port, SumOutputs_12_37_port, 
      SumOutputs_12_36_port, SumOutputs_12_35_port, SumOutputs_12_34_port, 
      SumOutputs_12_33_port, SumOutputs_12_32_port, SumOutputs_12_31_port, 
      SumOutputs_12_30_port, SumOutputs_12_29_port, SumOutputs_12_28_port, 
      SumOutputs_12_27_port, SumOutputs_12_26_port, SumOutputs_12_25_port, 
      SumOutputs_12_24_port, SumOutputs_12_23_port, SumOutputs_12_22_port, 
      SumOutputs_12_21_port, SumOutputs_12_20_port, SumOutputs_12_19_port, 
      SumOutputs_12_18_port, SumOutputs_12_17_port, SumOutputs_12_16_port, 
      SumOutputs_12_15_port, SumOutputs_12_14_port, SumOutputs_12_13_port, 
      SumOutputs_12_12_port, SumOutputs_12_11_port, SumOutputs_12_10_port, 
      SumOutputs_12_9_port, SumOutputs_12_8_port, SumOutputs_12_7_port, 
      SumOutputs_12_6_port, SumOutputs_12_5_port, SumOutputs_12_4_port, 
      SumOutputs_12_3_port, SumOutputs_12_2_port, SumOutputs_12_1_port, 
      SumOutputs_12_0_port, SumOutputs_11_63_port, SumOutputs_11_62_port, 
      SumOutputs_11_61_port, SumOutputs_11_60_port, SumOutputs_11_59_port, 
      SumOutputs_11_58_port, SumOutputs_11_57_port, SumOutputs_11_56_port, 
      SumOutputs_11_55_port, SumOutputs_11_54_port, SumOutputs_11_53_port, 
      SumOutputs_11_52_port, SumOutputs_11_51_port, SumOutputs_11_50_port, 
      SumOutputs_11_49_port, SumOutputs_11_48_port, SumOutputs_11_47_port, 
      SumOutputs_11_46_port, SumOutputs_11_45_port, SumOutputs_11_44_port, 
      SumOutputs_11_43_port, SumOutputs_11_42_port, SumOutputs_11_41_port, 
      SumOutputs_11_40_port, SumOutputs_11_39_port, SumOutputs_11_38_port, 
      SumOutputs_11_37_port, SumOutputs_11_36_port, SumOutputs_11_35_port, 
      SumOutputs_11_34_port, SumOutputs_11_33_port, SumOutputs_11_32_port, 
      SumOutputs_11_31_port, SumOutputs_11_30_port, SumOutputs_11_29_port, 
      SumOutputs_11_28_port, SumOutputs_11_27_port, SumOutputs_11_26_port, 
      SumOutputs_11_25_port, SumOutputs_11_24_port, SumOutputs_11_23_port, 
      SumOutputs_11_22_port, SumOutputs_11_21_port, SumOutputs_11_20_port, 
      SumOutputs_11_19_port, SumOutputs_11_18_port, SumOutputs_11_17_port, 
      SumOutputs_11_16_port, SumOutputs_11_15_port, SumOutputs_11_14_port, 
      SumOutputs_11_13_port, SumOutputs_11_12_port, SumOutputs_11_11_port, 
      SumOutputs_11_10_port, SumOutputs_11_9_port, SumOutputs_11_8_port, 
      SumOutputs_11_7_port, SumOutputs_11_6_port, SumOutputs_11_5_port, 
      SumOutputs_11_4_port, SumOutputs_11_3_port, SumOutputs_11_2_port, 
      SumOutputs_11_1_port, SumOutputs_11_0_port, SumOutputs_10_63_port, 
      SumOutputs_10_62_port, SumOutputs_10_61_port, SumOutputs_10_60_port, 
      SumOutputs_10_59_port, SumOutputs_10_58_port, SumOutputs_10_57_port, 
      SumOutputs_10_56_port, SumOutputs_10_55_port, SumOutputs_10_54_port, 
      SumOutputs_10_53_port, SumOutputs_10_52_port, SumOutputs_10_51_port, 
      SumOutputs_10_50_port, SumOutputs_10_49_port, SumOutputs_10_48_port, 
      SumOutputs_10_47_port, SumOutputs_10_46_port, SumOutputs_10_45_port, 
      SumOutputs_10_44_port, SumOutputs_10_43_port, SumOutputs_10_42_port, 
      SumOutputs_10_41_port, SumOutputs_10_40_port, SumOutputs_10_39_port, 
      SumOutputs_10_38_port, SumOutputs_10_37_port, SumOutputs_10_36_port, 
      SumOutputs_10_35_port, SumOutputs_10_34_port, SumOutputs_10_33_port, 
      SumOutputs_10_32_port, SumOutputs_10_31_port, SumOutputs_10_30_port, 
      SumOutputs_10_29_port, SumOutputs_10_28_port, SumOutputs_10_27_port, 
      SumOutputs_10_26_port, SumOutputs_10_25_port, SumOutputs_10_24_port, 
      SumOutputs_10_23_port, SumOutputs_10_22_port, SumOutputs_10_21_port, 
      SumOutputs_10_20_port, SumOutputs_10_19_port, SumOutputs_10_18_port, 
      SumOutputs_10_17_port, SumOutputs_10_16_port, SumOutputs_10_15_port, 
      SumOutputs_10_14_port, SumOutputs_10_13_port, SumOutputs_10_12_port, 
      SumOutputs_10_11_port, SumOutputs_10_10_port, SumOutputs_10_9_port, 
      SumOutputs_10_8_port, SumOutputs_10_7_port, SumOutputs_10_6_port, 
      SumOutputs_10_5_port, SumOutputs_10_4_port, SumOutputs_10_3_port, 
      SumOutputs_10_2_port, SumOutputs_10_1_port, SumOutputs_10_0_port, 
      SumOutputs_9_63_port, SumOutputs_9_62_port, SumOutputs_9_61_port, 
      SumOutputs_9_60_port, SumOutputs_9_59_port, SumOutputs_9_58_port, 
      SumOutputs_9_57_port, SumOutputs_9_56_port, SumOutputs_9_55_port, 
      SumOutputs_9_54_port, SumOutputs_9_53_port, SumOutputs_9_52_port, 
      SumOutputs_9_51_port, SumOutputs_9_50_port, SumOutputs_9_49_port, 
      SumOutputs_9_48_port, SumOutputs_9_47_port, SumOutputs_9_46_port, 
      SumOutputs_9_45_port, SumOutputs_9_44_port, SumOutputs_9_43_port, 
      SumOutputs_9_42_port, SumOutputs_9_41_port, SumOutputs_9_40_port, 
      SumOutputs_9_39_port, SumOutputs_9_38_port, SumOutputs_9_37_port, 
      SumOutputs_9_36_port, SumOutputs_9_35_port, SumOutputs_9_34_port, 
      SumOutputs_9_33_port, SumOutputs_9_32_port, SumOutputs_9_31_port, 
      SumOutputs_9_30_port, SumOutputs_9_29_port, SumOutputs_9_28_port, 
      SumOutputs_9_27_port, SumOutputs_9_26_port, SumOutputs_9_25_port, 
      SumOutputs_9_24_port, SumOutputs_9_23_port, SumOutputs_9_22_port, 
      SumOutputs_9_21_port, SumOutputs_9_20_port, SumOutputs_9_19_port, 
      SumOutputs_9_18_port, SumOutputs_9_17_port, SumOutputs_9_16_port, 
      SumOutputs_9_15_port, SumOutputs_9_14_port, SumOutputs_9_13_port, 
      SumOutputs_9_12_port, SumOutputs_9_11_port, SumOutputs_9_10_port, 
      SumOutputs_9_9_port, SumOutputs_9_8_port, SumOutputs_9_7_port, 
      SumOutputs_9_6_port, SumOutputs_9_5_port, SumOutputs_9_4_port, 
      SumOutputs_9_3_port, SumOutputs_9_2_port, SumOutputs_9_1_port, 
      SumOutputs_9_0_port, SumOutputs_8_63_port, SumOutputs_8_62_port, 
      SumOutputs_8_61_port, SumOutputs_8_60_port, SumOutputs_8_59_port, 
      SumOutputs_8_58_port, SumOutputs_8_57_port, SumOutputs_8_56_port, 
      SumOutputs_8_55_port, SumOutputs_8_54_port, SumOutputs_8_53_port, 
      SumOutputs_8_52_port, SumOutputs_8_51_port, SumOutputs_8_50_port, 
      SumOutputs_8_49_port, SumOutputs_8_48_port, SumOutputs_8_47_port, 
      SumOutputs_8_46_port, SumOutputs_8_45_port, SumOutputs_8_44_port, 
      SumOutputs_8_43_port, SumOutputs_8_42_port, SumOutputs_8_41_port, 
      SumOutputs_8_40_port, SumOutputs_8_39_port, SumOutputs_8_38_port, 
      SumOutputs_8_37_port, SumOutputs_8_36_port, SumOutputs_8_35_port, 
      SumOutputs_8_34_port, SumOutputs_8_33_port, SumOutputs_8_32_port, 
      SumOutputs_8_31_port, SumOutputs_8_30_port, SumOutputs_8_29_port, 
      SumOutputs_8_28_port, SumOutputs_8_27_port, SumOutputs_8_26_port, 
      SumOutputs_8_25_port, SumOutputs_8_24_port, SumOutputs_8_23_port, 
      SumOutputs_8_22_port, SumOutputs_8_21_port, SumOutputs_8_20_port, 
      SumOutputs_8_19_port, SumOutputs_8_18_port, SumOutputs_8_17_port, 
      SumOutputs_8_16_port, SumOutputs_8_15_port, SumOutputs_8_14_port, 
      SumOutputs_8_13_port, SumOutputs_8_12_port, SumOutputs_8_11_port, 
      SumOutputs_8_10_port, SumOutputs_8_9_port, SumOutputs_8_8_port, 
      SumOutputs_8_7_port, SumOutputs_8_6_port, SumOutputs_8_5_port, 
      SumOutputs_8_4_port, SumOutputs_8_3_port, SumOutputs_8_2_port, 
      SumOutputs_8_1_port, SumOutputs_8_0_port, n8, n9, n10, n11, n12, n13, n14
      , n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, 
      n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43
      , n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, 
      n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72
      , n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, 
      n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, 
      n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, 
      n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, 
      n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, 
      n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, 
      n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, 
      n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, 
      n173, n174, n175, n176, n177, n178, n179, n180, n181, n_1000, n_1001, 
      n_1002, n_1003, n_1004, n_1005, n_1006, n_1007, n_1008, n_1009, n_1010, 
      n_1011, n_1012, n_1013, n_1014, n_1015, n_1016, n_1017, n_1018, n_1019, 
      n_1020, n_1021, n_1022, n_1023, n_1024, n_1025, n_1026, n_1027, n_1028, 
      n_1029, n_1030, n_1031, n_1032, n_1033, n_1034, n_1035, n_1036, n_1037, 
      n_1038, n_1039, n_1040, n_1041, n_1042, n_1043, n_1044, n_1045, n_1046, 
      n_1047, n_1048, n_1049, n_1050, n_1051, n_1052, n_1053, n_1054, n_1055, 
      n_1056, n_1057, n_1058, n_1059, n_1060, n_1061, n_1062, n_1063, n_1064, 
      n_1065, n_1066, n_1067, n_1068, n_1069, n_1070, n_1071, n_1072, n_1073, 
      n_1074, n_1075, n_1076, n_1077, n_1078, n_1079, n_1080, n_1081, n_1082, 
      n_1083, n_1084, n_1085, n_1086, n_1087, n_1088, n_1089, n_1090, n_1091, 
      n_1092, n_1093, n_1094, n_1095, n_1096, n_1097, n_1098, n_1099, n_1100, 
      n_1101, n_1102, n_1103, n_1104, n_1105, n_1106, n_1107, n_1108, n_1109, 
      n_1110, n_1111, n_1112, n_1113, n_1114, n_1115, n_1116, n_1117, n_1118, 
      n_1119, n_1120, n_1121, n_1122, n_1123, n_1124, n_1125, n_1126, n_1127, 
      n_1128, n_1129, n_1130, n_1131, n_1132, n_1133, n_1134, n_1135, n_1136, 
      n_1137, n_1138, n_1139, n_1140, n_1141 : std_logic;

begin
   
   inverterI_0 : IV_64 port map( A => A(0), Y => A_complement_0_port);
   inverterI_1 : IV_127 port map( A => A(1), Y => A_complement_1_port);
   inverterI_2 : IV_126 port map( A => A(2), Y => A_complement_2_port);
   inverterI_3 : IV_125 port map( A => A(3), Y => A_complement_3_port);
   inverterI_4 : IV_124 port map( A => A(4), Y => A_complement_4_port);
   inverterI_5 : IV_123 port map( A => A(5), Y => A_complement_5_port);
   inverterI_6 : IV_122 port map( A => A(6), Y => A_complement_6_port);
   inverterI_7 : IV_121 port map( A => A(7), Y => A_complement_7_port);
   inverterI_8 : IV_120 port map( A => A(8), Y => A_complement_8_port);
   inverterI_9 : IV_119 port map( A => A(9), Y => A_complement_9_port);
   inverterI_10 : IV_118 port map( A => A(10), Y => A_complement_10_port);
   inverterI_11 : IV_117 port map( A => A(11), Y => A_complement_11_port);
   inverterI_12 : IV_116 port map( A => A(12), Y => A_complement_12_port);
   inverterI_13 : IV_115 port map( A => A(13), Y => A_complement_13_port);
   inverterI_14 : IV_114 port map( A => A(14), Y => A_complement_14_port);
   inverterI_15 : IV_113 port map( A => A(15), Y => A_complement_15_port);
   inverterI_16 : IV_112 port map( A => A(16), Y => A_complement_16_port);
   inverterI_17 : IV_111 port map( A => A(17), Y => A_complement_17_port);
   inverterI_18 : IV_110 port map( A => A(18), Y => A_complement_18_port);
   inverterI_19 : IV_109 port map( A => A(19), Y => A_complement_19_port);
   inverterI_20 : IV_108 port map( A => A(20), Y => A_complement_20_port);
   inverterI_21 : IV_107 port map( A => A(21), Y => A_complement_21_port);
   inverterI_22 : IV_106 port map( A => A(22), Y => A_complement_22_port);
   inverterI_23 : IV_105 port map( A => A(23), Y => A_complement_23_port);
   inverterI_24 : IV_104 port map( A => A(24), Y => A_complement_24_port);
   inverterI_25 : IV_103 port map( A => A(25), Y => A_complement_25_port);
   inverterI_26 : IV_102 port map( A => A(26), Y => A_complement_26_port);
   inverterI_27 : IV_101 port map( A => A(27), Y => A_complement_27_port);
   inverterI_28 : IV_100 port map( A => A(28), Y => A_complement_28_port);
   inverterI_29 : IV_99 port map( A => A(29), Y => A_complement_29_port);
   inverterI_30 : IV_98 port map( A => A(30), Y => A_complement_30_port);
   inverterI_31 : IV_97 port map( A => A(31), Y => A_complement_31_port);
   inverterI_32 : IV_96 port map( A => A(31), Y => A_complement_32_port);
   inverterI_33 : IV_95 port map( A => A(31), Y => A_complement_33_port);
   inverterI_34 : IV_94 port map( A => A(31), Y => A_complement_34_port);
   inverterI_35 : IV_93 port map( A => A(31), Y => A_complement_35_port);
   inverterI_36 : IV_92 port map( A => A(31), Y => A_complement_36_port);
   inverterI_37 : IV_91 port map( A => A(31), Y => A_complement_37_port);
   inverterI_38 : IV_90 port map( A => A(31), Y => A_complement_38_port);
   inverterI_39 : IV_89 port map( A => A(31), Y => A_complement_39_port);
   inverterI_40 : IV_88 port map( A => A(31), Y => A_complement_40_port);
   inverterI_41 : IV_87 port map( A => A(31), Y => A_complement_41_port);
   inverterI_42 : IV_86 port map( A => A(31), Y => A_complement_42_port);
   inverterI_43 : IV_85 port map( A => A(31), Y => A_complement_43_port);
   inverterI_44 : IV_84 port map( A => A(31), Y => A_complement_44_port);
   inverterI_45 : IV_83 port map( A => A(31), Y => A_complement_45_port);
   inverterI_46 : IV_82 port map( A => A(31), Y => A_complement_46_port);
   inverterI_47 : IV_81 port map( A => A(31), Y => A_complement_47_port);
   inverterI_48 : IV_80 port map( A => A(31), Y => A_complement_48_port);
   inverterI_49 : IV_79 port map( A => A(31), Y => A_complement_49_port);
   inverterI_50 : IV_78 port map( A => A(31), Y => A_complement_50_port);
   inverterI_51 : IV_77 port map( A => A(31), Y => A_complement_51_port);
   inverterI_52 : IV_76 port map( A => A(31), Y => A_complement_52_port);
   inverterI_53 : IV_75 port map( A => A(31), Y => A_complement_53_port);
   inverterI_54 : IV_74 port map( A => A(31), Y => A_complement_54_port);
   inverterI_55 : IV_73 port map( A => A(31), Y => A_complement_55_port);
   inverterI_56 : IV_72 port map( A => A(31), Y => A_complement_56_port);
   inverterI_57 : IV_71 port map( A => A(31), Y => A_complement_57_port);
   inverterI_58 : IV_70 port map( A => A(31), Y => A_complement_58_port);
   inverterI_59 : IV_69 port map( A => A(31), Y => A_complement_59_port);
   inverterI_60 : IV_68 port map( A => A(31), Y => A_complement_60_port);
   inverterI_61 : IV_67 port map( A => A(31), Y => A_complement_61_port);
   inverterI_62 : IV_66 port map( A => A(31), Y => A_complement_62_port);
   inverterI_63 : IV_65 port map( A => A(31), Y => A_complement_63_port);
   FinilizingNegativeSignal : RCA_NbitRca64_16 port map( A(63) => 
                           A_complement_63_port, A(62) => A_complement_62_port,
                           A(61) => A_complement_61_port, A(60) => 
                           A_complement_60_port, A(59) => A_complement_59_port,
                           A(58) => A_complement_58_port, A(57) => 
                           A_complement_57_port, A(56) => A_complement_56_port,
                           A(55) => A_complement_55_port, A(54) => 
                           A_complement_54_port, A(53) => A_complement_53_port,
                           A(52) => A_complement_52_port, A(51) => 
                           A_complement_51_port, A(50) => A_complement_50_port,
                           A(49) => A_complement_49_port, A(48) => 
                           A_complement_48_port, A(47) => A_complement_47_port,
                           A(46) => A_complement_46_port, A(45) => 
                           A_complement_45_port, A(44) => A_complement_44_port,
                           A(43) => A_complement_43_port, A(42) => 
                           A_complement_42_port, A(41) => A_complement_41_port,
                           A(40) => A_complement_40_port, A(39) => 
                           A_complement_39_port, A(38) => A_complement_38_port,
                           A(37) => A_complement_37_port, A(36) => 
                           A_complement_36_port, A(35) => A_complement_35_port,
                           A(34) => A_complement_34_port, A(33) => 
                           A_complement_33_port, A(32) => A_complement_32_port,
                           A(31) => A_complement_31_port, A(30) => 
                           A_complement_30_port, A(29) => A_complement_29_port,
                           A(28) => A_complement_28_port, A(27) => 
                           A_complement_27_port, A(26) => A_complement_26_port,
                           A(25) => A_complement_25_port, A(24) => 
                           A_complement_24_port, A(23) => A_complement_23_port,
                           A(22) => A_complement_22_port, A(21) => 
                           A_complement_21_port, A(20) => A_complement_20_port,
                           A(19) => A_complement_19_port, A(18) => 
                           A_complement_18_port, A(17) => A_complement_17_port,
                           A(16) => A_complement_16_port, A(15) => 
                           A_complement_15_port, A(14) => A_complement_14_port,
                           A(13) => A_complement_13_port, A(12) => 
                           A_complement_12_port, A(11) => A_complement_11_port,
                           A(10) => A_complement_10_port, A(9) => 
                           A_complement_9_port, A(8) => A_complement_8_port, 
                           A(7) => A_complement_7_port, A(6) => 
                           A_complement_6_port, A(5) => A_complement_5_port, 
                           A(4) => A_complement_4_port, A(3) => 
                           A_complement_3_port, A(2) => A_complement_2_port, 
                           A(1) => A_complement_1_port, A(0) => 
                           A_complement_0_port, B(63) => X_Logic0_port, B(62) 
                           => X_Logic0_port, B(61) => X_Logic0_port, B(60) => 
                           X_Logic0_port, B(59) => X_Logic0_port, B(58) => 
                           X_Logic0_port, B(57) => X_Logic0_port, B(56) => 
                           X_Logic0_port, B(55) => X_Logic0_port, B(54) => 
                           X_Logic0_port, B(53) => X_Logic0_port, B(52) => 
                           X_Logic0_port, B(51) => X_Logic0_port, B(50) => 
                           X_Logic0_port, B(49) => X_Logic0_port, B(48) => 
                           X_Logic0_port, B(47) => X_Logic0_port, B(46) => 
                           X_Logic0_port, B(45) => X_Logic0_port, B(44) => 
                           X_Logic0_port, B(43) => X_Logic0_port, B(42) => 
                           X_Logic0_port, B(41) => X_Logic0_port, B(40) => 
                           X_Logic0_port, B(39) => X_Logic0_port, B(38) => 
                           X_Logic0_port, B(37) => X_Logic0_port, B(36) => 
                           X_Logic0_port, B(35) => X_Logic0_port, B(34) => 
                           X_Logic0_port, B(33) => X_Logic0_port, B(32) => 
                           X_Logic0_port, B(31) => X_Logic0_port, B(30) => 
                           X_Logic0_port, B(29) => X_Logic0_port, B(28) => 
                           X_Logic0_port, B(27) => X_Logic0_port, B(26) => 
                           X_Logic0_port, B(25) => X_Logic0_port, B(24) => 
                           X_Logic0_port, B(23) => X_Logic0_port, B(22) => 
                           X_Logic0_port, B(21) => X_Logic0_port, B(20) => 
                           X_Logic0_port, B(19) => X_Logic0_port, B(18) => 
                           X_Logic0_port, B(17) => X_Logic0_port, B(16) => 
                           X_Logic0_port, B(15) => X_Logic0_port, B(14) => 
                           X_Logic0_port, B(13) => X_Logic0_port, B(12) => 
                           X_Logic0_port, B(11) => X_Logic0_port, B(10) => 
                           X_Logic0_port, B(9) => X_Logic0_port, B(8) => 
                           X_Logic0_port, B(7) => X_Logic0_port, B(6) => 
                           X_Logic0_port, B(5) => X_Logic0_port, B(4) => 
                           X_Logic0_port, B(3) => X_Logic0_port, B(2) => 
                           X_Logic0_port, B(1) => X_Logic0_port, B(0) => 
                           X_Logic0_port, Ci => X_Logic1_port, S(63) => 
                           negative_inputs_0_63_port, S(62) => 
                           negative_inputs_0_62_port, S(61) => 
                           negative_inputs_0_61_port, S(60) => 
                           negative_inputs_0_60_port, S(59) => 
                           negative_inputs_0_59_port, S(58) => 
                           negative_inputs_0_58_port, S(57) => 
                           negative_inputs_0_57_port, S(56) => 
                           negative_inputs_0_56_port, S(55) => 
                           negative_inputs_0_55_port, S(54) => 
                           negative_inputs_0_54_port, S(53) => 
                           negative_inputs_0_53_port, S(52) => 
                           negative_inputs_0_52_port, S(51) => 
                           negative_inputs_0_51_port, S(50) => 
                           negative_inputs_0_50_port, S(49) => 
                           negative_inputs_0_49_port, S(48) => 
                           negative_inputs_0_48_port, S(47) => 
                           negative_inputs_0_47_port, S(46) => 
                           negative_inputs_0_46_port, S(45) => 
                           negative_inputs_0_45_port, S(44) => 
                           negative_inputs_0_44_port, S(43) => 
                           negative_inputs_0_43_port, S(42) => 
                           negative_inputs_0_42_port, S(41) => 
                           negative_inputs_0_41_port, S(40) => 
                           negative_inputs_0_40_port, S(39) => 
                           negative_inputs_0_39_port, S(38) => 
                           negative_inputs_0_38_port, S(37) => 
                           negative_inputs_0_37_port, S(36) => 
                           negative_inputs_0_36_port, S(35) => 
                           negative_inputs_0_35_port, S(34) => 
                           negative_inputs_0_34_port, S(33) => 
                           negative_inputs_0_33_port, S(32) => 
                           negative_inputs_0_32_port, S(31) => 
                           negative_inputs_0_31_port, S(30) => 
                           negative_inputs_0_30_port, S(29) => 
                           negative_inputs_0_29_port, S(28) => 
                           negative_inputs_0_28_port, S(27) => 
                           negative_inputs_0_27_port, S(26) => 
                           negative_inputs_0_26_port, S(25) => 
                           negative_inputs_0_25_port, S(24) => 
                           negative_inputs_0_24_port, S(23) => 
                           negative_inputs_0_23_port, S(22) => 
                           negative_inputs_0_22_port, S(21) => 
                           negative_inputs_0_21_port, S(20) => 
                           negative_inputs_0_20_port, S(19) => 
                           negative_inputs_0_19_port, S(18) => 
                           negative_inputs_0_18_port, S(17) => 
                           negative_inputs_0_17_port, S(16) => 
                           negative_inputs_0_16_port, S(15) => 
                           negative_inputs_0_15_port, S(14) => 
                           negative_inputs_0_14_port, S(13) => 
                           negative_inputs_0_13_port, S(12) => 
                           negative_inputs_0_12_port, S(11) => 
                           negative_inputs_0_11_port, S(10) => 
                           negative_inputs_0_10_port, S(9) => 
                           negative_inputs_0_9_port, S(8) => 
                           negative_inputs_0_8_port, S(7) => 
                           negative_inputs_0_7_port, S(6) => 
                           negative_inputs_0_6_port, S(5) => 
                           negative_inputs_0_5_port, S(4) => 
                           negative_inputs_0_4_port, S(3) => 
                           negative_inputs_0_3_port, S(2) => 
                           negative_inputs_0_2_port, S(1) => 
                           negative_inputs_0_1_port, S(0) => 
                           negative_inputs_0_0_port, Co => n_1000);
   shifted_pos_1 : leftshifter_NbitShifter64_63 port map( shift_in(63) => A(31)
                           , shift_in(62) => A(31), shift_in(61) => A(31), 
                           shift_in(60) => A(31), shift_in(59) => A(31), 
                           shift_in(58) => A(31), shift_in(57) => A(31), 
                           shift_in(56) => A(31), shift_in(55) => A(31), 
                           shift_in(54) => A(31), shift_in(53) => A(31), 
                           shift_in(52) => A(31), shift_in(51) => A(31), 
                           shift_in(50) => A(31), shift_in(49) => A(31), 
                           shift_in(48) => A(31), shift_in(47) => A(31), 
                           shift_in(46) => A(31), shift_in(45) => A(31), 
                           shift_in(44) => A(31), shift_in(43) => A(31), 
                           shift_in(42) => A(31), shift_in(41) => A(31), 
                           shift_in(40) => A(31), shift_in(39) => A(31), 
                           shift_in(38) => A(31), shift_in(37) => A(31), 
                           shift_in(36) => A(31), shift_in(35) => A(31), 
                           shift_in(34) => A(31), shift_in(33) => A(31), 
                           shift_in(32) => A(31), shift_in(31) => A(31), 
                           shift_in(30) => A(30), shift_in(29) => A(29), 
                           shift_in(28) => A(28), shift_in(27) => A(27), 
                           shift_in(26) => A(26), shift_in(25) => A(25), 
                           shift_in(24) => A(24), shift_in(23) => A(23), 
                           shift_in(22) => A(22), shift_in(21) => A(21), 
                           shift_in(20) => A(20), shift_in(19) => A(19), 
                           shift_in(18) => A(18), shift_in(17) => A(17), 
                           shift_in(16) => A(16), shift_in(15) => A(15), 
                           shift_in(14) => A(14), shift_in(13) => A(13), 
                           shift_in(12) => A(12), shift_in(11) => A(11), 
                           shift_in(10) => A(10), shift_in(9) => A(9), 
                           shift_in(8) => A(8), shift_in(7) => A(7), 
                           shift_in(6) => A(6), shift_in(5) => A(5), 
                           shift_in(4) => A(4), shift_in(3) => A(3), 
                           shift_in(2) => A(2), shift_in(1) => n15, shift_in(0)
                           => n18, shift_out(63) => positive_inputs_1_63_port, 
                           shift_out(62) => positive_inputs_1_62_port, 
                           shift_out(61) => positive_inputs_1_61_port, 
                           shift_out(60) => positive_inputs_1_60_port, 
                           shift_out(59) => positive_inputs_1_59_port, 
                           shift_out(58) => positive_inputs_1_58_port, 
                           shift_out(57) => positive_inputs_1_57_port, 
                           shift_out(56) => positive_inputs_1_56_port, 
                           shift_out(55) => positive_inputs_1_55_port, 
                           shift_out(54) => positive_inputs_1_54_port, 
                           shift_out(53) => positive_inputs_1_53_port, 
                           shift_out(52) => positive_inputs_1_52_port, 
                           shift_out(51) => positive_inputs_1_51_port, 
                           shift_out(50) => positive_inputs_1_50_port, 
                           shift_out(49) => positive_inputs_1_49_port, 
                           shift_out(48) => positive_inputs_1_48_port, 
                           shift_out(47) => positive_inputs_1_47_port, 
                           shift_out(46) => positive_inputs_1_46_port, 
                           shift_out(45) => positive_inputs_1_45_port, 
                           shift_out(44) => positive_inputs_1_44_port, 
                           shift_out(43) => positive_inputs_1_43_port, 
                           shift_out(42) => positive_inputs_1_42_port, 
                           shift_out(41) => positive_inputs_1_41_port, 
                           shift_out(40) => positive_inputs_1_40_port, 
                           shift_out(39) => positive_inputs_1_39_port, 
                           shift_out(38) => positive_inputs_1_38_port, 
                           shift_out(37) => positive_inputs_1_37_port, 
                           shift_out(36) => positive_inputs_1_36_port, 
                           shift_out(35) => positive_inputs_1_35_port, 
                           shift_out(34) => positive_inputs_1_34_port, 
                           shift_out(33) => positive_inputs_1_33_port, 
                           shift_out(32) => positive_inputs_1_32_port, 
                           shift_out(31) => positive_inputs_1_31_port, 
                           shift_out(30) => positive_inputs_1_30_port, 
                           shift_out(29) => positive_inputs_1_29_port, 
                           shift_out(28) => positive_inputs_1_28_port, 
                           shift_out(27) => positive_inputs_1_27_port, 
                           shift_out(26) => positive_inputs_1_26_port, 
                           shift_out(25) => positive_inputs_1_25_port, 
                           shift_out(24) => positive_inputs_1_24_port, 
                           shift_out(23) => positive_inputs_1_23_port, 
                           shift_out(22) => positive_inputs_1_22_port, 
                           shift_out(21) => positive_inputs_1_21_port, 
                           shift_out(20) => positive_inputs_1_20_port, 
                           shift_out(19) => positive_inputs_1_19_port, 
                           shift_out(18) => positive_inputs_1_18_port, 
                           shift_out(17) => positive_inputs_1_17_port, 
                           shift_out(16) => positive_inputs_1_16_port, 
                           shift_out(15) => positive_inputs_1_15_port, 
                           shift_out(14) => positive_inputs_1_14_port, 
                           shift_out(13) => positive_inputs_1_13_port, 
                           shift_out(12) => positive_inputs_1_12_port, 
                           shift_out(11) => positive_inputs_1_11_port, 
                           shift_out(10) => positive_inputs_1_10_port, 
                           shift_out(9) => positive_inputs_1_9_port, 
                           shift_out(8) => positive_inputs_1_8_port, 
                           shift_out(7) => positive_inputs_1_7_port, 
                           shift_out(6) => positive_inputs_1_6_port, 
                           shift_out(5) => positive_inputs_1_5_port, 
                           shift_out(4) => positive_inputs_1_4_port, 
                           shift_out(3) => positive_inputs_1_3_port, 
                           shift_out(2) => positive_inputs_1_2_port, 
                           shift_out(1) => positive_inputs_1_1_port, 
                           shift_out(0) => n_1001);
   shifted_pos_2 : leftshifter_NbitShifter64_125 port map( shift_in(63) => 
                           positive_inputs_1_63_port, shift_in(62) => 
                           positive_inputs_1_62_port, shift_in(61) => 
                           positive_inputs_1_61_port, shift_in(60) => 
                           positive_inputs_1_60_port, shift_in(59) => 
                           positive_inputs_1_59_port, shift_in(58) => 
                           positive_inputs_1_58_port, shift_in(57) => 
                           positive_inputs_1_57_port, shift_in(56) => 
                           positive_inputs_1_56_port, shift_in(55) => 
                           positive_inputs_1_55_port, shift_in(54) => 
                           positive_inputs_1_54_port, shift_in(53) => 
                           positive_inputs_1_53_port, shift_in(52) => 
                           positive_inputs_1_52_port, shift_in(51) => 
                           positive_inputs_1_51_port, shift_in(50) => 
                           positive_inputs_1_50_port, shift_in(49) => 
                           positive_inputs_1_49_port, shift_in(48) => 
                           positive_inputs_1_48_port, shift_in(47) => 
                           positive_inputs_1_47_port, shift_in(46) => 
                           positive_inputs_1_46_port, shift_in(45) => 
                           positive_inputs_1_45_port, shift_in(44) => 
                           positive_inputs_1_44_port, shift_in(43) => 
                           positive_inputs_1_43_port, shift_in(42) => 
                           positive_inputs_1_42_port, shift_in(41) => 
                           positive_inputs_1_41_port, shift_in(40) => 
                           positive_inputs_1_40_port, shift_in(39) => 
                           positive_inputs_1_39_port, shift_in(38) => 
                           positive_inputs_1_38_port, shift_in(37) => n24, 
                           shift_in(36) => positive_inputs_1_36_port, 
                           shift_in(35) => positive_inputs_1_35_port, 
                           shift_in(34) => positive_inputs_1_34_port, 
                           shift_in(33) => positive_inputs_1_33_port, 
                           shift_in(32) => positive_inputs_1_32_port, 
                           shift_in(31) => positive_inputs_1_31_port, 
                           shift_in(30) => positive_inputs_1_30_port, 
                           shift_in(29) => positive_inputs_1_29_port, 
                           shift_in(28) => positive_inputs_1_28_port, 
                           shift_in(27) => positive_inputs_1_27_port, 
                           shift_in(26) => positive_inputs_1_26_port, 
                           shift_in(25) => positive_inputs_1_25_port, 
                           shift_in(24) => positive_inputs_1_24_port, 
                           shift_in(23) => positive_inputs_1_23_port, 
                           shift_in(22) => positive_inputs_1_22_port, 
                           shift_in(21) => positive_inputs_1_21_port, 
                           shift_in(20) => positive_inputs_1_20_port, 
                           shift_in(19) => positive_inputs_1_19_port, 
                           shift_in(18) => positive_inputs_1_18_port, 
                           shift_in(17) => positive_inputs_1_17_port, 
                           shift_in(16) => positive_inputs_1_16_port, 
                           shift_in(15) => positive_inputs_1_15_port, 
                           shift_in(14) => positive_inputs_1_14_port, 
                           shift_in(13) => positive_inputs_1_13_port, 
                           shift_in(12) => positive_inputs_1_12_port, 
                           shift_in(11) => positive_inputs_1_11_port, 
                           shift_in(10) => positive_inputs_1_10_port, 
                           shift_in(9) => positive_inputs_1_9_port, shift_in(8)
                           => positive_inputs_1_8_port, shift_in(7) => 
                           positive_inputs_1_7_port, shift_in(6) => 
                           positive_inputs_1_6_port, shift_in(5) => 
                           positive_inputs_1_5_port, shift_in(4) => 
                           positive_inputs_1_4_port, shift_in(3) => 
                           positive_inputs_1_3_port, shift_in(2) => 
                           positive_inputs_1_2_port, shift_in(1) => 
                           positive_inputs_1_1_port, shift_in(0) => n8, 
                           shift_out(63) => positive_inputs_2_63_port, 
                           shift_out(62) => positive_inputs_2_62_port, 
                           shift_out(61) => positive_inputs_2_61_port, 
                           shift_out(60) => positive_inputs_2_60_port, 
                           shift_out(59) => positive_inputs_2_59_port, 
                           shift_out(58) => positive_inputs_2_58_port, 
                           shift_out(57) => positive_inputs_2_57_port, 
                           shift_out(56) => positive_inputs_2_56_port, 
                           shift_out(55) => positive_inputs_2_55_port, 
                           shift_out(54) => positive_inputs_2_54_port, 
                           shift_out(53) => positive_inputs_2_53_port, 
                           shift_out(52) => positive_inputs_2_52_port, 
                           shift_out(51) => positive_inputs_2_51_port, 
                           shift_out(50) => positive_inputs_2_50_port, 
                           shift_out(49) => positive_inputs_2_49_port, 
                           shift_out(48) => positive_inputs_2_48_port, 
                           shift_out(47) => positive_inputs_2_47_port, 
                           shift_out(46) => positive_inputs_2_46_port, 
                           shift_out(45) => positive_inputs_2_45_port, 
                           shift_out(44) => positive_inputs_2_44_port, 
                           shift_out(43) => positive_inputs_2_43_port, 
                           shift_out(42) => positive_inputs_2_42_port, 
                           shift_out(41) => positive_inputs_2_41_port, 
                           shift_out(40) => positive_inputs_2_40_port, 
                           shift_out(39) => positive_inputs_2_39_port, 
                           shift_out(38) => positive_inputs_2_38_port, 
                           shift_out(37) => positive_inputs_2_37_port, 
                           shift_out(36) => positive_inputs_2_36_port, 
                           shift_out(35) => positive_inputs_2_35_port, 
                           shift_out(34) => positive_inputs_2_34_port, 
                           shift_out(33) => positive_inputs_2_33_port, 
                           shift_out(32) => positive_inputs_2_32_port, 
                           shift_out(31) => positive_inputs_2_31_port, 
                           shift_out(30) => positive_inputs_2_30_port, 
                           shift_out(29) => positive_inputs_2_29_port, 
                           shift_out(28) => positive_inputs_2_28_port, 
                           shift_out(27) => positive_inputs_2_27_port, 
                           shift_out(26) => positive_inputs_2_26_port, 
                           shift_out(25) => positive_inputs_2_25_port, 
                           shift_out(24) => positive_inputs_2_24_port, 
                           shift_out(23) => positive_inputs_2_23_port, 
                           shift_out(22) => positive_inputs_2_22_port, 
                           shift_out(21) => positive_inputs_2_21_port, 
                           shift_out(20) => positive_inputs_2_20_port, 
                           shift_out(19) => positive_inputs_2_19_port, 
                           shift_out(18) => positive_inputs_2_18_port, 
                           shift_out(17) => positive_inputs_2_17_port, 
                           shift_out(16) => positive_inputs_2_16_port, 
                           shift_out(15) => positive_inputs_2_15_port, 
                           shift_out(14) => positive_inputs_2_14_port, 
                           shift_out(13) => positive_inputs_2_13_port, 
                           shift_out(12) => positive_inputs_2_12_port, 
                           shift_out(11) => positive_inputs_2_11_port, 
                           shift_out(10) => positive_inputs_2_10_port, 
                           shift_out(9) => positive_inputs_2_9_port, 
                           shift_out(8) => positive_inputs_2_8_port, 
                           shift_out(7) => positive_inputs_2_7_port, 
                           shift_out(6) => positive_inputs_2_6_port, 
                           shift_out(5) => positive_inputs_2_5_port, 
                           shift_out(4) => positive_inputs_2_4_port, 
                           shift_out(3) => positive_inputs_2_3_port, 
                           shift_out(2) => positive_inputs_2_2_port, 
                           shift_out(1) => positive_inputs_2_1_port, 
                           shift_out(0) => n_1002);
   shifted_pos_3 : leftshifter_NbitShifter64_124 port map( shift_in(63) => 
                           positive_inputs_2_63_port, shift_in(62) => 
                           positive_inputs_2_62_port, shift_in(61) => 
                           positive_inputs_2_61_port, shift_in(60) => 
                           positive_inputs_2_60_port, shift_in(59) => 
                           positive_inputs_2_59_port, shift_in(58) => 
                           positive_inputs_2_58_port, shift_in(57) => 
                           positive_inputs_2_57_port, shift_in(56) => 
                           positive_inputs_2_56_port, shift_in(55) => 
                           positive_inputs_2_55_port, shift_in(54) => 
                           positive_inputs_2_54_port, shift_in(53) => 
                           positive_inputs_2_53_port, shift_in(52) => 
                           positive_inputs_2_52_port, shift_in(51) => 
                           positive_inputs_2_51_port, shift_in(50) => 
                           positive_inputs_2_50_port, shift_in(49) => 
                           positive_inputs_2_49_port, shift_in(48) => 
                           positive_inputs_2_48_port, shift_in(47) => n38, 
                           shift_in(46) => positive_inputs_2_46_port, 
                           shift_in(45) => positive_inputs_2_45_port, 
                           shift_in(44) => positive_inputs_2_44_port, 
                           shift_in(43) => positive_inputs_2_43_port, 
                           shift_in(42) => positive_inputs_2_42_port, 
                           shift_in(41) => positive_inputs_2_41_port, 
                           shift_in(40) => positive_inputs_2_40_port, 
                           shift_in(39) => positive_inputs_2_39_port, 
                           shift_in(38) => positive_inputs_2_38_port, 
                           shift_in(37) => n23, shift_in(36) => 
                           positive_inputs_2_36_port, shift_in(35) => 
                           positive_inputs_2_35_port, shift_in(34) => 
                           positive_inputs_2_34_port, shift_in(33) => 
                           positive_inputs_2_33_port, shift_in(32) => 
                           positive_inputs_2_32_port, shift_in(31) => 
                           positive_inputs_2_31_port, shift_in(30) => 
                           positive_inputs_2_30_port, shift_in(29) => 
                           positive_inputs_2_29_port, shift_in(28) => 
                           positive_inputs_2_28_port, shift_in(27) => 
                           positive_inputs_2_27_port, shift_in(26) => 
                           positive_inputs_2_26_port, shift_in(25) => 
                           positive_inputs_2_25_port, shift_in(24) => 
                           positive_inputs_2_24_port, shift_in(23) => 
                           positive_inputs_2_23_port, shift_in(22) => 
                           positive_inputs_2_22_port, shift_in(21) => 
                           positive_inputs_2_21_port, shift_in(20) => 
                           positive_inputs_2_20_port, shift_in(19) => 
                           positive_inputs_2_19_port, shift_in(18) => 
                           positive_inputs_2_18_port, shift_in(17) => 
                           positive_inputs_2_17_port, shift_in(16) => 
                           positive_inputs_2_16_port, shift_in(15) => 
                           positive_inputs_2_15_port, shift_in(14) => 
                           positive_inputs_2_14_port, shift_in(13) => 
                           positive_inputs_2_13_port, shift_in(12) => 
                           positive_inputs_2_12_port, shift_in(11) => 
                           positive_inputs_2_11_port, shift_in(10) => 
                           positive_inputs_2_10_port, shift_in(9) => 
                           positive_inputs_2_9_port, shift_in(8) => 
                           positive_inputs_2_8_port, shift_in(7) => 
                           positive_inputs_2_7_port, shift_in(6) => 
                           positive_inputs_2_6_port, shift_in(5) => 
                           positive_inputs_2_5_port, shift_in(4) => 
                           positive_inputs_2_4_port, shift_in(3) => 
                           positive_inputs_2_3_port, shift_in(2) => 
                           positive_inputs_2_2_port, shift_in(1) => 
                           positive_inputs_2_1_port, shift_in(0) => n8, 
                           shift_out(63) => positive_inputs_3_63_port, 
                           shift_out(62) => positive_inputs_3_62_port, 
                           shift_out(61) => positive_inputs_3_61_port, 
                           shift_out(60) => positive_inputs_3_60_port, 
                           shift_out(59) => positive_inputs_3_59_port, 
                           shift_out(58) => positive_inputs_3_58_port, 
                           shift_out(57) => positive_inputs_3_57_port, 
                           shift_out(56) => positive_inputs_3_56_port, 
                           shift_out(55) => positive_inputs_3_55_port, 
                           shift_out(54) => positive_inputs_3_54_port, 
                           shift_out(53) => positive_inputs_3_53_port, 
                           shift_out(52) => positive_inputs_3_52_port, 
                           shift_out(51) => positive_inputs_3_51_port, 
                           shift_out(50) => positive_inputs_3_50_port, 
                           shift_out(49) => positive_inputs_3_49_port, 
                           shift_out(48) => positive_inputs_3_48_port, 
                           shift_out(47) => positive_inputs_3_47_port, 
                           shift_out(46) => positive_inputs_3_46_port, 
                           shift_out(45) => positive_inputs_3_45_port, 
                           shift_out(44) => positive_inputs_3_44_port, 
                           shift_out(43) => positive_inputs_3_43_port, 
                           shift_out(42) => positive_inputs_3_42_port, 
                           shift_out(41) => positive_inputs_3_41_port, 
                           shift_out(40) => positive_inputs_3_40_port, 
                           shift_out(39) => positive_inputs_3_39_port, 
                           shift_out(38) => positive_inputs_3_38_port, 
                           shift_out(37) => positive_inputs_3_37_port, 
                           shift_out(36) => positive_inputs_3_36_port, 
                           shift_out(35) => positive_inputs_3_35_port, 
                           shift_out(34) => positive_inputs_3_34_port, 
                           shift_out(33) => positive_inputs_3_33_port, 
                           shift_out(32) => positive_inputs_3_32_port, 
                           shift_out(31) => positive_inputs_3_31_port, 
                           shift_out(30) => positive_inputs_3_30_port, 
                           shift_out(29) => positive_inputs_3_29_port, 
                           shift_out(28) => positive_inputs_3_28_port, 
                           shift_out(27) => positive_inputs_3_27_port, 
                           shift_out(26) => positive_inputs_3_26_port, 
                           shift_out(25) => positive_inputs_3_25_port, 
                           shift_out(24) => positive_inputs_3_24_port, 
                           shift_out(23) => positive_inputs_3_23_port, 
                           shift_out(22) => positive_inputs_3_22_port, 
                           shift_out(21) => positive_inputs_3_21_port, 
                           shift_out(20) => positive_inputs_3_20_port, 
                           shift_out(19) => positive_inputs_3_19_port, 
                           shift_out(18) => positive_inputs_3_18_port, 
                           shift_out(17) => positive_inputs_3_17_port, 
                           shift_out(16) => positive_inputs_3_16_port, 
                           shift_out(15) => positive_inputs_3_15_port, 
                           shift_out(14) => positive_inputs_3_14_port, 
                           shift_out(13) => positive_inputs_3_13_port, 
                           shift_out(12) => positive_inputs_3_12_port, 
                           shift_out(11) => positive_inputs_3_11_port, 
                           shift_out(10) => positive_inputs_3_10_port, 
                           shift_out(9) => positive_inputs_3_9_port, 
                           shift_out(8) => positive_inputs_3_8_port, 
                           shift_out(7) => positive_inputs_3_7_port, 
                           shift_out(6) => positive_inputs_3_6_port, 
                           shift_out(5) => positive_inputs_3_5_port, 
                           shift_out(4) => positive_inputs_3_4_port, 
                           shift_out(3) => positive_inputs_3_3_port, 
                           shift_out(2) => positive_inputs_3_2_port, 
                           shift_out(1) => positive_inputs_3_1_port, 
                           shift_out(0) => n_1003);
   shifted_pos_4 : leftshifter_NbitShifter64_123 port map( shift_in(63) => 
                           positive_inputs_3_63_port, shift_in(62) => 
                           positive_inputs_3_62_port, shift_in(61) => 
                           positive_inputs_3_61_port, shift_in(60) => 
                           positive_inputs_3_60_port, shift_in(59) => 
                           positive_inputs_3_59_port, shift_in(58) => 
                           positive_inputs_3_58_port, shift_in(57) => 
                           positive_inputs_3_57_port, shift_in(56) => 
                           positive_inputs_3_56_port, shift_in(55) => 
                           positive_inputs_3_55_port, shift_in(54) => 
                           positive_inputs_3_54_port, shift_in(53) => 
                           positive_inputs_3_53_port, shift_in(52) => 
                           positive_inputs_3_52_port, shift_in(51) => 
                           positive_inputs_3_51_port, shift_in(50) => 
                           positive_inputs_3_50_port, shift_in(49) => 
                           positive_inputs_3_49_port, shift_in(48) => 
                           positive_inputs_3_48_port, shift_in(47) => 
                           positive_inputs_3_47_port, shift_in(46) => 
                           positive_inputs_3_46_port, shift_in(45) => 
                           positive_inputs_3_45_port, shift_in(44) => 
                           positive_inputs_3_44_port, shift_in(43) => 
                           positive_inputs_3_43_port, shift_in(42) => 
                           positive_inputs_3_42_port, shift_in(41) => 
                           positive_inputs_3_41_port, shift_in(40) => 
                           positive_inputs_3_40_port, shift_in(39) => 
                           positive_inputs_3_39_port, shift_in(38) => 
                           positive_inputs_3_38_port, shift_in(37) => n22, 
                           shift_in(36) => positive_inputs_3_36_port, 
                           shift_in(35) => positive_inputs_3_35_port, 
                           shift_in(34) => positive_inputs_3_34_port, 
                           shift_in(33) => positive_inputs_3_33_port, 
                           shift_in(32) => positive_inputs_3_32_port, 
                           shift_in(31) => positive_inputs_3_31_port, 
                           shift_in(30) => positive_inputs_3_30_port, 
                           shift_in(29) => positive_inputs_3_29_port, 
                           shift_in(28) => positive_inputs_3_28_port, 
                           shift_in(27) => positive_inputs_3_27_port, 
                           shift_in(26) => positive_inputs_3_26_port, 
                           shift_in(25) => positive_inputs_3_25_port, 
                           shift_in(24) => positive_inputs_3_24_port, 
                           shift_in(23) => positive_inputs_3_23_port, 
                           shift_in(22) => positive_inputs_3_22_port, 
                           shift_in(21) => positive_inputs_3_21_port, 
                           shift_in(20) => positive_inputs_3_20_port, 
                           shift_in(19) => positive_inputs_3_19_port, 
                           shift_in(18) => positive_inputs_3_18_port, 
                           shift_in(17) => positive_inputs_3_17_port, 
                           shift_in(16) => positive_inputs_3_16_port, 
                           shift_in(15) => positive_inputs_3_15_port, 
                           shift_in(14) => positive_inputs_3_14_port, 
                           shift_in(13) => positive_inputs_3_13_port, 
                           shift_in(12) => positive_inputs_3_12_port, 
                           shift_in(11) => positive_inputs_3_11_port, 
                           shift_in(10) => positive_inputs_3_10_port, 
                           shift_in(9) => positive_inputs_3_9_port, shift_in(8)
                           => positive_inputs_3_8_port, shift_in(7) => 
                           positive_inputs_3_7_port, shift_in(6) => 
                           positive_inputs_3_6_port, shift_in(5) => 
                           positive_inputs_3_5_port, shift_in(4) => 
                           positive_inputs_3_4_port, shift_in(3) => 
                           positive_inputs_3_3_port, shift_in(2) => 
                           positive_inputs_3_2_port, shift_in(1) => 
                           positive_inputs_3_1_port, shift_in(0) => n8, 
                           shift_out(63) => positive_inputs_4_63_port, 
                           shift_out(62) => positive_inputs_4_62_port, 
                           shift_out(61) => positive_inputs_4_61_port, 
                           shift_out(60) => positive_inputs_4_60_port, 
                           shift_out(59) => positive_inputs_4_59_port, 
                           shift_out(58) => positive_inputs_4_58_port, 
                           shift_out(57) => positive_inputs_4_57_port, 
                           shift_out(56) => positive_inputs_4_56_port, 
                           shift_out(55) => positive_inputs_4_55_port, 
                           shift_out(54) => positive_inputs_4_54_port, 
                           shift_out(53) => positive_inputs_4_53_port, 
                           shift_out(52) => positive_inputs_4_52_port, 
                           shift_out(51) => positive_inputs_4_51_port, 
                           shift_out(50) => positive_inputs_4_50_port, 
                           shift_out(49) => positive_inputs_4_49_port, 
                           shift_out(48) => positive_inputs_4_48_port, 
                           shift_out(47) => positive_inputs_4_47_port, 
                           shift_out(46) => positive_inputs_4_46_port, 
                           shift_out(45) => positive_inputs_4_45_port, 
                           shift_out(44) => positive_inputs_4_44_port, 
                           shift_out(43) => positive_inputs_4_43_port, 
                           shift_out(42) => positive_inputs_4_42_port, 
                           shift_out(41) => positive_inputs_4_41_port, 
                           shift_out(40) => positive_inputs_4_40_port, 
                           shift_out(39) => positive_inputs_4_39_port, 
                           shift_out(38) => positive_inputs_4_38_port, 
                           shift_out(37) => positive_inputs_4_37_port, 
                           shift_out(36) => positive_inputs_4_36_port, 
                           shift_out(35) => positive_inputs_4_35_port, 
                           shift_out(34) => positive_inputs_4_34_port, 
                           shift_out(33) => positive_inputs_4_33_port, 
                           shift_out(32) => positive_inputs_4_32_port, 
                           shift_out(31) => positive_inputs_4_31_port, 
                           shift_out(30) => positive_inputs_4_30_port, 
                           shift_out(29) => positive_inputs_4_29_port, 
                           shift_out(28) => positive_inputs_4_28_port, 
                           shift_out(27) => positive_inputs_4_27_port, 
                           shift_out(26) => positive_inputs_4_26_port, 
                           shift_out(25) => positive_inputs_4_25_port, 
                           shift_out(24) => positive_inputs_4_24_port, 
                           shift_out(23) => positive_inputs_4_23_port, 
                           shift_out(22) => positive_inputs_4_22_port, 
                           shift_out(21) => positive_inputs_4_21_port, 
                           shift_out(20) => positive_inputs_4_20_port, 
                           shift_out(19) => positive_inputs_4_19_port, 
                           shift_out(18) => positive_inputs_4_18_port, 
                           shift_out(17) => positive_inputs_4_17_port, 
                           shift_out(16) => positive_inputs_4_16_port, 
                           shift_out(15) => positive_inputs_4_15_port, 
                           shift_out(14) => positive_inputs_4_14_port, 
                           shift_out(13) => positive_inputs_4_13_port, 
                           shift_out(12) => positive_inputs_4_12_port, 
                           shift_out(11) => positive_inputs_4_11_port, 
                           shift_out(10) => positive_inputs_4_10_port, 
                           shift_out(9) => positive_inputs_4_9_port, 
                           shift_out(8) => positive_inputs_4_8_port, 
                           shift_out(7) => positive_inputs_4_7_port, 
                           shift_out(6) => positive_inputs_4_6_port, 
                           shift_out(5) => positive_inputs_4_5_port, 
                           shift_out(4) => positive_inputs_4_4_port, 
                           shift_out(3) => positive_inputs_4_3_port, 
                           shift_out(2) => positive_inputs_4_2_port, 
                           shift_out(1) => positive_inputs_4_1_port, 
                           shift_out(0) => n_1004);
   shifted_pos_5 : leftshifter_NbitShifter64_122 port map( shift_in(63) => 
                           positive_inputs_4_63_port, shift_in(62) => 
                           positive_inputs_4_62_port, shift_in(61) => 
                           positive_inputs_4_61_port, shift_in(60) => 
                           positive_inputs_4_60_port, shift_in(59) => 
                           positive_inputs_4_59_port, shift_in(58) => 
                           positive_inputs_4_58_port, shift_in(57) => 
                           positive_inputs_4_57_port, shift_in(56) => 
                           positive_inputs_4_56_port, shift_in(55) => 
                           positive_inputs_4_55_port, shift_in(54) => 
                           positive_inputs_4_54_port, shift_in(53) => 
                           positive_inputs_4_53_port, shift_in(52) => 
                           positive_inputs_4_52_port, shift_in(51) => 
                           positive_inputs_4_51_port, shift_in(50) => 
                           positive_inputs_4_50_port, shift_in(49) => 
                           positive_inputs_4_49_port, shift_in(48) => 
                           positive_inputs_4_48_port, shift_in(47) => n37, 
                           shift_in(46) => positive_inputs_4_46_port, 
                           shift_in(45) => positive_inputs_4_45_port, 
                           shift_in(44) => positive_inputs_4_44_port, 
                           shift_in(43) => positive_inputs_4_43_port, 
                           shift_in(42) => positive_inputs_4_42_port, 
                           shift_in(41) => positive_inputs_4_41_port, 
                           shift_in(40) => positive_inputs_4_40_port, 
                           shift_in(39) => positive_inputs_4_39_port, 
                           shift_in(38) => positive_inputs_4_38_port, 
                           shift_in(37) => n21, shift_in(36) => 
                           positive_inputs_4_36_port, shift_in(35) => 
                           positive_inputs_4_35_port, shift_in(34) => 
                           positive_inputs_4_34_port, shift_in(33) => 
                           positive_inputs_4_33_port, shift_in(32) => 
                           positive_inputs_4_32_port, shift_in(31) => 
                           positive_inputs_4_31_port, shift_in(30) => 
                           positive_inputs_4_30_port, shift_in(29) => 
                           positive_inputs_4_29_port, shift_in(28) => 
                           positive_inputs_4_28_port, shift_in(27) => 
                           positive_inputs_4_27_port, shift_in(26) => 
                           positive_inputs_4_26_port, shift_in(25) => 
                           positive_inputs_4_25_port, shift_in(24) => 
                           positive_inputs_4_24_port, shift_in(23) => 
                           positive_inputs_4_23_port, shift_in(22) => 
                           positive_inputs_4_22_port, shift_in(21) => 
                           positive_inputs_4_21_port, shift_in(20) => 
                           positive_inputs_4_20_port, shift_in(19) => 
                           positive_inputs_4_19_port, shift_in(18) => 
                           positive_inputs_4_18_port, shift_in(17) => 
                           positive_inputs_4_17_port, shift_in(16) => 
                           positive_inputs_4_16_port, shift_in(15) => 
                           positive_inputs_4_15_port, shift_in(14) => 
                           positive_inputs_4_14_port, shift_in(13) => 
                           positive_inputs_4_13_port, shift_in(12) => 
                           positive_inputs_4_12_port, shift_in(11) => 
                           positive_inputs_4_11_port, shift_in(10) => 
                           positive_inputs_4_10_port, shift_in(9) => 
                           positive_inputs_4_9_port, shift_in(8) => 
                           positive_inputs_4_8_port, shift_in(7) => 
                           positive_inputs_4_7_port, shift_in(6) => 
                           positive_inputs_4_6_port, shift_in(5) => 
                           positive_inputs_4_5_port, shift_in(4) => 
                           positive_inputs_4_4_port, shift_in(3) => 
                           positive_inputs_4_3_port, shift_in(2) => 
                           positive_inputs_4_2_port, shift_in(1) => 
                           positive_inputs_4_1_port, shift_in(0) => n8, 
                           shift_out(63) => positive_inputs_5_63_port, 
                           shift_out(62) => positive_inputs_5_62_port, 
                           shift_out(61) => positive_inputs_5_61_port, 
                           shift_out(60) => positive_inputs_5_60_port, 
                           shift_out(59) => positive_inputs_5_59_port, 
                           shift_out(58) => positive_inputs_5_58_port, 
                           shift_out(57) => positive_inputs_5_57_port, 
                           shift_out(56) => positive_inputs_5_56_port, 
                           shift_out(55) => positive_inputs_5_55_port, 
                           shift_out(54) => positive_inputs_5_54_port, 
                           shift_out(53) => positive_inputs_5_53_port, 
                           shift_out(52) => positive_inputs_5_52_port, 
                           shift_out(51) => positive_inputs_5_51_port, 
                           shift_out(50) => positive_inputs_5_50_port, 
                           shift_out(49) => positive_inputs_5_49_port, 
                           shift_out(48) => positive_inputs_5_48_port, 
                           shift_out(47) => positive_inputs_5_47_port, 
                           shift_out(46) => positive_inputs_5_46_port, 
                           shift_out(45) => positive_inputs_5_45_port, 
                           shift_out(44) => positive_inputs_5_44_port, 
                           shift_out(43) => positive_inputs_5_43_port, 
                           shift_out(42) => positive_inputs_5_42_port, 
                           shift_out(41) => positive_inputs_5_41_port, 
                           shift_out(40) => positive_inputs_5_40_port, 
                           shift_out(39) => positive_inputs_5_39_port, 
                           shift_out(38) => positive_inputs_5_38_port, 
                           shift_out(37) => positive_inputs_5_37_port, 
                           shift_out(36) => positive_inputs_5_36_port, 
                           shift_out(35) => positive_inputs_5_35_port, 
                           shift_out(34) => positive_inputs_5_34_port, 
                           shift_out(33) => positive_inputs_5_33_port, 
                           shift_out(32) => positive_inputs_5_32_port, 
                           shift_out(31) => positive_inputs_5_31_port, 
                           shift_out(30) => positive_inputs_5_30_port, 
                           shift_out(29) => positive_inputs_5_29_port, 
                           shift_out(28) => positive_inputs_5_28_port, 
                           shift_out(27) => positive_inputs_5_27_port, 
                           shift_out(26) => positive_inputs_5_26_port, 
                           shift_out(25) => positive_inputs_5_25_port, 
                           shift_out(24) => positive_inputs_5_24_port, 
                           shift_out(23) => positive_inputs_5_23_port, 
                           shift_out(22) => positive_inputs_5_22_port, 
                           shift_out(21) => positive_inputs_5_21_port, 
                           shift_out(20) => positive_inputs_5_20_port, 
                           shift_out(19) => positive_inputs_5_19_port, 
                           shift_out(18) => positive_inputs_5_18_port, 
                           shift_out(17) => positive_inputs_5_17_port, 
                           shift_out(16) => positive_inputs_5_16_port, 
                           shift_out(15) => positive_inputs_5_15_port, 
                           shift_out(14) => positive_inputs_5_14_port, 
                           shift_out(13) => positive_inputs_5_13_port, 
                           shift_out(12) => positive_inputs_5_12_port, 
                           shift_out(11) => positive_inputs_5_11_port, 
                           shift_out(10) => positive_inputs_5_10_port, 
                           shift_out(9) => positive_inputs_5_9_port, 
                           shift_out(8) => positive_inputs_5_8_port, 
                           shift_out(7) => positive_inputs_5_7_port, 
                           shift_out(6) => positive_inputs_5_6_port, 
                           shift_out(5) => positive_inputs_5_5_port, 
                           shift_out(4) => positive_inputs_5_4_port, 
                           shift_out(3) => positive_inputs_5_3_port, 
                           shift_out(2) => positive_inputs_5_2_port, 
                           shift_out(1) => positive_inputs_5_1_port, 
                           shift_out(0) => n_1005);
   shifted_pos_6 : leftshifter_NbitShifter64_121 port map( shift_in(63) => 
                           positive_inputs_5_63_port, shift_in(62) => 
                           positive_inputs_5_62_port, shift_in(61) => 
                           positive_inputs_5_61_port, shift_in(60) => 
                           positive_inputs_5_60_port, shift_in(59) => 
                           positive_inputs_5_59_port, shift_in(58) => 
                           positive_inputs_5_58_port, shift_in(57) => 
                           positive_inputs_5_57_port, shift_in(56) => 
                           positive_inputs_5_56_port, shift_in(55) => 
                           positive_inputs_5_55_port, shift_in(54) => 
                           positive_inputs_5_54_port, shift_in(53) => 
                           positive_inputs_5_53_port, shift_in(52) => 
                           positive_inputs_5_52_port, shift_in(51) => 
                           positive_inputs_5_51_port, shift_in(50) => 
                           positive_inputs_5_50_port, shift_in(49) => 
                           positive_inputs_5_49_port, shift_in(48) => 
                           positive_inputs_5_48_port, shift_in(47) => n36, 
                           shift_in(46) => positive_inputs_5_46_port, 
                           shift_in(45) => positive_inputs_5_45_port, 
                           shift_in(44) => positive_inputs_5_44_port, 
                           shift_in(43) => positive_inputs_5_43_port, 
                           shift_in(42) => positive_inputs_5_42_port, 
                           shift_in(41) => positive_inputs_5_41_port, 
                           shift_in(40) => positive_inputs_5_40_port, 
                           shift_in(39) => positive_inputs_5_39_port, 
                           shift_in(38) => positive_inputs_5_38_port, 
                           shift_in(37) => n20, shift_in(36) => n19, 
                           shift_in(35) => n180, shift_in(34) => n178, 
                           shift_in(33) => n176, shift_in(32) => n174, 
                           shift_in(31) => n172, shift_in(30) => n170, 
                           shift_in(29) => n168, shift_in(28) => n166, 
                           shift_in(27) => n164, shift_in(26) => n162, 
                           shift_in(25) => n160, shift_in(24) => n158, 
                           shift_in(23) => n156, shift_in(22) => n154, 
                           shift_in(21) => n152, shift_in(20) => n150, 
                           shift_in(19) => n148, shift_in(18) => n146, 
                           shift_in(17) => n144, shift_in(16) => n142, 
                           shift_in(15) => n140, shift_in(14) => n138, 
                           shift_in(13) => n136, shift_in(12) => n134, 
                           shift_in(11) => n132, shift_in(10) => n130, 
                           shift_in(9) => n128, shift_in(8) => n126, 
                           shift_in(7) => n124, shift_in(6) => n122, 
                           shift_in(5) => n120, shift_in(4) => 
                           positive_inputs_5_4_port, shift_in(3) => 
                           positive_inputs_5_3_port, shift_in(2) => 
                           positive_inputs_5_2_port, shift_in(1) => 
                           positive_inputs_5_1_port, shift_in(0) => n8, 
                           shift_out(63) => positive_inputs_6_63_port, 
                           shift_out(62) => positive_inputs_6_62_port, 
                           shift_out(61) => positive_inputs_6_61_port, 
                           shift_out(60) => positive_inputs_6_60_port, 
                           shift_out(59) => positive_inputs_6_59_port, 
                           shift_out(58) => positive_inputs_6_58_port, 
                           shift_out(57) => positive_inputs_6_57_port, 
                           shift_out(56) => positive_inputs_6_56_port, 
                           shift_out(55) => positive_inputs_6_55_port, 
                           shift_out(54) => positive_inputs_6_54_port, 
                           shift_out(53) => positive_inputs_6_53_port, 
                           shift_out(52) => positive_inputs_6_52_port, 
                           shift_out(51) => positive_inputs_6_51_port, 
                           shift_out(50) => positive_inputs_6_50_port, 
                           shift_out(49) => positive_inputs_6_49_port, 
                           shift_out(48) => positive_inputs_6_48_port, 
                           shift_out(47) => positive_inputs_6_47_port, 
                           shift_out(46) => positive_inputs_6_46_port, 
                           shift_out(45) => positive_inputs_6_45_port, 
                           shift_out(44) => positive_inputs_6_44_port, 
                           shift_out(43) => positive_inputs_6_43_port, 
                           shift_out(42) => positive_inputs_6_42_port, 
                           shift_out(41) => positive_inputs_6_41_port, 
                           shift_out(40) => positive_inputs_6_40_port, 
                           shift_out(39) => positive_inputs_6_39_port, 
                           shift_out(38) => positive_inputs_6_38_port, 
                           shift_out(37) => positive_inputs_6_37_port, 
                           shift_out(36) => positive_inputs_6_36_port, 
                           shift_out(35) => positive_inputs_6_35_port, 
                           shift_out(34) => positive_inputs_6_34_port, 
                           shift_out(33) => positive_inputs_6_33_port, 
                           shift_out(32) => positive_inputs_6_32_port, 
                           shift_out(31) => positive_inputs_6_31_port, 
                           shift_out(30) => positive_inputs_6_30_port, 
                           shift_out(29) => positive_inputs_6_29_port, 
                           shift_out(28) => positive_inputs_6_28_port, 
                           shift_out(27) => positive_inputs_6_27_port, 
                           shift_out(26) => positive_inputs_6_26_port, 
                           shift_out(25) => positive_inputs_6_25_port, 
                           shift_out(24) => positive_inputs_6_24_port, 
                           shift_out(23) => positive_inputs_6_23_port, 
                           shift_out(22) => positive_inputs_6_22_port, 
                           shift_out(21) => positive_inputs_6_21_port, 
                           shift_out(20) => positive_inputs_6_20_port, 
                           shift_out(19) => positive_inputs_6_19_port, 
                           shift_out(18) => positive_inputs_6_18_port, 
                           shift_out(17) => positive_inputs_6_17_port, 
                           shift_out(16) => positive_inputs_6_16_port, 
                           shift_out(15) => positive_inputs_6_15_port, 
                           shift_out(14) => positive_inputs_6_14_port, 
                           shift_out(13) => positive_inputs_6_13_port, 
                           shift_out(12) => positive_inputs_6_12_port, 
                           shift_out(11) => positive_inputs_6_11_port, 
                           shift_out(10) => positive_inputs_6_10_port, 
                           shift_out(9) => positive_inputs_6_9_port, 
                           shift_out(8) => positive_inputs_6_8_port, 
                           shift_out(7) => positive_inputs_6_7_port, 
                           shift_out(6) => positive_inputs_6_6_port, 
                           shift_out(5) => positive_inputs_6_5_port, 
                           shift_out(4) => positive_inputs_6_4_port, 
                           shift_out(3) => positive_inputs_6_3_port, 
                           shift_out(2) => positive_inputs_6_2_port, 
                           shift_out(1) => positive_inputs_6_1_port, 
                           shift_out(0) => n_1006);
   shifted_pos_7 : leftshifter_NbitShifter64_120 port map( shift_in(63) => 
                           positive_inputs_6_63_port, shift_in(62) => 
                           positive_inputs_6_62_port, shift_in(61) => 
                           positive_inputs_6_61_port, shift_in(60) => 
                           positive_inputs_6_60_port, shift_in(59) => 
                           positive_inputs_6_59_port, shift_in(58) => 
                           positive_inputs_6_58_port, shift_in(57) => 
                           positive_inputs_6_57_port, shift_in(56) => 
                           positive_inputs_6_56_port, shift_in(55) => 
                           positive_inputs_6_55_port, shift_in(54) => 
                           positive_inputs_6_54_port, shift_in(53) => 
                           positive_inputs_6_53_port, shift_in(52) => 
                           positive_inputs_6_52_port, shift_in(51) => 
                           positive_inputs_6_51_port, shift_in(50) => 
                           positive_inputs_6_50_port, shift_in(49) => 
                           positive_inputs_6_49_port, shift_in(48) => 
                           positive_inputs_6_48_port, shift_in(47) => n35, 
                           shift_in(46) => positive_inputs_6_46_port, 
                           shift_in(45) => positive_inputs_6_45_port, 
                           shift_in(44) => positive_inputs_6_44_port, 
                           shift_in(43) => positive_inputs_6_43_port, 
                           shift_in(42) => positive_inputs_6_42_port, 
                           shift_in(41) => positive_inputs_6_41_port, 
                           shift_in(40) => positive_inputs_6_40_port, 
                           shift_in(39) => positive_inputs_6_39_port, 
                           shift_in(38) => positive_inputs_6_38_port, 
                           shift_in(37) => positive_inputs_6_37_port, 
                           shift_in(36) => positive_inputs_6_36_port, 
                           shift_in(35) => positive_inputs_6_35_port, 
                           shift_in(34) => positive_inputs_6_34_port, 
                           shift_in(33) => positive_inputs_6_33_port, 
                           shift_in(32) => positive_inputs_6_32_port, 
                           shift_in(31) => positive_inputs_6_31_port, 
                           shift_in(30) => positive_inputs_6_30_port, 
                           shift_in(29) => positive_inputs_6_29_port, 
                           shift_in(28) => positive_inputs_6_28_port, 
                           shift_in(27) => positive_inputs_6_27_port, 
                           shift_in(26) => positive_inputs_6_26_port, 
                           shift_in(25) => positive_inputs_6_25_port, 
                           shift_in(24) => positive_inputs_6_24_port, 
                           shift_in(23) => positive_inputs_6_23_port, 
                           shift_in(22) => positive_inputs_6_22_port, 
                           shift_in(21) => positive_inputs_6_21_port, 
                           shift_in(20) => positive_inputs_6_20_port, 
                           shift_in(19) => positive_inputs_6_19_port, 
                           shift_in(18) => positive_inputs_6_18_port, 
                           shift_in(17) => positive_inputs_6_17_port, 
                           shift_in(16) => positive_inputs_6_16_port, 
                           shift_in(15) => positive_inputs_6_15_port, 
                           shift_in(14) => positive_inputs_6_14_port, 
                           shift_in(13) => positive_inputs_6_13_port, 
                           shift_in(12) => positive_inputs_6_12_port, 
                           shift_in(11) => positive_inputs_6_11_port, 
                           shift_in(10) => positive_inputs_6_10_port, 
                           shift_in(9) => positive_inputs_6_9_port, shift_in(8)
                           => positive_inputs_6_8_port, shift_in(7) => 
                           positive_inputs_6_7_port, shift_in(6) => 
                           positive_inputs_6_6_port, shift_in(5) => 
                           positive_inputs_6_5_port, shift_in(4) => 
                           positive_inputs_6_4_port, shift_in(3) => 
                           positive_inputs_6_3_port, shift_in(2) => 
                           positive_inputs_6_2_port, shift_in(1) => 
                           positive_inputs_6_1_port, shift_in(0) => n8, 
                           shift_out(63) => positive_inputs_7_63_port, 
                           shift_out(62) => positive_inputs_7_62_port, 
                           shift_out(61) => positive_inputs_7_61_port, 
                           shift_out(60) => positive_inputs_7_60_port, 
                           shift_out(59) => positive_inputs_7_59_port, 
                           shift_out(58) => positive_inputs_7_58_port, 
                           shift_out(57) => positive_inputs_7_57_port, 
                           shift_out(56) => positive_inputs_7_56_port, 
                           shift_out(55) => positive_inputs_7_55_port, 
                           shift_out(54) => positive_inputs_7_54_port, 
                           shift_out(53) => positive_inputs_7_53_port, 
                           shift_out(52) => positive_inputs_7_52_port, 
                           shift_out(51) => positive_inputs_7_51_port, 
                           shift_out(50) => positive_inputs_7_50_port, 
                           shift_out(49) => positive_inputs_7_49_port, 
                           shift_out(48) => positive_inputs_7_48_port, 
                           shift_out(47) => positive_inputs_7_47_port, 
                           shift_out(46) => positive_inputs_7_46_port, 
                           shift_out(45) => positive_inputs_7_45_port, 
                           shift_out(44) => positive_inputs_7_44_port, 
                           shift_out(43) => positive_inputs_7_43_port, 
                           shift_out(42) => positive_inputs_7_42_port, 
                           shift_out(41) => positive_inputs_7_41_port, 
                           shift_out(40) => positive_inputs_7_40_port, 
                           shift_out(39) => positive_inputs_7_39_port, 
                           shift_out(38) => positive_inputs_7_38_port, 
                           shift_out(37) => positive_inputs_7_37_port, 
                           shift_out(36) => positive_inputs_7_36_port, 
                           shift_out(35) => positive_inputs_7_35_port, 
                           shift_out(34) => positive_inputs_7_34_port, 
                           shift_out(33) => positive_inputs_7_33_port, 
                           shift_out(32) => positive_inputs_7_32_port, 
                           shift_out(31) => positive_inputs_7_31_port, 
                           shift_out(30) => positive_inputs_7_30_port, 
                           shift_out(29) => positive_inputs_7_29_port, 
                           shift_out(28) => positive_inputs_7_28_port, 
                           shift_out(27) => positive_inputs_7_27_port, 
                           shift_out(26) => positive_inputs_7_26_port, 
                           shift_out(25) => positive_inputs_7_25_port, 
                           shift_out(24) => positive_inputs_7_24_port, 
                           shift_out(23) => positive_inputs_7_23_port, 
                           shift_out(22) => positive_inputs_7_22_port, 
                           shift_out(21) => positive_inputs_7_21_port, 
                           shift_out(20) => positive_inputs_7_20_port, 
                           shift_out(19) => positive_inputs_7_19_port, 
                           shift_out(18) => positive_inputs_7_18_port, 
                           shift_out(17) => positive_inputs_7_17_port, 
                           shift_out(16) => positive_inputs_7_16_port, 
                           shift_out(15) => positive_inputs_7_15_port, 
                           shift_out(14) => positive_inputs_7_14_port, 
                           shift_out(13) => positive_inputs_7_13_port, 
                           shift_out(12) => positive_inputs_7_12_port, 
                           shift_out(11) => positive_inputs_7_11_port, 
                           shift_out(10) => positive_inputs_7_10_port, 
                           shift_out(9) => positive_inputs_7_9_port, 
                           shift_out(8) => positive_inputs_7_8_port, 
                           shift_out(7) => positive_inputs_7_7_port, 
                           shift_out(6) => positive_inputs_7_6_port, 
                           shift_out(5) => positive_inputs_7_5_port, 
                           shift_out(4) => positive_inputs_7_4_port, 
                           shift_out(3) => positive_inputs_7_3_port, 
                           shift_out(2) => positive_inputs_7_2_port, 
                           shift_out(1) => positive_inputs_7_1_port, 
                           shift_out(0) => n_1007);
   shifted_pos_8 : leftshifter_NbitShifter64_119 port map( shift_in(63) => 
                           positive_inputs_7_63_port, shift_in(62) => 
                           positive_inputs_7_62_port, shift_in(61) => 
                           positive_inputs_7_61_port, shift_in(60) => 
                           positive_inputs_7_60_port, shift_in(59) => 
                           positive_inputs_7_59_port, shift_in(58) => 
                           positive_inputs_7_58_port, shift_in(57) => 
                           positive_inputs_7_57_port, shift_in(56) => 
                           positive_inputs_7_56_port, shift_in(55) => 
                           positive_inputs_7_55_port, shift_in(54) => 
                           positive_inputs_7_54_port, shift_in(53) => 
                           positive_inputs_7_53_port, shift_in(52) => 
                           positive_inputs_7_52_port, shift_in(51) => 
                           positive_inputs_7_51_port, shift_in(50) => 
                           positive_inputs_7_50_port, shift_in(49) => 
                           positive_inputs_7_49_port, shift_in(48) => 
                           positive_inputs_7_48_port, shift_in(47) => n34, 
                           shift_in(46) => positive_inputs_7_46_port, 
                           shift_in(45) => positive_inputs_7_45_port, 
                           shift_in(44) => positive_inputs_7_44_port, 
                           shift_in(43) => positive_inputs_7_43_port, 
                           shift_in(42) => positive_inputs_7_42_port, 
                           shift_in(41) => positive_inputs_7_41_port, 
                           shift_in(40) => positive_inputs_7_40_port, 
                           shift_in(39) => positive_inputs_7_39_port, 
                           shift_in(38) => positive_inputs_7_38_port, 
                           shift_in(37) => positive_inputs_7_37_port, 
                           shift_in(36) => positive_inputs_7_36_port, 
                           shift_in(35) => positive_inputs_7_35_port, 
                           shift_in(34) => positive_inputs_7_34_port, 
                           shift_in(33) => positive_inputs_7_33_port, 
                           shift_in(32) => positive_inputs_7_32_port, 
                           shift_in(31) => positive_inputs_7_31_port, 
                           shift_in(30) => positive_inputs_7_30_port, 
                           shift_in(29) => positive_inputs_7_29_port, 
                           shift_in(28) => positive_inputs_7_28_port, 
                           shift_in(27) => positive_inputs_7_27_port, 
                           shift_in(26) => positive_inputs_7_26_port, 
                           shift_in(25) => positive_inputs_7_25_port, 
                           shift_in(24) => positive_inputs_7_24_port, 
                           shift_in(23) => positive_inputs_7_23_port, 
                           shift_in(22) => positive_inputs_7_22_port, 
                           shift_in(21) => positive_inputs_7_21_port, 
                           shift_in(20) => positive_inputs_7_20_port, 
                           shift_in(19) => positive_inputs_7_19_port, 
                           shift_in(18) => positive_inputs_7_18_port, 
                           shift_in(17) => positive_inputs_7_17_port, 
                           shift_in(16) => positive_inputs_7_16_port, 
                           shift_in(15) => positive_inputs_7_15_port, 
                           shift_in(14) => positive_inputs_7_14_port, 
                           shift_in(13) => positive_inputs_7_13_port, 
                           shift_in(12) => positive_inputs_7_12_port, 
                           shift_in(11) => positive_inputs_7_11_port, 
                           shift_in(10) => positive_inputs_7_10_port, 
                           shift_in(9) => positive_inputs_7_9_port, shift_in(8)
                           => positive_inputs_7_8_port, shift_in(7) => 
                           positive_inputs_7_7_port, shift_in(6) => 
                           positive_inputs_7_6_port, shift_in(5) => 
                           positive_inputs_7_5_port, shift_in(4) => 
                           positive_inputs_7_4_port, shift_in(3) => 
                           positive_inputs_7_3_port, shift_in(2) => 
                           positive_inputs_7_2_port, shift_in(1) => 
                           positive_inputs_7_1_port, shift_in(0) => n8, 
                           shift_out(63) => positive_inputs_8_63_port, 
                           shift_out(62) => positive_inputs_8_62_port, 
                           shift_out(61) => positive_inputs_8_61_port, 
                           shift_out(60) => positive_inputs_8_60_port, 
                           shift_out(59) => positive_inputs_8_59_port, 
                           shift_out(58) => positive_inputs_8_58_port, 
                           shift_out(57) => positive_inputs_8_57_port, 
                           shift_out(56) => positive_inputs_8_56_port, 
                           shift_out(55) => positive_inputs_8_55_port, 
                           shift_out(54) => positive_inputs_8_54_port, 
                           shift_out(53) => positive_inputs_8_53_port, 
                           shift_out(52) => positive_inputs_8_52_port, 
                           shift_out(51) => positive_inputs_8_51_port, 
                           shift_out(50) => positive_inputs_8_50_port, 
                           shift_out(49) => positive_inputs_8_49_port, 
                           shift_out(48) => positive_inputs_8_48_port, 
                           shift_out(47) => positive_inputs_8_47_port, 
                           shift_out(46) => positive_inputs_8_46_port, 
                           shift_out(45) => positive_inputs_8_45_port, 
                           shift_out(44) => positive_inputs_8_44_port, 
                           shift_out(43) => positive_inputs_8_43_port, 
                           shift_out(42) => positive_inputs_8_42_port, 
                           shift_out(41) => positive_inputs_8_41_port, 
                           shift_out(40) => positive_inputs_8_40_port, 
                           shift_out(39) => positive_inputs_8_39_port, 
                           shift_out(38) => positive_inputs_8_38_port, 
                           shift_out(37) => positive_inputs_8_37_port, 
                           shift_out(36) => positive_inputs_8_36_port, 
                           shift_out(35) => positive_inputs_8_35_port, 
                           shift_out(34) => positive_inputs_8_34_port, 
                           shift_out(33) => positive_inputs_8_33_port, 
                           shift_out(32) => positive_inputs_8_32_port, 
                           shift_out(31) => positive_inputs_8_31_port, 
                           shift_out(30) => positive_inputs_8_30_port, 
                           shift_out(29) => positive_inputs_8_29_port, 
                           shift_out(28) => positive_inputs_8_28_port, 
                           shift_out(27) => positive_inputs_8_27_port, 
                           shift_out(26) => positive_inputs_8_26_port, 
                           shift_out(25) => positive_inputs_8_25_port, 
                           shift_out(24) => positive_inputs_8_24_port, 
                           shift_out(23) => positive_inputs_8_23_port, 
                           shift_out(22) => positive_inputs_8_22_port, 
                           shift_out(21) => positive_inputs_8_21_port, 
                           shift_out(20) => positive_inputs_8_20_port, 
                           shift_out(19) => positive_inputs_8_19_port, 
                           shift_out(18) => positive_inputs_8_18_port, 
                           shift_out(17) => positive_inputs_8_17_port, 
                           shift_out(16) => positive_inputs_8_16_port, 
                           shift_out(15) => positive_inputs_8_15_port, 
                           shift_out(14) => positive_inputs_8_14_port, 
                           shift_out(13) => positive_inputs_8_13_port, 
                           shift_out(12) => positive_inputs_8_12_port, 
                           shift_out(11) => positive_inputs_8_11_port, 
                           shift_out(10) => positive_inputs_8_10_port, 
                           shift_out(9) => positive_inputs_8_9_port, 
                           shift_out(8) => positive_inputs_8_8_port, 
                           shift_out(7) => positive_inputs_8_7_port, 
                           shift_out(6) => positive_inputs_8_6_port, 
                           shift_out(5) => positive_inputs_8_5_port, 
                           shift_out(4) => positive_inputs_8_4_port, 
                           shift_out(3) => positive_inputs_8_3_port, 
                           shift_out(2) => positive_inputs_8_2_port, 
                           shift_out(1) => positive_inputs_8_1_port, 
                           shift_out(0) => n_1008);
   shifted_pos_9 : leftshifter_NbitShifter64_118 port map( shift_in(63) => 
                           positive_inputs_8_63_port, shift_in(62) => 
                           positive_inputs_8_62_port, shift_in(61) => 
                           positive_inputs_8_61_port, shift_in(60) => 
                           positive_inputs_8_60_port, shift_in(59) => 
                           positive_inputs_8_59_port, shift_in(58) => 
                           positive_inputs_8_58_port, shift_in(57) => 
                           positive_inputs_8_57_port, shift_in(56) => 
                           positive_inputs_8_56_port, shift_in(55) => 
                           positive_inputs_8_55_port, shift_in(54) => 
                           positive_inputs_8_54_port, shift_in(53) => 
                           positive_inputs_8_53_port, shift_in(52) => 
                           positive_inputs_8_52_port, shift_in(51) => 
                           positive_inputs_8_51_port, shift_in(50) => 
                           positive_inputs_8_50_port, shift_in(49) => 
                           positive_inputs_8_49_port, shift_in(48) => 
                           positive_inputs_8_48_port, shift_in(47) => n33, 
                           shift_in(46) => positive_inputs_8_46_port, 
                           shift_in(45) => positive_inputs_8_45_port, 
                           shift_in(44) => positive_inputs_8_44_port, 
                           shift_in(43) => positive_inputs_8_43_port, 
                           shift_in(42) => positive_inputs_8_42_port, 
                           shift_in(41) => positive_inputs_8_41_port, 
                           shift_in(40) => positive_inputs_8_40_port, 
                           shift_in(39) => positive_inputs_8_39_port, 
                           shift_in(38) => positive_inputs_8_38_port, 
                           shift_in(37) => positive_inputs_8_37_port, 
                           shift_in(36) => positive_inputs_8_36_port, 
                           shift_in(35) => positive_inputs_8_35_port, 
                           shift_in(34) => positive_inputs_8_34_port, 
                           shift_in(33) => positive_inputs_8_33_port, 
                           shift_in(32) => positive_inputs_8_32_port, 
                           shift_in(31) => positive_inputs_8_31_port, 
                           shift_in(30) => positive_inputs_8_30_port, 
                           shift_in(29) => positive_inputs_8_29_port, 
                           shift_in(28) => positive_inputs_8_28_port, 
                           shift_in(27) => positive_inputs_8_27_port, 
                           shift_in(26) => positive_inputs_8_26_port, 
                           shift_in(25) => positive_inputs_8_25_port, 
                           shift_in(24) => positive_inputs_8_24_port, 
                           shift_in(23) => positive_inputs_8_23_port, 
                           shift_in(22) => positive_inputs_8_22_port, 
                           shift_in(21) => positive_inputs_8_21_port, 
                           shift_in(20) => positive_inputs_8_20_port, 
                           shift_in(19) => positive_inputs_8_19_port, 
                           shift_in(18) => positive_inputs_8_18_port, 
                           shift_in(17) => positive_inputs_8_17_port, 
                           shift_in(16) => positive_inputs_8_16_port, 
                           shift_in(15) => positive_inputs_8_15_port, 
                           shift_in(14) => positive_inputs_8_14_port, 
                           shift_in(13) => positive_inputs_8_13_port, 
                           shift_in(12) => positive_inputs_8_12_port, 
                           shift_in(11) => positive_inputs_8_11_port, 
                           shift_in(10) => positive_inputs_8_10_port, 
                           shift_in(9) => positive_inputs_8_9_port, shift_in(8)
                           => positive_inputs_8_8_port, shift_in(7) => 
                           positive_inputs_8_7_port, shift_in(6) => 
                           positive_inputs_8_6_port, shift_in(5) => 
                           positive_inputs_8_5_port, shift_in(4) => 
                           positive_inputs_8_4_port, shift_in(3) => 
                           positive_inputs_8_3_port, shift_in(2) => 
                           positive_inputs_8_2_port, shift_in(1) => 
                           positive_inputs_8_1_port, shift_in(0) => n8, 
                           shift_out(63) => positive_inputs_9_63_port, 
                           shift_out(62) => positive_inputs_9_62_port, 
                           shift_out(61) => positive_inputs_9_61_port, 
                           shift_out(60) => positive_inputs_9_60_port, 
                           shift_out(59) => positive_inputs_9_59_port, 
                           shift_out(58) => positive_inputs_9_58_port, 
                           shift_out(57) => positive_inputs_9_57_port, 
                           shift_out(56) => positive_inputs_9_56_port, 
                           shift_out(55) => positive_inputs_9_55_port, 
                           shift_out(54) => positive_inputs_9_54_port, 
                           shift_out(53) => positive_inputs_9_53_port, 
                           shift_out(52) => positive_inputs_9_52_port, 
                           shift_out(51) => positive_inputs_9_51_port, 
                           shift_out(50) => positive_inputs_9_50_port, 
                           shift_out(49) => positive_inputs_9_49_port, 
                           shift_out(48) => positive_inputs_9_48_port, 
                           shift_out(47) => positive_inputs_9_47_port, 
                           shift_out(46) => positive_inputs_9_46_port, 
                           shift_out(45) => positive_inputs_9_45_port, 
                           shift_out(44) => positive_inputs_9_44_port, 
                           shift_out(43) => positive_inputs_9_43_port, 
                           shift_out(42) => positive_inputs_9_42_port, 
                           shift_out(41) => positive_inputs_9_41_port, 
                           shift_out(40) => positive_inputs_9_40_port, 
                           shift_out(39) => positive_inputs_9_39_port, 
                           shift_out(38) => positive_inputs_9_38_port, 
                           shift_out(37) => positive_inputs_9_37_port, 
                           shift_out(36) => positive_inputs_9_36_port, 
                           shift_out(35) => positive_inputs_9_35_port, 
                           shift_out(34) => positive_inputs_9_34_port, 
                           shift_out(33) => positive_inputs_9_33_port, 
                           shift_out(32) => positive_inputs_9_32_port, 
                           shift_out(31) => positive_inputs_9_31_port, 
                           shift_out(30) => positive_inputs_9_30_port, 
                           shift_out(29) => positive_inputs_9_29_port, 
                           shift_out(28) => positive_inputs_9_28_port, 
                           shift_out(27) => positive_inputs_9_27_port, 
                           shift_out(26) => positive_inputs_9_26_port, 
                           shift_out(25) => positive_inputs_9_25_port, 
                           shift_out(24) => positive_inputs_9_24_port, 
                           shift_out(23) => positive_inputs_9_23_port, 
                           shift_out(22) => positive_inputs_9_22_port, 
                           shift_out(21) => positive_inputs_9_21_port, 
                           shift_out(20) => positive_inputs_9_20_port, 
                           shift_out(19) => positive_inputs_9_19_port, 
                           shift_out(18) => positive_inputs_9_18_port, 
                           shift_out(17) => positive_inputs_9_17_port, 
                           shift_out(16) => positive_inputs_9_16_port, 
                           shift_out(15) => positive_inputs_9_15_port, 
                           shift_out(14) => positive_inputs_9_14_port, 
                           shift_out(13) => positive_inputs_9_13_port, 
                           shift_out(12) => positive_inputs_9_12_port, 
                           shift_out(11) => positive_inputs_9_11_port, 
                           shift_out(10) => positive_inputs_9_10_port, 
                           shift_out(9) => positive_inputs_9_9_port, 
                           shift_out(8) => positive_inputs_9_8_port, 
                           shift_out(7) => positive_inputs_9_7_port, 
                           shift_out(6) => positive_inputs_9_6_port, 
                           shift_out(5) => positive_inputs_9_5_port, 
                           shift_out(4) => positive_inputs_9_4_port, 
                           shift_out(3) => positive_inputs_9_3_port, 
                           shift_out(2) => positive_inputs_9_2_port, 
                           shift_out(1) => positive_inputs_9_1_port, 
                           shift_out(0) => n_1009);
   shifted_pos_10 : leftshifter_NbitShifter64_117 port map( shift_in(63) => 
                           positive_inputs_9_63_port, shift_in(62) => 
                           positive_inputs_9_62_port, shift_in(61) => 
                           positive_inputs_9_61_port, shift_in(60) => 
                           positive_inputs_9_60_port, shift_in(59) => 
                           positive_inputs_9_59_port, shift_in(58) => 
                           positive_inputs_9_58_port, shift_in(57) => 
                           positive_inputs_9_57_port, shift_in(56) => 
                           positive_inputs_9_56_port, shift_in(55) => 
                           positive_inputs_9_55_port, shift_in(54) => 
                           positive_inputs_9_54_port, shift_in(53) => 
                           positive_inputs_9_53_port, shift_in(52) => 
                           positive_inputs_9_52_port, shift_in(51) => 
                           positive_inputs_9_51_port, shift_in(50) => 
                           positive_inputs_9_50_port, shift_in(49) => 
                           positive_inputs_9_49_port, shift_in(48) => 
                           positive_inputs_9_48_port, shift_in(47) => n32, 
                           shift_in(46) => positive_inputs_9_46_port, 
                           shift_in(45) => positive_inputs_9_45_port, 
                           shift_in(44) => positive_inputs_9_44_port, 
                           shift_in(43) => positive_inputs_9_43_port, 
                           shift_in(42) => positive_inputs_9_42_port, 
                           shift_in(41) => positive_inputs_9_41_port, 
                           shift_in(40) => positive_inputs_9_40_port, 
                           shift_in(39) => positive_inputs_9_39_port, 
                           shift_in(38) => positive_inputs_9_38_port, 
                           shift_in(37) => positive_inputs_9_37_port, 
                           shift_in(36) => positive_inputs_9_36_port, 
                           shift_in(35) => positive_inputs_9_35_port, 
                           shift_in(34) => positive_inputs_9_34_port, 
                           shift_in(33) => positive_inputs_9_33_port, 
                           shift_in(32) => positive_inputs_9_32_port, 
                           shift_in(31) => positive_inputs_9_31_port, 
                           shift_in(30) => positive_inputs_9_30_port, 
                           shift_in(29) => positive_inputs_9_29_port, 
                           shift_in(28) => positive_inputs_9_28_port, 
                           shift_in(27) => positive_inputs_9_27_port, 
                           shift_in(26) => positive_inputs_9_26_port, 
                           shift_in(25) => positive_inputs_9_25_port, 
                           shift_in(24) => positive_inputs_9_24_port, 
                           shift_in(23) => positive_inputs_9_23_port, 
                           shift_in(22) => positive_inputs_9_22_port, 
                           shift_in(21) => positive_inputs_9_21_port, 
                           shift_in(20) => positive_inputs_9_20_port, 
                           shift_in(19) => positive_inputs_9_19_port, 
                           shift_in(18) => positive_inputs_9_18_port, 
                           shift_in(17) => positive_inputs_9_17_port, 
                           shift_in(16) => positive_inputs_9_16_port, 
                           shift_in(15) => positive_inputs_9_15_port, 
                           shift_in(14) => positive_inputs_9_14_port, 
                           shift_in(13) => positive_inputs_9_13_port, 
                           shift_in(12) => positive_inputs_9_12_port, 
                           shift_in(11) => positive_inputs_9_11_port, 
                           shift_in(10) => positive_inputs_9_10_port, 
                           shift_in(9) => positive_inputs_9_9_port, shift_in(8)
                           => positive_inputs_9_8_port, shift_in(7) => 
                           positive_inputs_9_7_port, shift_in(6) => 
                           positive_inputs_9_6_port, shift_in(5) => 
                           positive_inputs_9_5_port, shift_in(4) => 
                           positive_inputs_9_4_port, shift_in(3) => 
                           positive_inputs_9_3_port, shift_in(2) => 
                           positive_inputs_9_2_port, shift_in(1) => 
                           positive_inputs_9_1_port, shift_in(0) => n8, 
                           shift_out(63) => positive_inputs_10_63_port, 
                           shift_out(62) => positive_inputs_10_62_port, 
                           shift_out(61) => positive_inputs_10_61_port, 
                           shift_out(60) => positive_inputs_10_60_port, 
                           shift_out(59) => positive_inputs_10_59_port, 
                           shift_out(58) => positive_inputs_10_58_port, 
                           shift_out(57) => positive_inputs_10_57_port, 
                           shift_out(56) => positive_inputs_10_56_port, 
                           shift_out(55) => positive_inputs_10_55_port, 
                           shift_out(54) => positive_inputs_10_54_port, 
                           shift_out(53) => positive_inputs_10_53_port, 
                           shift_out(52) => positive_inputs_10_52_port, 
                           shift_out(51) => positive_inputs_10_51_port, 
                           shift_out(50) => positive_inputs_10_50_port, 
                           shift_out(49) => positive_inputs_10_49_port, 
                           shift_out(48) => positive_inputs_10_48_port, 
                           shift_out(47) => positive_inputs_10_47_port, 
                           shift_out(46) => positive_inputs_10_46_port, 
                           shift_out(45) => positive_inputs_10_45_port, 
                           shift_out(44) => positive_inputs_10_44_port, 
                           shift_out(43) => positive_inputs_10_43_port, 
                           shift_out(42) => positive_inputs_10_42_port, 
                           shift_out(41) => positive_inputs_10_41_port, 
                           shift_out(40) => positive_inputs_10_40_port, 
                           shift_out(39) => positive_inputs_10_39_port, 
                           shift_out(38) => positive_inputs_10_38_port, 
                           shift_out(37) => positive_inputs_10_37_port, 
                           shift_out(36) => positive_inputs_10_36_port, 
                           shift_out(35) => positive_inputs_10_35_port, 
                           shift_out(34) => positive_inputs_10_34_port, 
                           shift_out(33) => positive_inputs_10_33_port, 
                           shift_out(32) => positive_inputs_10_32_port, 
                           shift_out(31) => positive_inputs_10_31_port, 
                           shift_out(30) => positive_inputs_10_30_port, 
                           shift_out(29) => positive_inputs_10_29_port, 
                           shift_out(28) => positive_inputs_10_28_port, 
                           shift_out(27) => positive_inputs_10_27_port, 
                           shift_out(26) => positive_inputs_10_26_port, 
                           shift_out(25) => positive_inputs_10_25_port, 
                           shift_out(24) => positive_inputs_10_24_port, 
                           shift_out(23) => positive_inputs_10_23_port, 
                           shift_out(22) => positive_inputs_10_22_port, 
                           shift_out(21) => positive_inputs_10_21_port, 
                           shift_out(20) => positive_inputs_10_20_port, 
                           shift_out(19) => positive_inputs_10_19_port, 
                           shift_out(18) => positive_inputs_10_18_port, 
                           shift_out(17) => positive_inputs_10_17_port, 
                           shift_out(16) => positive_inputs_10_16_port, 
                           shift_out(15) => positive_inputs_10_15_port, 
                           shift_out(14) => positive_inputs_10_14_port, 
                           shift_out(13) => positive_inputs_10_13_port, 
                           shift_out(12) => positive_inputs_10_12_port, 
                           shift_out(11) => positive_inputs_10_11_port, 
                           shift_out(10) => positive_inputs_10_10_port, 
                           shift_out(9) => positive_inputs_10_9_port, 
                           shift_out(8) => positive_inputs_10_8_port, 
                           shift_out(7) => positive_inputs_10_7_port, 
                           shift_out(6) => positive_inputs_10_6_port, 
                           shift_out(5) => positive_inputs_10_5_port, 
                           shift_out(4) => positive_inputs_10_4_port, 
                           shift_out(3) => positive_inputs_10_3_port, 
                           shift_out(2) => positive_inputs_10_2_port, 
                           shift_out(1) => positive_inputs_10_1_port, 
                           shift_out(0) => n_1010);
   shifted_pos_11 : leftshifter_NbitShifter64_116 port map( shift_in(63) => 
                           positive_inputs_10_63_port, shift_in(62) => 
                           positive_inputs_10_62_port, shift_in(61) => 
                           positive_inputs_10_61_port, shift_in(60) => 
                           positive_inputs_10_60_port, shift_in(59) => 
                           positive_inputs_10_59_port, shift_in(58) => 
                           positive_inputs_10_58_port, shift_in(57) => 
                           positive_inputs_10_57_port, shift_in(56) => 
                           positive_inputs_10_56_port, shift_in(55) => 
                           positive_inputs_10_55_port, shift_in(54) => 
                           positive_inputs_10_54_port, shift_in(53) => 
                           positive_inputs_10_53_port, shift_in(52) => 
                           positive_inputs_10_52_port, shift_in(51) => 
                           positive_inputs_10_51_port, shift_in(50) => 
                           positive_inputs_10_50_port, shift_in(49) => 
                           positive_inputs_10_49_port, shift_in(48) => 
                           positive_inputs_10_48_port, shift_in(47) => n31, 
                           shift_in(46) => positive_inputs_10_46_port, 
                           shift_in(45) => positive_inputs_10_45_port, 
                           shift_in(44) => positive_inputs_10_44_port, 
                           shift_in(43) => positive_inputs_10_43_port, 
                           shift_in(42) => positive_inputs_10_42_port, 
                           shift_in(41) => positive_inputs_10_41_port, 
                           shift_in(40) => positive_inputs_10_40_port, 
                           shift_in(39) => positive_inputs_10_39_port, 
                           shift_in(38) => positive_inputs_10_38_port, 
                           shift_in(37) => positive_inputs_10_37_port, 
                           shift_in(36) => positive_inputs_10_36_port, 
                           shift_in(35) => positive_inputs_10_35_port, 
                           shift_in(34) => positive_inputs_10_34_port, 
                           shift_in(33) => positive_inputs_10_33_port, 
                           shift_in(32) => positive_inputs_10_32_port, 
                           shift_in(31) => positive_inputs_10_31_port, 
                           shift_in(30) => positive_inputs_10_30_port, 
                           shift_in(29) => positive_inputs_10_29_port, 
                           shift_in(28) => positive_inputs_10_28_port, 
                           shift_in(27) => positive_inputs_10_27_port, 
                           shift_in(26) => positive_inputs_10_26_port, 
                           shift_in(25) => positive_inputs_10_25_port, 
                           shift_in(24) => positive_inputs_10_24_port, 
                           shift_in(23) => positive_inputs_10_23_port, 
                           shift_in(22) => positive_inputs_10_22_port, 
                           shift_in(21) => positive_inputs_10_21_port, 
                           shift_in(20) => positive_inputs_10_20_port, 
                           shift_in(19) => positive_inputs_10_19_port, 
                           shift_in(18) => positive_inputs_10_18_port, 
                           shift_in(17) => positive_inputs_10_17_port, 
                           shift_in(16) => positive_inputs_10_16_port, 
                           shift_in(15) => positive_inputs_10_15_port, 
                           shift_in(14) => positive_inputs_10_14_port, 
                           shift_in(13) => positive_inputs_10_13_port, 
                           shift_in(12) => positive_inputs_10_12_port, 
                           shift_in(11) => positive_inputs_10_11_port, 
                           shift_in(10) => positive_inputs_10_10_port, 
                           shift_in(9) => positive_inputs_10_9_port, 
                           shift_in(8) => positive_inputs_10_8_port, 
                           shift_in(7) => positive_inputs_10_7_port, 
                           shift_in(6) => positive_inputs_10_6_port, 
                           shift_in(5) => positive_inputs_10_5_port, 
                           shift_in(4) => positive_inputs_10_4_port, 
                           shift_in(3) => positive_inputs_10_3_port, 
                           shift_in(2) => positive_inputs_10_2_port, 
                           shift_in(1) => positive_inputs_10_1_port, 
                           shift_in(0) => n8, shift_out(63) => 
                           positive_inputs_11_63_port, shift_out(62) => 
                           positive_inputs_11_62_port, shift_out(61) => 
                           positive_inputs_11_61_port, shift_out(60) => 
                           positive_inputs_11_60_port, shift_out(59) => 
                           positive_inputs_11_59_port, shift_out(58) => 
                           positive_inputs_11_58_port, shift_out(57) => 
                           positive_inputs_11_57_port, shift_out(56) => 
                           positive_inputs_11_56_port, shift_out(55) => 
                           positive_inputs_11_55_port, shift_out(54) => 
                           positive_inputs_11_54_port, shift_out(53) => 
                           positive_inputs_11_53_port, shift_out(52) => 
                           positive_inputs_11_52_port, shift_out(51) => 
                           positive_inputs_11_51_port, shift_out(50) => 
                           positive_inputs_11_50_port, shift_out(49) => 
                           positive_inputs_11_49_port, shift_out(48) => 
                           positive_inputs_11_48_port, shift_out(47) => 
                           positive_inputs_11_47_port, shift_out(46) => 
                           positive_inputs_11_46_port, shift_out(45) => 
                           positive_inputs_11_45_port, shift_out(44) => 
                           positive_inputs_11_44_port, shift_out(43) => 
                           positive_inputs_11_43_port, shift_out(42) => 
                           positive_inputs_11_42_port, shift_out(41) => 
                           positive_inputs_11_41_port, shift_out(40) => 
                           positive_inputs_11_40_port, shift_out(39) => 
                           positive_inputs_11_39_port, shift_out(38) => 
                           positive_inputs_11_38_port, shift_out(37) => 
                           positive_inputs_11_37_port, shift_out(36) => 
                           positive_inputs_11_36_port, shift_out(35) => 
                           positive_inputs_11_35_port, shift_out(34) => 
                           positive_inputs_11_34_port, shift_out(33) => 
                           positive_inputs_11_33_port, shift_out(32) => 
                           positive_inputs_11_32_port, shift_out(31) => 
                           positive_inputs_11_31_port, shift_out(30) => 
                           positive_inputs_11_30_port, shift_out(29) => 
                           positive_inputs_11_29_port, shift_out(28) => 
                           positive_inputs_11_28_port, shift_out(27) => 
                           positive_inputs_11_27_port, shift_out(26) => 
                           positive_inputs_11_26_port, shift_out(25) => 
                           positive_inputs_11_25_port, shift_out(24) => 
                           positive_inputs_11_24_port, shift_out(23) => 
                           positive_inputs_11_23_port, shift_out(22) => 
                           positive_inputs_11_22_port, shift_out(21) => 
                           positive_inputs_11_21_port, shift_out(20) => 
                           positive_inputs_11_20_port, shift_out(19) => 
                           positive_inputs_11_19_port, shift_out(18) => 
                           positive_inputs_11_18_port, shift_out(17) => 
                           positive_inputs_11_17_port, shift_out(16) => 
                           positive_inputs_11_16_port, shift_out(15) => 
                           positive_inputs_11_15_port, shift_out(14) => 
                           positive_inputs_11_14_port, shift_out(13) => 
                           positive_inputs_11_13_port, shift_out(12) => 
                           positive_inputs_11_12_port, shift_out(11) => 
                           positive_inputs_11_11_port, shift_out(10) => 
                           positive_inputs_11_10_port, shift_out(9) => 
                           positive_inputs_11_9_port, shift_out(8) => 
                           positive_inputs_11_8_port, shift_out(7) => 
                           positive_inputs_11_7_port, shift_out(6) => 
                           positive_inputs_11_6_port, shift_out(5) => 
                           positive_inputs_11_5_port, shift_out(4) => 
                           positive_inputs_11_4_port, shift_out(3) => 
                           positive_inputs_11_3_port, shift_out(2) => 
                           positive_inputs_11_2_port, shift_out(1) => 
                           positive_inputs_11_1_port, shift_out(0) => n_1011);
   shifted_pos_12 : leftshifter_NbitShifter64_115 port map( shift_in(63) => 
                           positive_inputs_11_63_port, shift_in(62) => 
                           positive_inputs_11_62_port, shift_in(61) => 
                           positive_inputs_11_61_port, shift_in(60) => 
                           positive_inputs_11_60_port, shift_in(59) => 
                           positive_inputs_11_59_port, shift_in(58) => 
                           positive_inputs_11_58_port, shift_in(57) => 
                           positive_inputs_11_57_port, shift_in(56) => 
                           positive_inputs_11_56_port, shift_in(55) => 
                           positive_inputs_11_55_port, shift_in(54) => 
                           positive_inputs_11_54_port, shift_in(53) => 
                           positive_inputs_11_53_port, shift_in(52) => 
                           positive_inputs_11_52_port, shift_in(51) => 
                           positive_inputs_11_51_port, shift_in(50) => 
                           positive_inputs_11_50_port, shift_in(49) => 
                           positive_inputs_11_49_port, shift_in(48) => 
                           positive_inputs_11_48_port, shift_in(47) => n30, 
                           shift_in(46) => positive_inputs_11_46_port, 
                           shift_in(45) => positive_inputs_11_45_port, 
                           shift_in(44) => positive_inputs_11_44_port, 
                           shift_in(43) => positive_inputs_11_43_port, 
                           shift_in(42) => positive_inputs_11_42_port, 
                           shift_in(41) => positive_inputs_11_41_port, 
                           shift_in(40) => positive_inputs_11_40_port, 
                           shift_in(39) => positive_inputs_11_39_port, 
                           shift_in(38) => positive_inputs_11_38_port, 
                           shift_in(37) => positive_inputs_11_37_port, 
                           shift_in(36) => positive_inputs_11_36_port, 
                           shift_in(35) => positive_inputs_11_35_port, 
                           shift_in(34) => positive_inputs_11_34_port, 
                           shift_in(33) => positive_inputs_11_33_port, 
                           shift_in(32) => positive_inputs_11_32_port, 
                           shift_in(31) => positive_inputs_11_31_port, 
                           shift_in(30) => positive_inputs_11_30_port, 
                           shift_in(29) => positive_inputs_11_29_port, 
                           shift_in(28) => positive_inputs_11_28_port, 
                           shift_in(27) => positive_inputs_11_27_port, 
                           shift_in(26) => positive_inputs_11_26_port, 
                           shift_in(25) => positive_inputs_11_25_port, 
                           shift_in(24) => positive_inputs_11_24_port, 
                           shift_in(23) => positive_inputs_11_23_port, 
                           shift_in(22) => positive_inputs_11_22_port, 
                           shift_in(21) => positive_inputs_11_21_port, 
                           shift_in(20) => positive_inputs_11_20_port, 
                           shift_in(19) => positive_inputs_11_19_port, 
                           shift_in(18) => positive_inputs_11_18_port, 
                           shift_in(17) => positive_inputs_11_17_port, 
                           shift_in(16) => positive_inputs_11_16_port, 
                           shift_in(15) => positive_inputs_11_15_port, 
                           shift_in(14) => positive_inputs_11_14_port, 
                           shift_in(13) => positive_inputs_11_13_port, 
                           shift_in(12) => positive_inputs_11_12_port, 
                           shift_in(11) => positive_inputs_11_11_port, 
                           shift_in(10) => positive_inputs_11_10_port, 
                           shift_in(9) => positive_inputs_11_9_port, 
                           shift_in(8) => positive_inputs_11_8_port, 
                           shift_in(7) => positive_inputs_11_7_port, 
                           shift_in(6) => positive_inputs_11_6_port, 
                           shift_in(5) => positive_inputs_11_5_port, 
                           shift_in(4) => positive_inputs_11_4_port, 
                           shift_in(3) => positive_inputs_11_3_port, 
                           shift_in(2) => positive_inputs_11_2_port, 
                           shift_in(1) => positive_inputs_11_1_port, 
                           shift_in(0) => n8, shift_out(63) => 
                           positive_inputs_12_63_port, shift_out(62) => 
                           positive_inputs_12_62_port, shift_out(61) => 
                           positive_inputs_12_61_port, shift_out(60) => 
                           positive_inputs_12_60_port, shift_out(59) => 
                           positive_inputs_12_59_port, shift_out(58) => 
                           positive_inputs_12_58_port, shift_out(57) => 
                           positive_inputs_12_57_port, shift_out(56) => 
                           positive_inputs_12_56_port, shift_out(55) => 
                           positive_inputs_12_55_port, shift_out(54) => 
                           positive_inputs_12_54_port, shift_out(53) => 
                           positive_inputs_12_53_port, shift_out(52) => 
                           positive_inputs_12_52_port, shift_out(51) => 
                           positive_inputs_12_51_port, shift_out(50) => 
                           positive_inputs_12_50_port, shift_out(49) => 
                           positive_inputs_12_49_port, shift_out(48) => 
                           positive_inputs_12_48_port, shift_out(47) => 
                           positive_inputs_12_47_port, shift_out(46) => 
                           positive_inputs_12_46_port, shift_out(45) => 
                           positive_inputs_12_45_port, shift_out(44) => 
                           positive_inputs_12_44_port, shift_out(43) => 
                           positive_inputs_12_43_port, shift_out(42) => 
                           positive_inputs_12_42_port, shift_out(41) => 
                           positive_inputs_12_41_port, shift_out(40) => 
                           positive_inputs_12_40_port, shift_out(39) => 
                           positive_inputs_12_39_port, shift_out(38) => 
                           positive_inputs_12_38_port, shift_out(37) => 
                           positive_inputs_12_37_port, shift_out(36) => 
                           positive_inputs_12_36_port, shift_out(35) => 
                           positive_inputs_12_35_port, shift_out(34) => 
                           positive_inputs_12_34_port, shift_out(33) => 
                           positive_inputs_12_33_port, shift_out(32) => 
                           positive_inputs_12_32_port, shift_out(31) => 
                           positive_inputs_12_31_port, shift_out(30) => 
                           positive_inputs_12_30_port, shift_out(29) => 
                           positive_inputs_12_29_port, shift_out(28) => 
                           positive_inputs_12_28_port, shift_out(27) => 
                           positive_inputs_12_27_port, shift_out(26) => 
                           positive_inputs_12_26_port, shift_out(25) => 
                           positive_inputs_12_25_port, shift_out(24) => 
                           positive_inputs_12_24_port, shift_out(23) => 
                           positive_inputs_12_23_port, shift_out(22) => 
                           positive_inputs_12_22_port, shift_out(21) => 
                           positive_inputs_12_21_port, shift_out(20) => 
                           positive_inputs_12_20_port, shift_out(19) => 
                           positive_inputs_12_19_port, shift_out(18) => 
                           positive_inputs_12_18_port, shift_out(17) => 
                           positive_inputs_12_17_port, shift_out(16) => 
                           positive_inputs_12_16_port, shift_out(15) => 
                           positive_inputs_12_15_port, shift_out(14) => 
                           positive_inputs_12_14_port, shift_out(13) => 
                           positive_inputs_12_13_port, shift_out(12) => 
                           positive_inputs_12_12_port, shift_out(11) => 
                           positive_inputs_12_11_port, shift_out(10) => 
                           positive_inputs_12_10_port, shift_out(9) => 
                           positive_inputs_12_9_port, shift_out(8) => 
                           positive_inputs_12_8_port, shift_out(7) => 
                           positive_inputs_12_7_port, shift_out(6) => 
                           positive_inputs_12_6_port, shift_out(5) => 
                           positive_inputs_12_5_port, shift_out(4) => 
                           positive_inputs_12_4_port, shift_out(3) => 
                           positive_inputs_12_3_port, shift_out(2) => 
                           positive_inputs_12_2_port, shift_out(1) => 
                           positive_inputs_12_1_port, shift_out(0) => n_1012);
   shifted_pos_13 : leftshifter_NbitShifter64_114 port map( shift_in(63) => 
                           positive_inputs_12_63_port, shift_in(62) => 
                           positive_inputs_12_62_port, shift_in(61) => 
                           positive_inputs_12_61_port, shift_in(60) => 
                           positive_inputs_12_60_port, shift_in(59) => 
                           positive_inputs_12_59_port, shift_in(58) => 
                           positive_inputs_12_58_port, shift_in(57) => 
                           positive_inputs_12_57_port, shift_in(56) => 
                           positive_inputs_12_56_port, shift_in(55) => 
                           positive_inputs_12_55_port, shift_in(54) => 
                           positive_inputs_12_54_port, shift_in(53) => 
                           positive_inputs_12_53_port, shift_in(52) => 
                           positive_inputs_12_52_port, shift_in(51) => 
                           positive_inputs_12_51_port, shift_in(50) => 
                           positive_inputs_12_50_port, shift_in(49) => 
                           positive_inputs_12_49_port, shift_in(48) => 
                           positive_inputs_12_48_port, shift_in(47) => n29, 
                           shift_in(46) => positive_inputs_12_46_port, 
                           shift_in(45) => positive_inputs_12_45_port, 
                           shift_in(44) => positive_inputs_12_44_port, 
                           shift_in(43) => positive_inputs_12_43_port, 
                           shift_in(42) => positive_inputs_12_42_port, 
                           shift_in(41) => positive_inputs_12_41_port, 
                           shift_in(40) => positive_inputs_12_40_port, 
                           shift_in(39) => positive_inputs_12_39_port, 
                           shift_in(38) => positive_inputs_12_38_port, 
                           shift_in(37) => positive_inputs_12_37_port, 
                           shift_in(36) => positive_inputs_12_36_port, 
                           shift_in(35) => positive_inputs_12_35_port, 
                           shift_in(34) => positive_inputs_12_34_port, 
                           shift_in(33) => positive_inputs_12_33_port, 
                           shift_in(32) => positive_inputs_12_32_port, 
                           shift_in(31) => positive_inputs_12_31_port, 
                           shift_in(30) => positive_inputs_12_30_port, 
                           shift_in(29) => positive_inputs_12_29_port, 
                           shift_in(28) => positive_inputs_12_28_port, 
                           shift_in(27) => positive_inputs_12_27_port, 
                           shift_in(26) => positive_inputs_12_26_port, 
                           shift_in(25) => positive_inputs_12_25_port, 
                           shift_in(24) => positive_inputs_12_24_port, 
                           shift_in(23) => positive_inputs_12_23_port, 
                           shift_in(22) => positive_inputs_12_22_port, 
                           shift_in(21) => positive_inputs_12_21_port, 
                           shift_in(20) => positive_inputs_12_20_port, 
                           shift_in(19) => positive_inputs_12_19_port, 
                           shift_in(18) => positive_inputs_12_18_port, 
                           shift_in(17) => positive_inputs_12_17_port, 
                           shift_in(16) => positive_inputs_12_16_port, 
                           shift_in(15) => positive_inputs_12_15_port, 
                           shift_in(14) => positive_inputs_12_14_port, 
                           shift_in(13) => positive_inputs_12_13_port, 
                           shift_in(12) => positive_inputs_12_12_port, 
                           shift_in(11) => positive_inputs_12_11_port, 
                           shift_in(10) => positive_inputs_12_10_port, 
                           shift_in(9) => positive_inputs_12_9_port, 
                           shift_in(8) => positive_inputs_12_8_port, 
                           shift_in(7) => positive_inputs_12_7_port, 
                           shift_in(6) => positive_inputs_12_6_port, 
                           shift_in(5) => positive_inputs_12_5_port, 
                           shift_in(4) => positive_inputs_12_4_port, 
                           shift_in(3) => positive_inputs_12_3_port, 
                           shift_in(2) => positive_inputs_12_2_port, 
                           shift_in(1) => positive_inputs_12_1_port, 
                           shift_in(0) => n8, shift_out(63) => 
                           positive_inputs_13_63_port, shift_out(62) => 
                           positive_inputs_13_62_port, shift_out(61) => 
                           positive_inputs_13_61_port, shift_out(60) => 
                           positive_inputs_13_60_port, shift_out(59) => 
                           positive_inputs_13_59_port, shift_out(58) => 
                           positive_inputs_13_58_port, shift_out(57) => 
                           positive_inputs_13_57_port, shift_out(56) => 
                           positive_inputs_13_56_port, shift_out(55) => 
                           positive_inputs_13_55_port, shift_out(54) => 
                           positive_inputs_13_54_port, shift_out(53) => 
                           positive_inputs_13_53_port, shift_out(52) => 
                           positive_inputs_13_52_port, shift_out(51) => 
                           positive_inputs_13_51_port, shift_out(50) => 
                           positive_inputs_13_50_port, shift_out(49) => 
                           positive_inputs_13_49_port, shift_out(48) => 
                           positive_inputs_13_48_port, shift_out(47) => 
                           positive_inputs_13_47_port, shift_out(46) => 
                           positive_inputs_13_46_port, shift_out(45) => 
                           positive_inputs_13_45_port, shift_out(44) => 
                           positive_inputs_13_44_port, shift_out(43) => 
                           positive_inputs_13_43_port, shift_out(42) => 
                           positive_inputs_13_42_port, shift_out(41) => 
                           positive_inputs_13_41_port, shift_out(40) => 
                           positive_inputs_13_40_port, shift_out(39) => 
                           positive_inputs_13_39_port, shift_out(38) => 
                           positive_inputs_13_38_port, shift_out(37) => 
                           positive_inputs_13_37_port, shift_out(36) => 
                           positive_inputs_13_36_port, shift_out(35) => 
                           positive_inputs_13_35_port, shift_out(34) => 
                           positive_inputs_13_34_port, shift_out(33) => 
                           positive_inputs_13_33_port, shift_out(32) => 
                           positive_inputs_13_32_port, shift_out(31) => 
                           positive_inputs_13_31_port, shift_out(30) => 
                           positive_inputs_13_30_port, shift_out(29) => 
                           positive_inputs_13_29_port, shift_out(28) => 
                           positive_inputs_13_28_port, shift_out(27) => 
                           positive_inputs_13_27_port, shift_out(26) => 
                           positive_inputs_13_26_port, shift_out(25) => 
                           positive_inputs_13_25_port, shift_out(24) => 
                           positive_inputs_13_24_port, shift_out(23) => 
                           positive_inputs_13_23_port, shift_out(22) => 
                           positive_inputs_13_22_port, shift_out(21) => 
                           positive_inputs_13_21_port, shift_out(20) => 
                           positive_inputs_13_20_port, shift_out(19) => 
                           positive_inputs_13_19_port, shift_out(18) => 
                           positive_inputs_13_18_port, shift_out(17) => 
                           positive_inputs_13_17_port, shift_out(16) => 
                           positive_inputs_13_16_port, shift_out(15) => 
                           positive_inputs_13_15_port, shift_out(14) => 
                           positive_inputs_13_14_port, shift_out(13) => 
                           positive_inputs_13_13_port, shift_out(12) => 
                           positive_inputs_13_12_port, shift_out(11) => 
                           positive_inputs_13_11_port, shift_out(10) => 
                           positive_inputs_13_10_port, shift_out(9) => 
                           positive_inputs_13_9_port, shift_out(8) => 
                           positive_inputs_13_8_port, shift_out(7) => 
                           positive_inputs_13_7_port, shift_out(6) => 
                           positive_inputs_13_6_port, shift_out(5) => 
                           positive_inputs_13_5_port, shift_out(4) => 
                           positive_inputs_13_4_port, shift_out(3) => 
                           positive_inputs_13_3_port, shift_out(2) => 
                           positive_inputs_13_2_port, shift_out(1) => 
                           positive_inputs_13_1_port, shift_out(0) => n_1013);
   shifted_pos_14 : leftshifter_NbitShifter64_113 port map( shift_in(63) => 
                           positive_inputs_13_63_port, shift_in(62) => 
                           positive_inputs_13_62_port, shift_in(61) => 
                           positive_inputs_13_61_port, shift_in(60) => 
                           positive_inputs_13_60_port, shift_in(59) => 
                           positive_inputs_13_59_port, shift_in(58) => 
                           positive_inputs_13_58_port, shift_in(57) => 
                           positive_inputs_13_57_port, shift_in(56) => 
                           positive_inputs_13_56_port, shift_in(55) => 
                           positive_inputs_13_55_port, shift_in(54) => 
                           positive_inputs_13_54_port, shift_in(53) => 
                           positive_inputs_13_53_port, shift_in(52) => 
                           positive_inputs_13_52_port, shift_in(51) => 
                           positive_inputs_13_51_port, shift_in(50) => 
                           positive_inputs_13_50_port, shift_in(49) => 
                           positive_inputs_13_49_port, shift_in(48) => 
                           positive_inputs_13_48_port, shift_in(47) => n28, 
                           shift_in(46) => positive_inputs_13_46_port, 
                           shift_in(45) => positive_inputs_13_45_port, 
                           shift_in(44) => positive_inputs_13_44_port, 
                           shift_in(43) => positive_inputs_13_43_port, 
                           shift_in(42) => positive_inputs_13_42_port, 
                           shift_in(41) => positive_inputs_13_41_port, 
                           shift_in(40) => positive_inputs_13_40_port, 
                           shift_in(39) => positive_inputs_13_39_port, 
                           shift_in(38) => positive_inputs_13_38_port, 
                           shift_in(37) => positive_inputs_13_37_port, 
                           shift_in(36) => positive_inputs_13_36_port, 
                           shift_in(35) => positive_inputs_13_35_port, 
                           shift_in(34) => positive_inputs_13_34_port, 
                           shift_in(33) => positive_inputs_13_33_port, 
                           shift_in(32) => positive_inputs_13_32_port, 
                           shift_in(31) => positive_inputs_13_31_port, 
                           shift_in(30) => positive_inputs_13_30_port, 
                           shift_in(29) => positive_inputs_13_29_port, 
                           shift_in(28) => positive_inputs_13_28_port, 
                           shift_in(27) => positive_inputs_13_27_port, 
                           shift_in(26) => positive_inputs_13_26_port, 
                           shift_in(25) => positive_inputs_13_25_port, 
                           shift_in(24) => positive_inputs_13_24_port, 
                           shift_in(23) => positive_inputs_13_23_port, 
                           shift_in(22) => positive_inputs_13_22_port, 
                           shift_in(21) => positive_inputs_13_21_port, 
                           shift_in(20) => positive_inputs_13_20_port, 
                           shift_in(19) => positive_inputs_13_19_port, 
                           shift_in(18) => positive_inputs_13_18_port, 
                           shift_in(17) => positive_inputs_13_17_port, 
                           shift_in(16) => positive_inputs_13_16_port, 
                           shift_in(15) => positive_inputs_13_15_port, 
                           shift_in(14) => positive_inputs_13_14_port, 
                           shift_in(13) => positive_inputs_13_13_port, 
                           shift_in(12) => positive_inputs_13_12_port, 
                           shift_in(11) => positive_inputs_13_11_port, 
                           shift_in(10) => positive_inputs_13_10_port, 
                           shift_in(9) => positive_inputs_13_9_port, 
                           shift_in(8) => positive_inputs_13_8_port, 
                           shift_in(7) => positive_inputs_13_7_port, 
                           shift_in(6) => positive_inputs_13_6_port, 
                           shift_in(5) => positive_inputs_13_5_port, 
                           shift_in(4) => positive_inputs_13_4_port, 
                           shift_in(3) => positive_inputs_13_3_port, 
                           shift_in(2) => positive_inputs_13_2_port, 
                           shift_in(1) => positive_inputs_13_1_port, 
                           shift_in(0) => n8, shift_out(63) => 
                           positive_inputs_14_63_port, shift_out(62) => 
                           positive_inputs_14_62_port, shift_out(61) => 
                           positive_inputs_14_61_port, shift_out(60) => 
                           positive_inputs_14_60_port, shift_out(59) => 
                           positive_inputs_14_59_port, shift_out(58) => 
                           positive_inputs_14_58_port, shift_out(57) => 
                           positive_inputs_14_57_port, shift_out(56) => 
                           positive_inputs_14_56_port, shift_out(55) => 
                           positive_inputs_14_55_port, shift_out(54) => 
                           positive_inputs_14_54_port, shift_out(53) => 
                           positive_inputs_14_53_port, shift_out(52) => 
                           positive_inputs_14_52_port, shift_out(51) => 
                           positive_inputs_14_51_port, shift_out(50) => 
                           positive_inputs_14_50_port, shift_out(49) => 
                           positive_inputs_14_49_port, shift_out(48) => 
                           positive_inputs_14_48_port, shift_out(47) => 
                           positive_inputs_14_47_port, shift_out(46) => 
                           positive_inputs_14_46_port, shift_out(45) => 
                           positive_inputs_14_45_port, shift_out(44) => 
                           positive_inputs_14_44_port, shift_out(43) => 
                           positive_inputs_14_43_port, shift_out(42) => 
                           positive_inputs_14_42_port, shift_out(41) => 
                           positive_inputs_14_41_port, shift_out(40) => 
                           positive_inputs_14_40_port, shift_out(39) => 
                           positive_inputs_14_39_port, shift_out(38) => 
                           positive_inputs_14_38_port, shift_out(37) => 
                           positive_inputs_14_37_port, shift_out(36) => 
                           positive_inputs_14_36_port, shift_out(35) => 
                           positive_inputs_14_35_port, shift_out(34) => 
                           positive_inputs_14_34_port, shift_out(33) => 
                           positive_inputs_14_33_port, shift_out(32) => 
                           positive_inputs_14_32_port, shift_out(31) => 
                           positive_inputs_14_31_port, shift_out(30) => 
                           positive_inputs_14_30_port, shift_out(29) => 
                           positive_inputs_14_29_port, shift_out(28) => 
                           positive_inputs_14_28_port, shift_out(27) => 
                           positive_inputs_14_27_port, shift_out(26) => 
                           positive_inputs_14_26_port, shift_out(25) => 
                           positive_inputs_14_25_port, shift_out(24) => 
                           positive_inputs_14_24_port, shift_out(23) => 
                           positive_inputs_14_23_port, shift_out(22) => 
                           positive_inputs_14_22_port, shift_out(21) => 
                           positive_inputs_14_21_port, shift_out(20) => 
                           positive_inputs_14_20_port, shift_out(19) => 
                           positive_inputs_14_19_port, shift_out(18) => 
                           positive_inputs_14_18_port, shift_out(17) => 
                           positive_inputs_14_17_port, shift_out(16) => 
                           positive_inputs_14_16_port, shift_out(15) => 
                           positive_inputs_14_15_port, shift_out(14) => 
                           positive_inputs_14_14_port, shift_out(13) => 
                           positive_inputs_14_13_port, shift_out(12) => 
                           positive_inputs_14_12_port, shift_out(11) => 
                           positive_inputs_14_11_port, shift_out(10) => 
                           positive_inputs_14_10_port, shift_out(9) => 
                           positive_inputs_14_9_port, shift_out(8) => 
                           positive_inputs_14_8_port, shift_out(7) => 
                           positive_inputs_14_7_port, shift_out(6) => 
                           positive_inputs_14_6_port, shift_out(5) => 
                           positive_inputs_14_5_port, shift_out(4) => 
                           positive_inputs_14_4_port, shift_out(3) => 
                           positive_inputs_14_3_port, shift_out(2) => 
                           positive_inputs_14_2_port, shift_out(1) => 
                           positive_inputs_14_1_port, shift_out(0) => n_1014);
   shifted_pos_15 : leftshifter_NbitShifter64_112 port map( shift_in(63) => 
                           positive_inputs_14_63_port, shift_in(62) => 
                           positive_inputs_14_62_port, shift_in(61) => 
                           positive_inputs_14_61_port, shift_in(60) => 
                           positive_inputs_14_60_port, shift_in(59) => 
                           positive_inputs_14_59_port, shift_in(58) => 
                           positive_inputs_14_58_port, shift_in(57) => 
                           positive_inputs_14_57_port, shift_in(56) => 
                           positive_inputs_14_56_port, shift_in(55) => 
                           positive_inputs_14_55_port, shift_in(54) => 
                           positive_inputs_14_54_port, shift_in(53) => 
                           positive_inputs_14_53_port, shift_in(52) => 
                           positive_inputs_14_52_port, shift_in(51) => 
                           positive_inputs_14_51_port, shift_in(50) => 
                           positive_inputs_14_50_port, shift_in(49) => 
                           positive_inputs_14_49_port, shift_in(48) => 
                           positive_inputs_14_48_port, shift_in(47) => n27, 
                           shift_in(46) => positive_inputs_14_46_port, 
                           shift_in(45) => positive_inputs_14_45_port, 
                           shift_in(44) => positive_inputs_14_44_port, 
                           shift_in(43) => positive_inputs_14_43_port, 
                           shift_in(42) => positive_inputs_14_42_port, 
                           shift_in(41) => positive_inputs_14_41_port, 
                           shift_in(40) => positive_inputs_14_40_port, 
                           shift_in(39) => positive_inputs_14_39_port, 
                           shift_in(38) => positive_inputs_14_38_port, 
                           shift_in(37) => positive_inputs_14_37_port, 
                           shift_in(36) => positive_inputs_14_36_port, 
                           shift_in(35) => positive_inputs_14_35_port, 
                           shift_in(34) => positive_inputs_14_34_port, 
                           shift_in(33) => positive_inputs_14_33_port, 
                           shift_in(32) => positive_inputs_14_32_port, 
                           shift_in(31) => positive_inputs_14_31_port, 
                           shift_in(30) => positive_inputs_14_30_port, 
                           shift_in(29) => positive_inputs_14_29_port, 
                           shift_in(28) => positive_inputs_14_28_port, 
                           shift_in(27) => positive_inputs_14_27_port, 
                           shift_in(26) => positive_inputs_14_26_port, 
                           shift_in(25) => positive_inputs_14_25_port, 
                           shift_in(24) => positive_inputs_14_24_port, 
                           shift_in(23) => positive_inputs_14_23_port, 
                           shift_in(22) => positive_inputs_14_22_port, 
                           shift_in(21) => positive_inputs_14_21_port, 
                           shift_in(20) => positive_inputs_14_20_port, 
                           shift_in(19) => positive_inputs_14_19_port, 
                           shift_in(18) => positive_inputs_14_18_port, 
                           shift_in(17) => positive_inputs_14_17_port, 
                           shift_in(16) => positive_inputs_14_16_port, 
                           shift_in(15) => positive_inputs_14_15_port, 
                           shift_in(14) => positive_inputs_14_14_port, 
                           shift_in(13) => positive_inputs_14_13_port, 
                           shift_in(12) => positive_inputs_14_12_port, 
                           shift_in(11) => positive_inputs_14_11_port, 
                           shift_in(10) => positive_inputs_14_10_port, 
                           shift_in(9) => positive_inputs_14_9_port, 
                           shift_in(8) => positive_inputs_14_8_port, 
                           shift_in(7) => positive_inputs_14_7_port, 
                           shift_in(6) => positive_inputs_14_6_port, 
                           shift_in(5) => positive_inputs_14_5_port, 
                           shift_in(4) => positive_inputs_14_4_port, 
                           shift_in(3) => positive_inputs_14_3_port, 
                           shift_in(2) => positive_inputs_14_2_port, 
                           shift_in(1) => positive_inputs_14_1_port, 
                           shift_in(0) => n8, shift_out(63) => 
                           positive_inputs_15_63_port, shift_out(62) => 
                           positive_inputs_15_62_port, shift_out(61) => 
                           positive_inputs_15_61_port, shift_out(60) => 
                           positive_inputs_15_60_port, shift_out(59) => 
                           positive_inputs_15_59_port, shift_out(58) => 
                           positive_inputs_15_58_port, shift_out(57) => 
                           positive_inputs_15_57_port, shift_out(56) => 
                           positive_inputs_15_56_port, shift_out(55) => 
                           positive_inputs_15_55_port, shift_out(54) => 
                           positive_inputs_15_54_port, shift_out(53) => 
                           positive_inputs_15_53_port, shift_out(52) => 
                           positive_inputs_15_52_port, shift_out(51) => 
                           positive_inputs_15_51_port, shift_out(50) => 
                           positive_inputs_15_50_port, shift_out(49) => 
                           positive_inputs_15_49_port, shift_out(48) => 
                           positive_inputs_15_48_port, shift_out(47) => 
                           positive_inputs_15_47_port, shift_out(46) => 
                           positive_inputs_15_46_port, shift_out(45) => 
                           positive_inputs_15_45_port, shift_out(44) => 
                           positive_inputs_15_44_port, shift_out(43) => 
                           positive_inputs_15_43_port, shift_out(42) => 
                           positive_inputs_15_42_port, shift_out(41) => 
                           positive_inputs_15_41_port, shift_out(40) => 
                           positive_inputs_15_40_port, shift_out(39) => 
                           positive_inputs_15_39_port, shift_out(38) => 
                           positive_inputs_15_38_port, shift_out(37) => 
                           positive_inputs_15_37_port, shift_out(36) => 
                           positive_inputs_15_36_port, shift_out(35) => 
                           positive_inputs_15_35_port, shift_out(34) => 
                           positive_inputs_15_34_port, shift_out(33) => 
                           positive_inputs_15_33_port, shift_out(32) => 
                           positive_inputs_15_32_port, shift_out(31) => 
                           positive_inputs_15_31_port, shift_out(30) => 
                           positive_inputs_15_30_port, shift_out(29) => 
                           positive_inputs_15_29_port, shift_out(28) => 
                           positive_inputs_15_28_port, shift_out(27) => 
                           positive_inputs_15_27_port, shift_out(26) => 
                           positive_inputs_15_26_port, shift_out(25) => 
                           positive_inputs_15_25_port, shift_out(24) => 
                           positive_inputs_15_24_port, shift_out(23) => 
                           positive_inputs_15_23_port, shift_out(22) => 
                           positive_inputs_15_22_port, shift_out(21) => 
                           positive_inputs_15_21_port, shift_out(20) => 
                           positive_inputs_15_20_port, shift_out(19) => 
                           positive_inputs_15_19_port, shift_out(18) => 
                           positive_inputs_15_18_port, shift_out(17) => 
                           positive_inputs_15_17_port, shift_out(16) => 
                           positive_inputs_15_16_port, shift_out(15) => 
                           positive_inputs_15_15_port, shift_out(14) => 
                           positive_inputs_15_14_port, shift_out(13) => 
                           positive_inputs_15_13_port, shift_out(12) => 
                           positive_inputs_15_12_port, shift_out(11) => 
                           positive_inputs_15_11_port, shift_out(10) => 
                           positive_inputs_15_10_port, shift_out(9) => 
                           positive_inputs_15_9_port, shift_out(8) => 
                           positive_inputs_15_8_port, shift_out(7) => 
                           positive_inputs_15_7_port, shift_out(6) => 
                           positive_inputs_15_6_port, shift_out(5) => 
                           positive_inputs_15_5_port, shift_out(4) => 
                           positive_inputs_15_4_port, shift_out(3) => 
                           positive_inputs_15_3_port, shift_out(2) => 
                           positive_inputs_15_2_port, shift_out(1) => 
                           positive_inputs_15_1_port, shift_out(0) => n_1015);
   shifted_pos_16 : leftshifter_NbitShifter64_111 port map( shift_in(63) => 
                           positive_inputs_15_63_port, shift_in(62) => 
                           positive_inputs_15_62_port, shift_in(61) => 
                           positive_inputs_15_61_port, shift_in(60) => 
                           positive_inputs_15_60_port, shift_in(59) => 
                           positive_inputs_15_59_port, shift_in(58) => 
                           positive_inputs_15_58_port, shift_in(57) => 
                           positive_inputs_15_57_port, shift_in(56) => 
                           positive_inputs_15_56_port, shift_in(55) => 
                           positive_inputs_15_55_port, shift_in(54) => 
                           positive_inputs_15_54_port, shift_in(53) => 
                           positive_inputs_15_53_port, shift_in(52) => 
                           positive_inputs_15_52_port, shift_in(51) => 
                           positive_inputs_15_51_port, shift_in(50) => 
                           positive_inputs_15_50_port, shift_in(49) => 
                           positive_inputs_15_49_port, shift_in(48) => 
                           positive_inputs_15_48_port, shift_in(47) => n26, 
                           shift_in(46) => n25, shift_in(45) => n181, 
                           shift_in(44) => n179, shift_in(43) => n177, 
                           shift_in(42) => n175, shift_in(41) => n173, 
                           shift_in(40) => n171, shift_in(39) => n169, 
                           shift_in(38) => n167, shift_in(37) => n165, 
                           shift_in(36) => n163, shift_in(35) => n161, 
                           shift_in(34) => n159, shift_in(33) => n157, 
                           shift_in(32) => n155, shift_in(31) => n153, 
                           shift_in(30) => n151, shift_in(29) => n149, 
                           shift_in(28) => n147, shift_in(27) => n145, 
                           shift_in(26) => n143, shift_in(25) => n141, 
                           shift_in(24) => n139, shift_in(23) => n137, 
                           shift_in(22) => n135, shift_in(21) => n133, 
                           shift_in(20) => n131, shift_in(19) => n129, 
                           shift_in(18) => n127, shift_in(17) => n125, 
                           shift_in(16) => n123, shift_in(15) => n121, 
                           shift_in(14) => positive_inputs_15_14_port, 
                           shift_in(13) => positive_inputs_15_13_port, 
                           shift_in(12) => positive_inputs_15_12_port, 
                           shift_in(11) => positive_inputs_15_11_port, 
                           shift_in(10) => positive_inputs_15_10_port, 
                           shift_in(9) => positive_inputs_15_9_port, 
                           shift_in(8) => positive_inputs_15_8_port, 
                           shift_in(7) => positive_inputs_15_7_port, 
                           shift_in(6) => positive_inputs_15_6_port, 
                           shift_in(5) => positive_inputs_15_5_port, 
                           shift_in(4) => positive_inputs_15_4_port, 
                           shift_in(3) => positive_inputs_15_3_port, 
                           shift_in(2) => positive_inputs_15_2_port, 
                           shift_in(1) => positive_inputs_15_1_port, 
                           shift_in(0) => n8, shift_out(63) => 
                           positive_inputs_16_63_port, shift_out(62) => 
                           positive_inputs_16_62_port, shift_out(61) => 
                           positive_inputs_16_61_port, shift_out(60) => 
                           positive_inputs_16_60_port, shift_out(59) => 
                           positive_inputs_16_59_port, shift_out(58) => 
                           positive_inputs_16_58_port, shift_out(57) => 
                           positive_inputs_16_57_port, shift_out(56) => 
                           positive_inputs_16_56_port, shift_out(55) => 
                           positive_inputs_16_55_port, shift_out(54) => 
                           positive_inputs_16_54_port, shift_out(53) => 
                           positive_inputs_16_53_port, shift_out(52) => 
                           positive_inputs_16_52_port, shift_out(51) => 
                           positive_inputs_16_51_port, shift_out(50) => 
                           positive_inputs_16_50_port, shift_out(49) => 
                           positive_inputs_16_49_port, shift_out(48) => 
                           positive_inputs_16_48_port, shift_out(47) => 
                           positive_inputs_16_47_port, shift_out(46) => 
                           positive_inputs_16_46_port, shift_out(45) => 
                           positive_inputs_16_45_port, shift_out(44) => 
                           positive_inputs_16_44_port, shift_out(43) => 
                           positive_inputs_16_43_port, shift_out(42) => 
                           positive_inputs_16_42_port, shift_out(41) => 
                           positive_inputs_16_41_port, shift_out(40) => 
                           positive_inputs_16_40_port, shift_out(39) => 
                           positive_inputs_16_39_port, shift_out(38) => 
                           positive_inputs_16_38_port, shift_out(37) => 
                           positive_inputs_16_37_port, shift_out(36) => 
                           positive_inputs_16_36_port, shift_out(35) => 
                           positive_inputs_16_35_port, shift_out(34) => 
                           positive_inputs_16_34_port, shift_out(33) => 
                           positive_inputs_16_33_port, shift_out(32) => 
                           positive_inputs_16_32_port, shift_out(31) => 
                           positive_inputs_16_31_port, shift_out(30) => 
                           positive_inputs_16_30_port, shift_out(29) => 
                           positive_inputs_16_29_port, shift_out(28) => 
                           positive_inputs_16_28_port, shift_out(27) => 
                           positive_inputs_16_27_port, shift_out(26) => 
                           positive_inputs_16_26_port, shift_out(25) => 
                           positive_inputs_16_25_port, shift_out(24) => 
                           positive_inputs_16_24_port, shift_out(23) => 
                           positive_inputs_16_23_port, shift_out(22) => 
                           positive_inputs_16_22_port, shift_out(21) => 
                           positive_inputs_16_21_port, shift_out(20) => 
                           positive_inputs_16_20_port, shift_out(19) => 
                           positive_inputs_16_19_port, shift_out(18) => 
                           positive_inputs_16_18_port, shift_out(17) => 
                           positive_inputs_16_17_port, shift_out(16) => 
                           positive_inputs_16_16_port, shift_out(15) => 
                           positive_inputs_16_15_port, shift_out(14) => 
                           positive_inputs_16_14_port, shift_out(13) => 
                           positive_inputs_16_13_port, shift_out(12) => 
                           positive_inputs_16_12_port, shift_out(11) => 
                           positive_inputs_16_11_port, shift_out(10) => 
                           positive_inputs_16_10_port, shift_out(9) => 
                           positive_inputs_16_9_port, shift_out(8) => 
                           positive_inputs_16_8_port, shift_out(7) => 
                           positive_inputs_16_7_port, shift_out(6) => 
                           positive_inputs_16_6_port, shift_out(5) => 
                           positive_inputs_16_5_port, shift_out(4) => 
                           positive_inputs_16_4_port, shift_out(3) => 
                           positive_inputs_16_3_port, shift_out(2) => 
                           positive_inputs_16_2_port, shift_out(1) => 
                           positive_inputs_16_1_port, shift_out(0) => n_1016);
   shifted_pos_17 : leftshifter_NbitShifter64_110 port map( shift_in(63) => 
                           positive_inputs_16_63_port, shift_in(62) => 
                           positive_inputs_16_62_port, shift_in(61) => 
                           positive_inputs_16_61_port, shift_in(60) => 
                           positive_inputs_16_60_port, shift_in(59) => 
                           positive_inputs_16_59_port, shift_in(58) => 
                           positive_inputs_16_58_port, shift_in(57) => 
                           positive_inputs_16_57_port, shift_in(56) => 
                           positive_inputs_16_56_port, shift_in(55) => 
                           positive_inputs_16_55_port, shift_in(54) => 
                           positive_inputs_16_54_port, shift_in(53) => 
                           positive_inputs_16_53_port, shift_in(52) => 
                           positive_inputs_16_52_port, shift_in(51) => 
                           positive_inputs_16_51_port, shift_in(50) => 
                           positive_inputs_16_50_port, shift_in(49) => 
                           positive_inputs_16_49_port, shift_in(48) => 
                           positive_inputs_16_48_port, shift_in(47) => 
                           positive_inputs_16_47_port, shift_in(46) => 
                           positive_inputs_16_46_port, shift_in(45) => 
                           positive_inputs_16_45_port, shift_in(44) => 
                           positive_inputs_16_44_port, shift_in(43) => 
                           positive_inputs_16_43_port, shift_in(42) => 
                           positive_inputs_16_42_port, shift_in(41) => 
                           positive_inputs_16_41_port, shift_in(40) => 
                           positive_inputs_16_40_port, shift_in(39) => 
                           positive_inputs_16_39_port, shift_in(38) => 
                           positive_inputs_16_38_port, shift_in(37) => 
                           positive_inputs_16_37_port, shift_in(36) => 
                           positive_inputs_16_36_port, shift_in(35) => 
                           positive_inputs_16_35_port, shift_in(34) => 
                           positive_inputs_16_34_port, shift_in(33) => 
                           positive_inputs_16_33_port, shift_in(32) => 
                           positive_inputs_16_32_port, shift_in(31) => 
                           positive_inputs_16_31_port, shift_in(30) => 
                           positive_inputs_16_30_port, shift_in(29) => 
                           positive_inputs_16_29_port, shift_in(28) => 
                           positive_inputs_16_28_port, shift_in(27) => 
                           positive_inputs_16_27_port, shift_in(26) => 
                           positive_inputs_16_26_port, shift_in(25) => 
                           positive_inputs_16_25_port, shift_in(24) => 
                           positive_inputs_16_24_port, shift_in(23) => 
                           positive_inputs_16_23_port, shift_in(22) => 
                           positive_inputs_16_22_port, shift_in(21) => 
                           positive_inputs_16_21_port, shift_in(20) => 
                           positive_inputs_16_20_port, shift_in(19) => 
                           positive_inputs_16_19_port, shift_in(18) => 
                           positive_inputs_16_18_port, shift_in(17) => 
                           positive_inputs_16_17_port, shift_in(16) => 
                           positive_inputs_16_16_port, shift_in(15) => 
                           positive_inputs_16_15_port, shift_in(14) => 
                           positive_inputs_16_14_port, shift_in(13) => 
                           positive_inputs_16_13_port, shift_in(12) => 
                           positive_inputs_16_12_port, shift_in(11) => 
                           positive_inputs_16_11_port, shift_in(10) => 
                           positive_inputs_16_10_port, shift_in(9) => 
                           positive_inputs_16_9_port, shift_in(8) => 
                           positive_inputs_16_8_port, shift_in(7) => 
                           positive_inputs_16_7_port, shift_in(6) => 
                           positive_inputs_16_6_port, shift_in(5) => 
                           positive_inputs_16_5_port, shift_in(4) => 
                           positive_inputs_16_4_port, shift_in(3) => 
                           positive_inputs_16_3_port, shift_in(2) => 
                           positive_inputs_16_2_port, shift_in(1) => 
                           positive_inputs_16_1_port, shift_in(0) => n8, 
                           shift_out(63) => positive_inputs_17_63_port, 
                           shift_out(62) => positive_inputs_17_62_port, 
                           shift_out(61) => positive_inputs_17_61_port, 
                           shift_out(60) => positive_inputs_17_60_port, 
                           shift_out(59) => positive_inputs_17_59_port, 
                           shift_out(58) => positive_inputs_17_58_port, 
                           shift_out(57) => positive_inputs_17_57_port, 
                           shift_out(56) => positive_inputs_17_56_port, 
                           shift_out(55) => positive_inputs_17_55_port, 
                           shift_out(54) => positive_inputs_17_54_port, 
                           shift_out(53) => positive_inputs_17_53_port, 
                           shift_out(52) => positive_inputs_17_52_port, 
                           shift_out(51) => positive_inputs_17_51_port, 
                           shift_out(50) => positive_inputs_17_50_port, 
                           shift_out(49) => positive_inputs_17_49_port, 
                           shift_out(48) => positive_inputs_17_48_port, 
                           shift_out(47) => positive_inputs_17_47_port, 
                           shift_out(46) => positive_inputs_17_46_port, 
                           shift_out(45) => positive_inputs_17_45_port, 
                           shift_out(44) => positive_inputs_17_44_port, 
                           shift_out(43) => positive_inputs_17_43_port, 
                           shift_out(42) => positive_inputs_17_42_port, 
                           shift_out(41) => positive_inputs_17_41_port, 
                           shift_out(40) => positive_inputs_17_40_port, 
                           shift_out(39) => positive_inputs_17_39_port, 
                           shift_out(38) => positive_inputs_17_38_port, 
                           shift_out(37) => positive_inputs_17_37_port, 
                           shift_out(36) => positive_inputs_17_36_port, 
                           shift_out(35) => positive_inputs_17_35_port, 
                           shift_out(34) => positive_inputs_17_34_port, 
                           shift_out(33) => positive_inputs_17_33_port, 
                           shift_out(32) => positive_inputs_17_32_port, 
                           shift_out(31) => positive_inputs_17_31_port, 
                           shift_out(30) => positive_inputs_17_30_port, 
                           shift_out(29) => positive_inputs_17_29_port, 
                           shift_out(28) => positive_inputs_17_28_port, 
                           shift_out(27) => positive_inputs_17_27_port, 
                           shift_out(26) => positive_inputs_17_26_port, 
                           shift_out(25) => positive_inputs_17_25_port, 
                           shift_out(24) => positive_inputs_17_24_port, 
                           shift_out(23) => positive_inputs_17_23_port, 
                           shift_out(22) => positive_inputs_17_22_port, 
                           shift_out(21) => positive_inputs_17_21_port, 
                           shift_out(20) => positive_inputs_17_20_port, 
                           shift_out(19) => positive_inputs_17_19_port, 
                           shift_out(18) => positive_inputs_17_18_port, 
                           shift_out(17) => positive_inputs_17_17_port, 
                           shift_out(16) => positive_inputs_17_16_port, 
                           shift_out(15) => positive_inputs_17_15_port, 
                           shift_out(14) => positive_inputs_17_14_port, 
                           shift_out(13) => positive_inputs_17_13_port, 
                           shift_out(12) => positive_inputs_17_12_port, 
                           shift_out(11) => positive_inputs_17_11_port, 
                           shift_out(10) => positive_inputs_17_10_port, 
                           shift_out(9) => positive_inputs_17_9_port, 
                           shift_out(8) => positive_inputs_17_8_port, 
                           shift_out(7) => positive_inputs_17_7_port, 
                           shift_out(6) => positive_inputs_17_6_port, 
                           shift_out(5) => positive_inputs_17_5_port, 
                           shift_out(4) => positive_inputs_17_4_port, 
                           shift_out(3) => positive_inputs_17_3_port, 
                           shift_out(2) => positive_inputs_17_2_port, 
                           shift_out(1) => positive_inputs_17_1_port, 
                           shift_out(0) => n_1017);
   shifted_pos_18 : leftshifter_NbitShifter64_109 port map( shift_in(63) => 
                           positive_inputs_17_63_port, shift_in(62) => 
                           positive_inputs_17_62_port, shift_in(61) => 
                           positive_inputs_17_61_port, shift_in(60) => 
                           positive_inputs_17_60_port, shift_in(59) => 
                           positive_inputs_17_59_port, shift_in(58) => 
                           positive_inputs_17_58_port, shift_in(57) => 
                           positive_inputs_17_57_port, shift_in(56) => 
                           positive_inputs_17_56_port, shift_in(55) => 
                           positive_inputs_17_55_port, shift_in(54) => 
                           positive_inputs_17_54_port, shift_in(53) => 
                           positive_inputs_17_53_port, shift_in(52) => 
                           positive_inputs_17_52_port, shift_in(51) => 
                           positive_inputs_17_51_port, shift_in(50) => 
                           positive_inputs_17_50_port, shift_in(49) => 
                           positive_inputs_17_49_port, shift_in(48) => 
                           positive_inputs_17_48_port, shift_in(47) => 
                           positive_inputs_17_47_port, shift_in(46) => 
                           positive_inputs_17_46_port, shift_in(45) => 
                           positive_inputs_17_45_port, shift_in(44) => 
                           positive_inputs_17_44_port, shift_in(43) => 
                           positive_inputs_17_43_port, shift_in(42) => 
                           positive_inputs_17_42_port, shift_in(41) => 
                           positive_inputs_17_41_port, shift_in(40) => 
                           positive_inputs_17_40_port, shift_in(39) => 
                           positive_inputs_17_39_port, shift_in(38) => 
                           positive_inputs_17_38_port, shift_in(37) => 
                           positive_inputs_17_37_port, shift_in(36) => 
                           positive_inputs_17_36_port, shift_in(35) => 
                           positive_inputs_17_35_port, shift_in(34) => 
                           positive_inputs_17_34_port, shift_in(33) => 
                           positive_inputs_17_33_port, shift_in(32) => 
                           positive_inputs_17_32_port, shift_in(31) => 
                           positive_inputs_17_31_port, shift_in(30) => 
                           positive_inputs_17_30_port, shift_in(29) => 
                           positive_inputs_17_29_port, shift_in(28) => 
                           positive_inputs_17_28_port, shift_in(27) => 
                           positive_inputs_17_27_port, shift_in(26) => 
                           positive_inputs_17_26_port, shift_in(25) => 
                           positive_inputs_17_25_port, shift_in(24) => 
                           positive_inputs_17_24_port, shift_in(23) => 
                           positive_inputs_17_23_port, shift_in(22) => 
                           positive_inputs_17_22_port, shift_in(21) => 
                           positive_inputs_17_21_port, shift_in(20) => 
                           positive_inputs_17_20_port, shift_in(19) => 
                           positive_inputs_17_19_port, shift_in(18) => 
                           positive_inputs_17_18_port, shift_in(17) => 
                           positive_inputs_17_17_port, shift_in(16) => 
                           positive_inputs_17_16_port, shift_in(15) => 
                           positive_inputs_17_15_port, shift_in(14) => 
                           positive_inputs_17_14_port, shift_in(13) => 
                           positive_inputs_17_13_port, shift_in(12) => 
                           positive_inputs_17_12_port, shift_in(11) => 
                           positive_inputs_17_11_port, shift_in(10) => 
                           positive_inputs_17_10_port, shift_in(9) => 
                           positive_inputs_17_9_port, shift_in(8) => 
                           positive_inputs_17_8_port, shift_in(7) => 
                           positive_inputs_17_7_port, shift_in(6) => 
                           positive_inputs_17_6_port, shift_in(5) => 
                           positive_inputs_17_5_port, shift_in(4) => 
                           positive_inputs_17_4_port, shift_in(3) => 
                           positive_inputs_17_3_port, shift_in(2) => 
                           positive_inputs_17_2_port, shift_in(1) => 
                           positive_inputs_17_1_port, shift_in(0) => n8, 
                           shift_out(63) => positive_inputs_18_63_port, 
                           shift_out(62) => positive_inputs_18_62_port, 
                           shift_out(61) => positive_inputs_18_61_port, 
                           shift_out(60) => positive_inputs_18_60_port, 
                           shift_out(59) => positive_inputs_18_59_port, 
                           shift_out(58) => positive_inputs_18_58_port, 
                           shift_out(57) => positive_inputs_18_57_port, 
                           shift_out(56) => positive_inputs_18_56_port, 
                           shift_out(55) => positive_inputs_18_55_port, 
                           shift_out(54) => positive_inputs_18_54_port, 
                           shift_out(53) => positive_inputs_18_53_port, 
                           shift_out(52) => positive_inputs_18_52_port, 
                           shift_out(51) => positive_inputs_18_51_port, 
                           shift_out(50) => positive_inputs_18_50_port, 
                           shift_out(49) => positive_inputs_18_49_port, 
                           shift_out(48) => positive_inputs_18_48_port, 
                           shift_out(47) => positive_inputs_18_47_port, 
                           shift_out(46) => positive_inputs_18_46_port, 
                           shift_out(45) => positive_inputs_18_45_port, 
                           shift_out(44) => positive_inputs_18_44_port, 
                           shift_out(43) => positive_inputs_18_43_port, 
                           shift_out(42) => positive_inputs_18_42_port, 
                           shift_out(41) => positive_inputs_18_41_port, 
                           shift_out(40) => positive_inputs_18_40_port, 
                           shift_out(39) => positive_inputs_18_39_port, 
                           shift_out(38) => positive_inputs_18_38_port, 
                           shift_out(37) => positive_inputs_18_37_port, 
                           shift_out(36) => positive_inputs_18_36_port, 
                           shift_out(35) => positive_inputs_18_35_port, 
                           shift_out(34) => positive_inputs_18_34_port, 
                           shift_out(33) => positive_inputs_18_33_port, 
                           shift_out(32) => positive_inputs_18_32_port, 
                           shift_out(31) => positive_inputs_18_31_port, 
                           shift_out(30) => positive_inputs_18_30_port, 
                           shift_out(29) => positive_inputs_18_29_port, 
                           shift_out(28) => positive_inputs_18_28_port, 
                           shift_out(27) => positive_inputs_18_27_port, 
                           shift_out(26) => positive_inputs_18_26_port, 
                           shift_out(25) => positive_inputs_18_25_port, 
                           shift_out(24) => positive_inputs_18_24_port, 
                           shift_out(23) => positive_inputs_18_23_port, 
                           shift_out(22) => positive_inputs_18_22_port, 
                           shift_out(21) => positive_inputs_18_21_port, 
                           shift_out(20) => positive_inputs_18_20_port, 
                           shift_out(19) => positive_inputs_18_19_port, 
                           shift_out(18) => positive_inputs_18_18_port, 
                           shift_out(17) => positive_inputs_18_17_port, 
                           shift_out(16) => positive_inputs_18_16_port, 
                           shift_out(15) => positive_inputs_18_15_port, 
                           shift_out(14) => positive_inputs_18_14_port, 
                           shift_out(13) => positive_inputs_18_13_port, 
                           shift_out(12) => positive_inputs_18_12_port, 
                           shift_out(11) => positive_inputs_18_11_port, 
                           shift_out(10) => positive_inputs_18_10_port, 
                           shift_out(9) => positive_inputs_18_9_port, 
                           shift_out(8) => positive_inputs_18_8_port, 
                           shift_out(7) => positive_inputs_18_7_port, 
                           shift_out(6) => positive_inputs_18_6_port, 
                           shift_out(5) => positive_inputs_18_5_port, 
                           shift_out(4) => positive_inputs_18_4_port, 
                           shift_out(3) => positive_inputs_18_3_port, 
                           shift_out(2) => positive_inputs_18_2_port, 
                           shift_out(1) => positive_inputs_18_1_port, 
                           shift_out(0) => n_1018);
   shifted_pos_19 : leftshifter_NbitShifter64_108 port map( shift_in(63) => 
                           positive_inputs_18_63_port, shift_in(62) => 
                           positive_inputs_18_62_port, shift_in(61) => 
                           positive_inputs_18_61_port, shift_in(60) => 
                           positive_inputs_18_60_port, shift_in(59) => 
                           positive_inputs_18_59_port, shift_in(58) => 
                           positive_inputs_18_58_port, shift_in(57) => 
                           positive_inputs_18_57_port, shift_in(56) => 
                           positive_inputs_18_56_port, shift_in(55) => 
                           positive_inputs_18_55_port, shift_in(54) => 
                           positive_inputs_18_54_port, shift_in(53) => 
                           positive_inputs_18_53_port, shift_in(52) => 
                           positive_inputs_18_52_port, shift_in(51) => 
                           positive_inputs_18_51_port, shift_in(50) => 
                           positive_inputs_18_50_port, shift_in(49) => 
                           positive_inputs_18_49_port, shift_in(48) => 
                           positive_inputs_18_48_port, shift_in(47) => 
                           positive_inputs_18_47_port, shift_in(46) => 
                           positive_inputs_18_46_port, shift_in(45) => 
                           positive_inputs_18_45_port, shift_in(44) => 
                           positive_inputs_18_44_port, shift_in(43) => 
                           positive_inputs_18_43_port, shift_in(42) => 
                           positive_inputs_18_42_port, shift_in(41) => 
                           positive_inputs_18_41_port, shift_in(40) => 
                           positive_inputs_18_40_port, shift_in(39) => 
                           positive_inputs_18_39_port, shift_in(38) => 
                           positive_inputs_18_38_port, shift_in(37) => 
                           positive_inputs_18_37_port, shift_in(36) => 
                           positive_inputs_18_36_port, shift_in(35) => 
                           positive_inputs_18_35_port, shift_in(34) => 
                           positive_inputs_18_34_port, shift_in(33) => 
                           positive_inputs_18_33_port, shift_in(32) => 
                           positive_inputs_18_32_port, shift_in(31) => 
                           positive_inputs_18_31_port, shift_in(30) => 
                           positive_inputs_18_30_port, shift_in(29) => 
                           positive_inputs_18_29_port, shift_in(28) => 
                           positive_inputs_18_28_port, shift_in(27) => 
                           positive_inputs_18_27_port, shift_in(26) => 
                           positive_inputs_18_26_port, shift_in(25) => 
                           positive_inputs_18_25_port, shift_in(24) => 
                           positive_inputs_18_24_port, shift_in(23) => 
                           positive_inputs_18_23_port, shift_in(22) => 
                           positive_inputs_18_22_port, shift_in(21) => 
                           positive_inputs_18_21_port, shift_in(20) => 
                           positive_inputs_18_20_port, shift_in(19) => 
                           positive_inputs_18_19_port, shift_in(18) => 
                           positive_inputs_18_18_port, shift_in(17) => 
                           positive_inputs_18_17_port, shift_in(16) => 
                           positive_inputs_18_16_port, shift_in(15) => 
                           positive_inputs_18_15_port, shift_in(14) => 
                           positive_inputs_18_14_port, shift_in(13) => 
                           positive_inputs_18_13_port, shift_in(12) => 
                           positive_inputs_18_12_port, shift_in(11) => 
                           positive_inputs_18_11_port, shift_in(10) => 
                           positive_inputs_18_10_port, shift_in(9) => 
                           positive_inputs_18_9_port, shift_in(8) => 
                           positive_inputs_18_8_port, shift_in(7) => 
                           positive_inputs_18_7_port, shift_in(6) => 
                           positive_inputs_18_6_port, shift_in(5) => 
                           positive_inputs_18_5_port, shift_in(4) => 
                           positive_inputs_18_4_port, shift_in(3) => 
                           positive_inputs_18_3_port, shift_in(2) => 
                           positive_inputs_18_2_port, shift_in(1) => 
                           positive_inputs_18_1_port, shift_in(0) => n8, 
                           shift_out(63) => positive_inputs_19_63_port, 
                           shift_out(62) => positive_inputs_19_62_port, 
                           shift_out(61) => positive_inputs_19_61_port, 
                           shift_out(60) => positive_inputs_19_60_port, 
                           shift_out(59) => positive_inputs_19_59_port, 
                           shift_out(58) => positive_inputs_19_58_port, 
                           shift_out(57) => positive_inputs_19_57_port, 
                           shift_out(56) => positive_inputs_19_56_port, 
                           shift_out(55) => positive_inputs_19_55_port, 
                           shift_out(54) => positive_inputs_19_54_port, 
                           shift_out(53) => positive_inputs_19_53_port, 
                           shift_out(52) => positive_inputs_19_52_port, 
                           shift_out(51) => positive_inputs_19_51_port, 
                           shift_out(50) => positive_inputs_19_50_port, 
                           shift_out(49) => positive_inputs_19_49_port, 
                           shift_out(48) => positive_inputs_19_48_port, 
                           shift_out(47) => positive_inputs_19_47_port, 
                           shift_out(46) => positive_inputs_19_46_port, 
                           shift_out(45) => positive_inputs_19_45_port, 
                           shift_out(44) => positive_inputs_19_44_port, 
                           shift_out(43) => positive_inputs_19_43_port, 
                           shift_out(42) => positive_inputs_19_42_port, 
                           shift_out(41) => positive_inputs_19_41_port, 
                           shift_out(40) => positive_inputs_19_40_port, 
                           shift_out(39) => positive_inputs_19_39_port, 
                           shift_out(38) => positive_inputs_19_38_port, 
                           shift_out(37) => positive_inputs_19_37_port, 
                           shift_out(36) => positive_inputs_19_36_port, 
                           shift_out(35) => positive_inputs_19_35_port, 
                           shift_out(34) => positive_inputs_19_34_port, 
                           shift_out(33) => positive_inputs_19_33_port, 
                           shift_out(32) => positive_inputs_19_32_port, 
                           shift_out(31) => positive_inputs_19_31_port, 
                           shift_out(30) => positive_inputs_19_30_port, 
                           shift_out(29) => positive_inputs_19_29_port, 
                           shift_out(28) => positive_inputs_19_28_port, 
                           shift_out(27) => positive_inputs_19_27_port, 
                           shift_out(26) => positive_inputs_19_26_port, 
                           shift_out(25) => positive_inputs_19_25_port, 
                           shift_out(24) => positive_inputs_19_24_port, 
                           shift_out(23) => positive_inputs_19_23_port, 
                           shift_out(22) => positive_inputs_19_22_port, 
                           shift_out(21) => positive_inputs_19_21_port, 
                           shift_out(20) => positive_inputs_19_20_port, 
                           shift_out(19) => positive_inputs_19_19_port, 
                           shift_out(18) => positive_inputs_19_18_port, 
                           shift_out(17) => positive_inputs_19_17_port, 
                           shift_out(16) => positive_inputs_19_16_port, 
                           shift_out(15) => positive_inputs_19_15_port, 
                           shift_out(14) => positive_inputs_19_14_port, 
                           shift_out(13) => positive_inputs_19_13_port, 
                           shift_out(12) => positive_inputs_19_12_port, 
                           shift_out(11) => positive_inputs_19_11_port, 
                           shift_out(10) => positive_inputs_19_10_port, 
                           shift_out(9) => positive_inputs_19_9_port, 
                           shift_out(8) => positive_inputs_19_8_port, 
                           shift_out(7) => positive_inputs_19_7_port, 
                           shift_out(6) => positive_inputs_19_6_port, 
                           shift_out(5) => positive_inputs_19_5_port, 
                           shift_out(4) => positive_inputs_19_4_port, 
                           shift_out(3) => positive_inputs_19_3_port, 
                           shift_out(2) => positive_inputs_19_2_port, 
                           shift_out(1) => positive_inputs_19_1_port, 
                           shift_out(0) => n_1019);
   shifted_pos_20 : leftshifter_NbitShifter64_107 port map( shift_in(63) => 
                           positive_inputs_19_63_port, shift_in(62) => 
                           positive_inputs_19_62_port, shift_in(61) => 
                           positive_inputs_19_61_port, shift_in(60) => 
                           positive_inputs_19_60_port, shift_in(59) => 
                           positive_inputs_19_59_port, shift_in(58) => 
                           positive_inputs_19_58_port, shift_in(57) => 
                           positive_inputs_19_57_port, shift_in(56) => 
                           positive_inputs_19_56_port, shift_in(55) => 
                           positive_inputs_19_55_port, shift_in(54) => 
                           positive_inputs_19_54_port, shift_in(53) => 
                           positive_inputs_19_53_port, shift_in(52) => 
                           positive_inputs_19_52_port, shift_in(51) => 
                           positive_inputs_19_51_port, shift_in(50) => 
                           positive_inputs_19_50_port, shift_in(49) => 
                           positive_inputs_19_49_port, shift_in(48) => 
                           positive_inputs_19_48_port, shift_in(47) => 
                           positive_inputs_19_47_port, shift_in(46) => 
                           positive_inputs_19_46_port, shift_in(45) => 
                           positive_inputs_19_45_port, shift_in(44) => 
                           positive_inputs_19_44_port, shift_in(43) => 
                           positive_inputs_19_43_port, shift_in(42) => 
                           positive_inputs_19_42_port, shift_in(41) => 
                           positive_inputs_19_41_port, shift_in(40) => 
                           positive_inputs_19_40_port, shift_in(39) => 
                           positive_inputs_19_39_port, shift_in(38) => 
                           positive_inputs_19_38_port, shift_in(37) => 
                           positive_inputs_19_37_port, shift_in(36) => 
                           positive_inputs_19_36_port, shift_in(35) => 
                           positive_inputs_19_35_port, shift_in(34) => 
                           positive_inputs_19_34_port, shift_in(33) => 
                           positive_inputs_19_33_port, shift_in(32) => 
                           positive_inputs_19_32_port, shift_in(31) => 
                           positive_inputs_19_31_port, shift_in(30) => 
                           positive_inputs_19_30_port, shift_in(29) => 
                           positive_inputs_19_29_port, shift_in(28) => 
                           positive_inputs_19_28_port, shift_in(27) => 
                           positive_inputs_19_27_port, shift_in(26) => 
                           positive_inputs_19_26_port, shift_in(25) => 
                           positive_inputs_19_25_port, shift_in(24) => 
                           positive_inputs_19_24_port, shift_in(23) => 
                           positive_inputs_19_23_port, shift_in(22) => 
                           positive_inputs_19_22_port, shift_in(21) => 
                           positive_inputs_19_21_port, shift_in(20) => 
                           positive_inputs_19_20_port, shift_in(19) => 
                           positive_inputs_19_19_port, shift_in(18) => 
                           positive_inputs_19_18_port, shift_in(17) => 
                           positive_inputs_19_17_port, shift_in(16) => 
                           positive_inputs_19_16_port, shift_in(15) => 
                           positive_inputs_19_15_port, shift_in(14) => 
                           positive_inputs_19_14_port, shift_in(13) => 
                           positive_inputs_19_13_port, shift_in(12) => 
                           positive_inputs_19_12_port, shift_in(11) => 
                           positive_inputs_19_11_port, shift_in(10) => 
                           positive_inputs_19_10_port, shift_in(9) => 
                           positive_inputs_19_9_port, shift_in(8) => 
                           positive_inputs_19_8_port, shift_in(7) => 
                           positive_inputs_19_7_port, shift_in(6) => 
                           positive_inputs_19_6_port, shift_in(5) => 
                           positive_inputs_19_5_port, shift_in(4) => 
                           positive_inputs_19_4_port, shift_in(3) => 
                           positive_inputs_19_3_port, shift_in(2) => 
                           positive_inputs_19_2_port, shift_in(1) => 
                           positive_inputs_19_1_port, shift_in(0) => n8, 
                           shift_out(63) => positive_inputs_20_63_port, 
                           shift_out(62) => positive_inputs_20_62_port, 
                           shift_out(61) => positive_inputs_20_61_port, 
                           shift_out(60) => positive_inputs_20_60_port, 
                           shift_out(59) => positive_inputs_20_59_port, 
                           shift_out(58) => positive_inputs_20_58_port, 
                           shift_out(57) => positive_inputs_20_57_port, 
                           shift_out(56) => positive_inputs_20_56_port, 
                           shift_out(55) => positive_inputs_20_55_port, 
                           shift_out(54) => positive_inputs_20_54_port, 
                           shift_out(53) => positive_inputs_20_53_port, 
                           shift_out(52) => positive_inputs_20_52_port, 
                           shift_out(51) => positive_inputs_20_51_port, 
                           shift_out(50) => positive_inputs_20_50_port, 
                           shift_out(49) => positive_inputs_20_49_port, 
                           shift_out(48) => positive_inputs_20_48_port, 
                           shift_out(47) => positive_inputs_20_47_port, 
                           shift_out(46) => positive_inputs_20_46_port, 
                           shift_out(45) => positive_inputs_20_45_port, 
                           shift_out(44) => positive_inputs_20_44_port, 
                           shift_out(43) => positive_inputs_20_43_port, 
                           shift_out(42) => positive_inputs_20_42_port, 
                           shift_out(41) => positive_inputs_20_41_port, 
                           shift_out(40) => positive_inputs_20_40_port, 
                           shift_out(39) => positive_inputs_20_39_port, 
                           shift_out(38) => positive_inputs_20_38_port, 
                           shift_out(37) => positive_inputs_20_37_port, 
                           shift_out(36) => positive_inputs_20_36_port, 
                           shift_out(35) => positive_inputs_20_35_port, 
                           shift_out(34) => positive_inputs_20_34_port, 
                           shift_out(33) => positive_inputs_20_33_port, 
                           shift_out(32) => positive_inputs_20_32_port, 
                           shift_out(31) => positive_inputs_20_31_port, 
                           shift_out(30) => positive_inputs_20_30_port, 
                           shift_out(29) => positive_inputs_20_29_port, 
                           shift_out(28) => positive_inputs_20_28_port, 
                           shift_out(27) => positive_inputs_20_27_port, 
                           shift_out(26) => positive_inputs_20_26_port, 
                           shift_out(25) => positive_inputs_20_25_port, 
                           shift_out(24) => positive_inputs_20_24_port, 
                           shift_out(23) => positive_inputs_20_23_port, 
                           shift_out(22) => positive_inputs_20_22_port, 
                           shift_out(21) => positive_inputs_20_21_port, 
                           shift_out(20) => positive_inputs_20_20_port, 
                           shift_out(19) => positive_inputs_20_19_port, 
                           shift_out(18) => positive_inputs_20_18_port, 
                           shift_out(17) => positive_inputs_20_17_port, 
                           shift_out(16) => positive_inputs_20_16_port, 
                           shift_out(15) => positive_inputs_20_15_port, 
                           shift_out(14) => positive_inputs_20_14_port, 
                           shift_out(13) => positive_inputs_20_13_port, 
                           shift_out(12) => positive_inputs_20_12_port, 
                           shift_out(11) => positive_inputs_20_11_port, 
                           shift_out(10) => positive_inputs_20_10_port, 
                           shift_out(9) => positive_inputs_20_9_port, 
                           shift_out(8) => positive_inputs_20_8_port, 
                           shift_out(7) => positive_inputs_20_7_port, 
                           shift_out(6) => positive_inputs_20_6_port, 
                           shift_out(5) => positive_inputs_20_5_port, 
                           shift_out(4) => positive_inputs_20_4_port, 
                           shift_out(3) => positive_inputs_20_3_port, 
                           shift_out(2) => positive_inputs_20_2_port, 
                           shift_out(1) => positive_inputs_20_1_port, 
                           shift_out(0) => n_1020);
   shifted_pos_21 : leftshifter_NbitShifter64_106 port map( shift_in(63) => 
                           positive_inputs_20_63_port, shift_in(62) => 
                           positive_inputs_20_62_port, shift_in(61) => 
                           positive_inputs_20_61_port, shift_in(60) => 
                           positive_inputs_20_60_port, shift_in(59) => 
                           positive_inputs_20_59_port, shift_in(58) => 
                           positive_inputs_20_58_port, shift_in(57) => 
                           positive_inputs_20_57_port, shift_in(56) => 
                           positive_inputs_20_56_port, shift_in(55) => 
                           positive_inputs_20_55_port, shift_in(54) => 
                           positive_inputs_20_54_port, shift_in(53) => 
                           positive_inputs_20_53_port, shift_in(52) => 
                           positive_inputs_20_52_port, shift_in(51) => 
                           positive_inputs_20_51_port, shift_in(50) => 
                           positive_inputs_20_50_port, shift_in(49) => 
                           positive_inputs_20_49_port, shift_in(48) => 
                           positive_inputs_20_48_port, shift_in(47) => 
                           positive_inputs_20_47_port, shift_in(46) => 
                           positive_inputs_20_46_port, shift_in(45) => 
                           positive_inputs_20_45_port, shift_in(44) => 
                           positive_inputs_20_44_port, shift_in(43) => 
                           positive_inputs_20_43_port, shift_in(42) => 
                           positive_inputs_20_42_port, shift_in(41) => 
                           positive_inputs_20_41_port, shift_in(40) => 
                           positive_inputs_20_40_port, shift_in(39) => 
                           positive_inputs_20_39_port, shift_in(38) => 
                           positive_inputs_20_38_port, shift_in(37) => 
                           positive_inputs_20_37_port, shift_in(36) => 
                           positive_inputs_20_36_port, shift_in(35) => 
                           positive_inputs_20_35_port, shift_in(34) => 
                           positive_inputs_20_34_port, shift_in(33) => 
                           positive_inputs_20_33_port, shift_in(32) => 
                           positive_inputs_20_32_port, shift_in(31) => 
                           positive_inputs_20_31_port, shift_in(30) => 
                           positive_inputs_20_30_port, shift_in(29) => 
                           positive_inputs_20_29_port, shift_in(28) => 
                           positive_inputs_20_28_port, shift_in(27) => 
                           positive_inputs_20_27_port, shift_in(26) => 
                           positive_inputs_20_26_port, shift_in(25) => 
                           positive_inputs_20_25_port, shift_in(24) => 
                           positive_inputs_20_24_port, shift_in(23) => 
                           positive_inputs_20_23_port, shift_in(22) => 
                           positive_inputs_20_22_port, shift_in(21) => 
                           positive_inputs_20_21_port, shift_in(20) => 
                           positive_inputs_20_20_port, shift_in(19) => 
                           positive_inputs_20_19_port, shift_in(18) => 
                           positive_inputs_20_18_port, shift_in(17) => 
                           positive_inputs_20_17_port, shift_in(16) => 
                           positive_inputs_20_16_port, shift_in(15) => 
                           positive_inputs_20_15_port, shift_in(14) => 
                           positive_inputs_20_14_port, shift_in(13) => 
                           positive_inputs_20_13_port, shift_in(12) => 
                           positive_inputs_20_12_port, shift_in(11) => 
                           positive_inputs_20_11_port, shift_in(10) => 
                           positive_inputs_20_10_port, shift_in(9) => 
                           positive_inputs_20_9_port, shift_in(8) => 
                           positive_inputs_20_8_port, shift_in(7) => 
                           positive_inputs_20_7_port, shift_in(6) => 
                           positive_inputs_20_6_port, shift_in(5) => 
                           positive_inputs_20_5_port, shift_in(4) => 
                           positive_inputs_20_4_port, shift_in(3) => 
                           positive_inputs_20_3_port, shift_in(2) => 
                           positive_inputs_20_2_port, shift_in(1) => 
                           positive_inputs_20_1_port, shift_in(0) => n8, 
                           shift_out(63) => positive_inputs_21_63_port, 
                           shift_out(62) => positive_inputs_21_62_port, 
                           shift_out(61) => positive_inputs_21_61_port, 
                           shift_out(60) => positive_inputs_21_60_port, 
                           shift_out(59) => positive_inputs_21_59_port, 
                           shift_out(58) => positive_inputs_21_58_port, 
                           shift_out(57) => positive_inputs_21_57_port, 
                           shift_out(56) => positive_inputs_21_56_port, 
                           shift_out(55) => positive_inputs_21_55_port, 
                           shift_out(54) => positive_inputs_21_54_port, 
                           shift_out(53) => positive_inputs_21_53_port, 
                           shift_out(52) => positive_inputs_21_52_port, 
                           shift_out(51) => positive_inputs_21_51_port, 
                           shift_out(50) => positive_inputs_21_50_port, 
                           shift_out(49) => positive_inputs_21_49_port, 
                           shift_out(48) => positive_inputs_21_48_port, 
                           shift_out(47) => positive_inputs_21_47_port, 
                           shift_out(46) => positive_inputs_21_46_port, 
                           shift_out(45) => positive_inputs_21_45_port, 
                           shift_out(44) => positive_inputs_21_44_port, 
                           shift_out(43) => positive_inputs_21_43_port, 
                           shift_out(42) => positive_inputs_21_42_port, 
                           shift_out(41) => positive_inputs_21_41_port, 
                           shift_out(40) => positive_inputs_21_40_port, 
                           shift_out(39) => positive_inputs_21_39_port, 
                           shift_out(38) => positive_inputs_21_38_port, 
                           shift_out(37) => positive_inputs_21_37_port, 
                           shift_out(36) => positive_inputs_21_36_port, 
                           shift_out(35) => positive_inputs_21_35_port, 
                           shift_out(34) => positive_inputs_21_34_port, 
                           shift_out(33) => positive_inputs_21_33_port, 
                           shift_out(32) => positive_inputs_21_32_port, 
                           shift_out(31) => positive_inputs_21_31_port, 
                           shift_out(30) => positive_inputs_21_30_port, 
                           shift_out(29) => positive_inputs_21_29_port, 
                           shift_out(28) => positive_inputs_21_28_port, 
                           shift_out(27) => positive_inputs_21_27_port, 
                           shift_out(26) => positive_inputs_21_26_port, 
                           shift_out(25) => positive_inputs_21_25_port, 
                           shift_out(24) => positive_inputs_21_24_port, 
                           shift_out(23) => positive_inputs_21_23_port, 
                           shift_out(22) => positive_inputs_21_22_port, 
                           shift_out(21) => positive_inputs_21_21_port, 
                           shift_out(20) => positive_inputs_21_20_port, 
                           shift_out(19) => positive_inputs_21_19_port, 
                           shift_out(18) => positive_inputs_21_18_port, 
                           shift_out(17) => positive_inputs_21_17_port, 
                           shift_out(16) => positive_inputs_21_16_port, 
                           shift_out(15) => positive_inputs_21_15_port, 
                           shift_out(14) => positive_inputs_21_14_port, 
                           shift_out(13) => positive_inputs_21_13_port, 
                           shift_out(12) => positive_inputs_21_12_port, 
                           shift_out(11) => positive_inputs_21_11_port, 
                           shift_out(10) => positive_inputs_21_10_port, 
                           shift_out(9) => positive_inputs_21_9_port, 
                           shift_out(8) => positive_inputs_21_8_port, 
                           shift_out(7) => positive_inputs_21_7_port, 
                           shift_out(6) => positive_inputs_21_6_port, 
                           shift_out(5) => positive_inputs_21_5_port, 
                           shift_out(4) => positive_inputs_21_4_port, 
                           shift_out(3) => positive_inputs_21_3_port, 
                           shift_out(2) => positive_inputs_21_2_port, 
                           shift_out(1) => positive_inputs_21_1_port, 
                           shift_out(0) => n_1021);
   shifted_pos_22 : leftshifter_NbitShifter64_105 port map( shift_in(63) => 
                           positive_inputs_21_63_port, shift_in(62) => 
                           positive_inputs_21_62_port, shift_in(61) => 
                           positive_inputs_21_61_port, shift_in(60) => 
                           positive_inputs_21_60_port, shift_in(59) => 
                           positive_inputs_21_59_port, shift_in(58) => 
                           positive_inputs_21_58_port, shift_in(57) => 
                           positive_inputs_21_57_port, shift_in(56) => 
                           positive_inputs_21_56_port, shift_in(55) => 
                           positive_inputs_21_55_port, shift_in(54) => 
                           positive_inputs_21_54_port, shift_in(53) => 
                           positive_inputs_21_53_port, shift_in(52) => 
                           positive_inputs_21_52_port, shift_in(51) => 
                           positive_inputs_21_51_port, shift_in(50) => 
                           positive_inputs_21_50_port, shift_in(49) => 
                           positive_inputs_21_49_port, shift_in(48) => 
                           positive_inputs_21_48_port, shift_in(47) => 
                           positive_inputs_21_47_port, shift_in(46) => 
                           positive_inputs_21_46_port, shift_in(45) => 
                           positive_inputs_21_45_port, shift_in(44) => 
                           positive_inputs_21_44_port, shift_in(43) => 
                           positive_inputs_21_43_port, shift_in(42) => 
                           positive_inputs_21_42_port, shift_in(41) => 
                           positive_inputs_21_41_port, shift_in(40) => 
                           positive_inputs_21_40_port, shift_in(39) => 
                           positive_inputs_21_39_port, shift_in(38) => 
                           positive_inputs_21_38_port, shift_in(37) => 
                           positive_inputs_21_37_port, shift_in(36) => 
                           positive_inputs_21_36_port, shift_in(35) => 
                           positive_inputs_21_35_port, shift_in(34) => 
                           positive_inputs_21_34_port, shift_in(33) => 
                           positive_inputs_21_33_port, shift_in(32) => 
                           positive_inputs_21_32_port, shift_in(31) => 
                           positive_inputs_21_31_port, shift_in(30) => 
                           positive_inputs_21_30_port, shift_in(29) => 
                           positive_inputs_21_29_port, shift_in(28) => 
                           positive_inputs_21_28_port, shift_in(27) => 
                           positive_inputs_21_27_port, shift_in(26) => 
                           positive_inputs_21_26_port, shift_in(25) => 
                           positive_inputs_21_25_port, shift_in(24) => 
                           positive_inputs_21_24_port, shift_in(23) => 
                           positive_inputs_21_23_port, shift_in(22) => 
                           positive_inputs_21_22_port, shift_in(21) => 
                           positive_inputs_21_21_port, shift_in(20) => 
                           positive_inputs_21_20_port, shift_in(19) => 
                           positive_inputs_21_19_port, shift_in(18) => 
                           positive_inputs_21_18_port, shift_in(17) => 
                           positive_inputs_21_17_port, shift_in(16) => 
                           positive_inputs_21_16_port, shift_in(15) => 
                           positive_inputs_21_15_port, shift_in(14) => 
                           positive_inputs_21_14_port, shift_in(13) => 
                           positive_inputs_21_13_port, shift_in(12) => 
                           positive_inputs_21_12_port, shift_in(11) => 
                           positive_inputs_21_11_port, shift_in(10) => 
                           positive_inputs_21_10_port, shift_in(9) => 
                           positive_inputs_21_9_port, shift_in(8) => 
                           positive_inputs_21_8_port, shift_in(7) => 
                           positive_inputs_21_7_port, shift_in(6) => 
                           positive_inputs_21_6_port, shift_in(5) => 
                           positive_inputs_21_5_port, shift_in(4) => 
                           positive_inputs_21_4_port, shift_in(3) => 
                           positive_inputs_21_3_port, shift_in(2) => 
                           positive_inputs_21_2_port, shift_in(1) => 
                           positive_inputs_21_1_port, shift_in(0) => n8, 
                           shift_out(63) => positive_inputs_22_63_port, 
                           shift_out(62) => positive_inputs_22_62_port, 
                           shift_out(61) => positive_inputs_22_61_port, 
                           shift_out(60) => positive_inputs_22_60_port, 
                           shift_out(59) => positive_inputs_22_59_port, 
                           shift_out(58) => positive_inputs_22_58_port, 
                           shift_out(57) => positive_inputs_22_57_port, 
                           shift_out(56) => positive_inputs_22_56_port, 
                           shift_out(55) => positive_inputs_22_55_port, 
                           shift_out(54) => positive_inputs_22_54_port, 
                           shift_out(53) => positive_inputs_22_53_port, 
                           shift_out(52) => positive_inputs_22_52_port, 
                           shift_out(51) => positive_inputs_22_51_port, 
                           shift_out(50) => positive_inputs_22_50_port, 
                           shift_out(49) => positive_inputs_22_49_port, 
                           shift_out(48) => positive_inputs_22_48_port, 
                           shift_out(47) => positive_inputs_22_47_port, 
                           shift_out(46) => positive_inputs_22_46_port, 
                           shift_out(45) => positive_inputs_22_45_port, 
                           shift_out(44) => positive_inputs_22_44_port, 
                           shift_out(43) => positive_inputs_22_43_port, 
                           shift_out(42) => positive_inputs_22_42_port, 
                           shift_out(41) => positive_inputs_22_41_port, 
                           shift_out(40) => positive_inputs_22_40_port, 
                           shift_out(39) => positive_inputs_22_39_port, 
                           shift_out(38) => positive_inputs_22_38_port, 
                           shift_out(37) => positive_inputs_22_37_port, 
                           shift_out(36) => positive_inputs_22_36_port, 
                           shift_out(35) => positive_inputs_22_35_port, 
                           shift_out(34) => positive_inputs_22_34_port, 
                           shift_out(33) => positive_inputs_22_33_port, 
                           shift_out(32) => positive_inputs_22_32_port, 
                           shift_out(31) => positive_inputs_22_31_port, 
                           shift_out(30) => positive_inputs_22_30_port, 
                           shift_out(29) => positive_inputs_22_29_port, 
                           shift_out(28) => positive_inputs_22_28_port, 
                           shift_out(27) => positive_inputs_22_27_port, 
                           shift_out(26) => positive_inputs_22_26_port, 
                           shift_out(25) => positive_inputs_22_25_port, 
                           shift_out(24) => positive_inputs_22_24_port, 
                           shift_out(23) => positive_inputs_22_23_port, 
                           shift_out(22) => positive_inputs_22_22_port, 
                           shift_out(21) => positive_inputs_22_21_port, 
                           shift_out(20) => positive_inputs_22_20_port, 
                           shift_out(19) => positive_inputs_22_19_port, 
                           shift_out(18) => positive_inputs_22_18_port, 
                           shift_out(17) => positive_inputs_22_17_port, 
                           shift_out(16) => positive_inputs_22_16_port, 
                           shift_out(15) => positive_inputs_22_15_port, 
                           shift_out(14) => positive_inputs_22_14_port, 
                           shift_out(13) => positive_inputs_22_13_port, 
                           shift_out(12) => positive_inputs_22_12_port, 
                           shift_out(11) => positive_inputs_22_11_port, 
                           shift_out(10) => positive_inputs_22_10_port, 
                           shift_out(9) => positive_inputs_22_9_port, 
                           shift_out(8) => positive_inputs_22_8_port, 
                           shift_out(7) => positive_inputs_22_7_port, 
                           shift_out(6) => positive_inputs_22_6_port, 
                           shift_out(5) => positive_inputs_22_5_port, 
                           shift_out(4) => positive_inputs_22_4_port, 
                           shift_out(3) => positive_inputs_22_3_port, 
                           shift_out(2) => positive_inputs_22_2_port, 
                           shift_out(1) => positive_inputs_22_1_port, 
                           shift_out(0) => n_1022);
   shifted_pos_23 : leftshifter_NbitShifter64_104 port map( shift_in(63) => 
                           positive_inputs_22_63_port, shift_in(62) => 
                           positive_inputs_22_62_port, shift_in(61) => 
                           positive_inputs_22_61_port, shift_in(60) => 
                           positive_inputs_22_60_port, shift_in(59) => 
                           positive_inputs_22_59_port, shift_in(58) => 
                           positive_inputs_22_58_port, shift_in(57) => 
                           positive_inputs_22_57_port, shift_in(56) => 
                           positive_inputs_22_56_port, shift_in(55) => 
                           positive_inputs_22_55_port, shift_in(54) => 
                           positive_inputs_22_54_port, shift_in(53) => 
                           positive_inputs_22_53_port, shift_in(52) => 
                           positive_inputs_22_52_port, shift_in(51) => 
                           positive_inputs_22_51_port, shift_in(50) => 
                           positive_inputs_22_50_port, shift_in(49) => 
                           positive_inputs_22_49_port, shift_in(48) => 
                           positive_inputs_22_48_port, shift_in(47) => 
                           positive_inputs_22_47_port, shift_in(46) => 
                           positive_inputs_22_46_port, shift_in(45) => 
                           positive_inputs_22_45_port, shift_in(44) => 
                           positive_inputs_22_44_port, shift_in(43) => 
                           positive_inputs_22_43_port, shift_in(42) => 
                           positive_inputs_22_42_port, shift_in(41) => 
                           positive_inputs_22_41_port, shift_in(40) => 
                           positive_inputs_22_40_port, shift_in(39) => 
                           positive_inputs_22_39_port, shift_in(38) => 
                           positive_inputs_22_38_port, shift_in(37) => 
                           positive_inputs_22_37_port, shift_in(36) => 
                           positive_inputs_22_36_port, shift_in(35) => 
                           positive_inputs_22_35_port, shift_in(34) => 
                           positive_inputs_22_34_port, shift_in(33) => 
                           positive_inputs_22_33_port, shift_in(32) => 
                           positive_inputs_22_32_port, shift_in(31) => 
                           positive_inputs_22_31_port, shift_in(30) => 
                           positive_inputs_22_30_port, shift_in(29) => 
                           positive_inputs_22_29_port, shift_in(28) => 
                           positive_inputs_22_28_port, shift_in(27) => 
                           positive_inputs_22_27_port, shift_in(26) => 
                           positive_inputs_22_26_port, shift_in(25) => 
                           positive_inputs_22_25_port, shift_in(24) => 
                           positive_inputs_22_24_port, shift_in(23) => 
                           positive_inputs_22_23_port, shift_in(22) => 
                           positive_inputs_22_22_port, shift_in(21) => 
                           positive_inputs_22_21_port, shift_in(20) => 
                           positive_inputs_22_20_port, shift_in(19) => 
                           positive_inputs_22_19_port, shift_in(18) => 
                           positive_inputs_22_18_port, shift_in(17) => 
                           positive_inputs_22_17_port, shift_in(16) => 
                           positive_inputs_22_16_port, shift_in(15) => 
                           positive_inputs_22_15_port, shift_in(14) => 
                           positive_inputs_22_14_port, shift_in(13) => 
                           positive_inputs_22_13_port, shift_in(12) => 
                           positive_inputs_22_12_port, shift_in(11) => 
                           positive_inputs_22_11_port, shift_in(10) => 
                           positive_inputs_22_10_port, shift_in(9) => 
                           positive_inputs_22_9_port, shift_in(8) => 
                           positive_inputs_22_8_port, shift_in(7) => 
                           positive_inputs_22_7_port, shift_in(6) => 
                           positive_inputs_22_6_port, shift_in(5) => 
                           positive_inputs_22_5_port, shift_in(4) => 
                           positive_inputs_22_4_port, shift_in(3) => 
                           positive_inputs_22_3_port, shift_in(2) => 
                           positive_inputs_22_2_port, shift_in(1) => 
                           positive_inputs_22_1_port, shift_in(0) => n8, 
                           shift_out(63) => positive_inputs_23_63_port, 
                           shift_out(62) => positive_inputs_23_62_port, 
                           shift_out(61) => positive_inputs_23_61_port, 
                           shift_out(60) => positive_inputs_23_60_port, 
                           shift_out(59) => positive_inputs_23_59_port, 
                           shift_out(58) => positive_inputs_23_58_port, 
                           shift_out(57) => positive_inputs_23_57_port, 
                           shift_out(56) => positive_inputs_23_56_port, 
                           shift_out(55) => positive_inputs_23_55_port, 
                           shift_out(54) => positive_inputs_23_54_port, 
                           shift_out(53) => positive_inputs_23_53_port, 
                           shift_out(52) => positive_inputs_23_52_port, 
                           shift_out(51) => positive_inputs_23_51_port, 
                           shift_out(50) => positive_inputs_23_50_port, 
                           shift_out(49) => positive_inputs_23_49_port, 
                           shift_out(48) => positive_inputs_23_48_port, 
                           shift_out(47) => positive_inputs_23_47_port, 
                           shift_out(46) => positive_inputs_23_46_port, 
                           shift_out(45) => positive_inputs_23_45_port, 
                           shift_out(44) => positive_inputs_23_44_port, 
                           shift_out(43) => positive_inputs_23_43_port, 
                           shift_out(42) => positive_inputs_23_42_port, 
                           shift_out(41) => positive_inputs_23_41_port, 
                           shift_out(40) => positive_inputs_23_40_port, 
                           shift_out(39) => positive_inputs_23_39_port, 
                           shift_out(38) => positive_inputs_23_38_port, 
                           shift_out(37) => positive_inputs_23_37_port, 
                           shift_out(36) => positive_inputs_23_36_port, 
                           shift_out(35) => positive_inputs_23_35_port, 
                           shift_out(34) => positive_inputs_23_34_port, 
                           shift_out(33) => positive_inputs_23_33_port, 
                           shift_out(32) => positive_inputs_23_32_port, 
                           shift_out(31) => positive_inputs_23_31_port, 
                           shift_out(30) => positive_inputs_23_30_port, 
                           shift_out(29) => positive_inputs_23_29_port, 
                           shift_out(28) => positive_inputs_23_28_port, 
                           shift_out(27) => positive_inputs_23_27_port, 
                           shift_out(26) => positive_inputs_23_26_port, 
                           shift_out(25) => positive_inputs_23_25_port, 
                           shift_out(24) => positive_inputs_23_24_port, 
                           shift_out(23) => positive_inputs_23_23_port, 
                           shift_out(22) => positive_inputs_23_22_port, 
                           shift_out(21) => positive_inputs_23_21_port, 
                           shift_out(20) => positive_inputs_23_20_port, 
                           shift_out(19) => positive_inputs_23_19_port, 
                           shift_out(18) => positive_inputs_23_18_port, 
                           shift_out(17) => positive_inputs_23_17_port, 
                           shift_out(16) => positive_inputs_23_16_port, 
                           shift_out(15) => positive_inputs_23_15_port, 
                           shift_out(14) => positive_inputs_23_14_port, 
                           shift_out(13) => positive_inputs_23_13_port, 
                           shift_out(12) => positive_inputs_23_12_port, 
                           shift_out(11) => positive_inputs_23_11_port, 
                           shift_out(10) => positive_inputs_23_10_port, 
                           shift_out(9) => positive_inputs_23_9_port, 
                           shift_out(8) => positive_inputs_23_8_port, 
                           shift_out(7) => positive_inputs_23_7_port, 
                           shift_out(6) => positive_inputs_23_6_port, 
                           shift_out(5) => positive_inputs_23_5_port, 
                           shift_out(4) => positive_inputs_23_4_port, 
                           shift_out(3) => positive_inputs_23_3_port, 
                           shift_out(2) => positive_inputs_23_2_port, 
                           shift_out(1) => positive_inputs_23_1_port, 
                           shift_out(0) => n_1023);
   shifted_pos_24 : leftshifter_NbitShifter64_103 port map( shift_in(63) => 
                           positive_inputs_23_63_port, shift_in(62) => 
                           positive_inputs_23_62_port, shift_in(61) => 
                           positive_inputs_23_61_port, shift_in(60) => 
                           positive_inputs_23_60_port, shift_in(59) => 
                           positive_inputs_23_59_port, shift_in(58) => 
                           positive_inputs_23_58_port, shift_in(57) => 
                           positive_inputs_23_57_port, shift_in(56) => 
                           positive_inputs_23_56_port, shift_in(55) => 
                           positive_inputs_23_55_port, shift_in(54) => 
                           positive_inputs_23_54_port, shift_in(53) => 
                           positive_inputs_23_53_port, shift_in(52) => 
                           positive_inputs_23_52_port, shift_in(51) => 
                           positive_inputs_23_51_port, shift_in(50) => 
                           positive_inputs_23_50_port, shift_in(49) => 
                           positive_inputs_23_49_port, shift_in(48) => 
                           positive_inputs_23_48_port, shift_in(47) => 
                           positive_inputs_23_47_port, shift_in(46) => 
                           positive_inputs_23_46_port, shift_in(45) => 
                           positive_inputs_23_45_port, shift_in(44) => 
                           positive_inputs_23_44_port, shift_in(43) => 
                           positive_inputs_23_43_port, shift_in(42) => 
                           positive_inputs_23_42_port, shift_in(41) => 
                           positive_inputs_23_41_port, shift_in(40) => 
                           positive_inputs_23_40_port, shift_in(39) => 
                           positive_inputs_23_39_port, shift_in(38) => 
                           positive_inputs_23_38_port, shift_in(37) => 
                           positive_inputs_23_37_port, shift_in(36) => 
                           positive_inputs_23_36_port, shift_in(35) => 
                           positive_inputs_23_35_port, shift_in(34) => 
                           positive_inputs_23_34_port, shift_in(33) => 
                           positive_inputs_23_33_port, shift_in(32) => 
                           positive_inputs_23_32_port, shift_in(31) => 
                           positive_inputs_23_31_port, shift_in(30) => 
                           positive_inputs_23_30_port, shift_in(29) => 
                           positive_inputs_23_29_port, shift_in(28) => 
                           positive_inputs_23_28_port, shift_in(27) => 
                           positive_inputs_23_27_port, shift_in(26) => 
                           positive_inputs_23_26_port, shift_in(25) => 
                           positive_inputs_23_25_port, shift_in(24) => 
                           positive_inputs_23_24_port, shift_in(23) => 
                           positive_inputs_23_23_port, shift_in(22) => 
                           positive_inputs_23_22_port, shift_in(21) => 
                           positive_inputs_23_21_port, shift_in(20) => 
                           positive_inputs_23_20_port, shift_in(19) => 
                           positive_inputs_23_19_port, shift_in(18) => 
                           positive_inputs_23_18_port, shift_in(17) => 
                           positive_inputs_23_17_port, shift_in(16) => 
                           positive_inputs_23_16_port, shift_in(15) => 
                           positive_inputs_23_15_port, shift_in(14) => 
                           positive_inputs_23_14_port, shift_in(13) => 
                           positive_inputs_23_13_port, shift_in(12) => 
                           positive_inputs_23_12_port, shift_in(11) => 
                           positive_inputs_23_11_port, shift_in(10) => 
                           positive_inputs_23_10_port, shift_in(9) => 
                           positive_inputs_23_9_port, shift_in(8) => 
                           positive_inputs_23_8_port, shift_in(7) => 
                           positive_inputs_23_7_port, shift_in(6) => 
                           positive_inputs_23_6_port, shift_in(5) => 
                           positive_inputs_23_5_port, shift_in(4) => 
                           positive_inputs_23_4_port, shift_in(3) => 
                           positive_inputs_23_3_port, shift_in(2) => 
                           positive_inputs_23_2_port, shift_in(1) => 
                           positive_inputs_23_1_port, shift_in(0) => n8, 
                           shift_out(63) => positive_inputs_24_63_port, 
                           shift_out(62) => positive_inputs_24_62_port, 
                           shift_out(61) => positive_inputs_24_61_port, 
                           shift_out(60) => positive_inputs_24_60_port, 
                           shift_out(59) => positive_inputs_24_59_port, 
                           shift_out(58) => positive_inputs_24_58_port, 
                           shift_out(57) => positive_inputs_24_57_port, 
                           shift_out(56) => positive_inputs_24_56_port, 
                           shift_out(55) => positive_inputs_24_55_port, 
                           shift_out(54) => positive_inputs_24_54_port, 
                           shift_out(53) => positive_inputs_24_53_port, 
                           shift_out(52) => positive_inputs_24_52_port, 
                           shift_out(51) => positive_inputs_24_51_port, 
                           shift_out(50) => positive_inputs_24_50_port, 
                           shift_out(49) => positive_inputs_24_49_port, 
                           shift_out(48) => positive_inputs_24_48_port, 
                           shift_out(47) => positive_inputs_24_47_port, 
                           shift_out(46) => positive_inputs_24_46_port, 
                           shift_out(45) => positive_inputs_24_45_port, 
                           shift_out(44) => positive_inputs_24_44_port, 
                           shift_out(43) => positive_inputs_24_43_port, 
                           shift_out(42) => positive_inputs_24_42_port, 
                           shift_out(41) => positive_inputs_24_41_port, 
                           shift_out(40) => positive_inputs_24_40_port, 
                           shift_out(39) => positive_inputs_24_39_port, 
                           shift_out(38) => positive_inputs_24_38_port, 
                           shift_out(37) => positive_inputs_24_37_port, 
                           shift_out(36) => positive_inputs_24_36_port, 
                           shift_out(35) => positive_inputs_24_35_port, 
                           shift_out(34) => positive_inputs_24_34_port, 
                           shift_out(33) => positive_inputs_24_33_port, 
                           shift_out(32) => positive_inputs_24_32_port, 
                           shift_out(31) => positive_inputs_24_31_port, 
                           shift_out(30) => positive_inputs_24_30_port, 
                           shift_out(29) => positive_inputs_24_29_port, 
                           shift_out(28) => positive_inputs_24_28_port, 
                           shift_out(27) => positive_inputs_24_27_port, 
                           shift_out(26) => positive_inputs_24_26_port, 
                           shift_out(25) => positive_inputs_24_25_port, 
                           shift_out(24) => positive_inputs_24_24_port, 
                           shift_out(23) => positive_inputs_24_23_port, 
                           shift_out(22) => positive_inputs_24_22_port, 
                           shift_out(21) => positive_inputs_24_21_port, 
                           shift_out(20) => positive_inputs_24_20_port, 
                           shift_out(19) => positive_inputs_24_19_port, 
                           shift_out(18) => positive_inputs_24_18_port, 
                           shift_out(17) => positive_inputs_24_17_port, 
                           shift_out(16) => positive_inputs_24_16_port, 
                           shift_out(15) => positive_inputs_24_15_port, 
                           shift_out(14) => positive_inputs_24_14_port, 
                           shift_out(13) => positive_inputs_24_13_port, 
                           shift_out(12) => positive_inputs_24_12_port, 
                           shift_out(11) => positive_inputs_24_11_port, 
                           shift_out(10) => positive_inputs_24_10_port, 
                           shift_out(9) => positive_inputs_24_9_port, 
                           shift_out(8) => positive_inputs_24_8_port, 
                           shift_out(7) => positive_inputs_24_7_port, 
                           shift_out(6) => positive_inputs_24_6_port, 
                           shift_out(5) => positive_inputs_24_5_port, 
                           shift_out(4) => positive_inputs_24_4_port, 
                           shift_out(3) => positive_inputs_24_3_port, 
                           shift_out(2) => positive_inputs_24_2_port, 
                           shift_out(1) => positive_inputs_24_1_port, 
                           shift_out(0) => n_1024);
   shifted_pos_25 : leftshifter_NbitShifter64_102 port map( shift_in(63) => 
                           positive_inputs_24_63_port, shift_in(62) => 
                           positive_inputs_24_62_port, shift_in(61) => 
                           positive_inputs_24_61_port, shift_in(60) => 
                           positive_inputs_24_60_port, shift_in(59) => 
                           positive_inputs_24_59_port, shift_in(58) => 
                           positive_inputs_24_58_port, shift_in(57) => 
                           positive_inputs_24_57_port, shift_in(56) => 
                           positive_inputs_24_56_port, shift_in(55) => 
                           positive_inputs_24_55_port, shift_in(54) => 
                           positive_inputs_24_54_port, shift_in(53) => 
                           positive_inputs_24_53_port, shift_in(52) => 
                           positive_inputs_24_52_port, shift_in(51) => 
                           positive_inputs_24_51_port, shift_in(50) => 
                           positive_inputs_24_50_port, shift_in(49) => 
                           positive_inputs_24_49_port, shift_in(48) => 
                           positive_inputs_24_48_port, shift_in(47) => 
                           positive_inputs_24_47_port, shift_in(46) => 
                           positive_inputs_24_46_port, shift_in(45) => 
                           positive_inputs_24_45_port, shift_in(44) => 
                           positive_inputs_24_44_port, shift_in(43) => 
                           positive_inputs_24_43_port, shift_in(42) => 
                           positive_inputs_24_42_port, shift_in(41) => 
                           positive_inputs_24_41_port, shift_in(40) => 
                           positive_inputs_24_40_port, shift_in(39) => 
                           positive_inputs_24_39_port, shift_in(38) => 
                           positive_inputs_24_38_port, shift_in(37) => 
                           positive_inputs_24_37_port, shift_in(36) => 
                           positive_inputs_24_36_port, shift_in(35) => 
                           positive_inputs_24_35_port, shift_in(34) => 
                           positive_inputs_24_34_port, shift_in(33) => 
                           positive_inputs_24_33_port, shift_in(32) => 
                           positive_inputs_24_32_port, shift_in(31) => 
                           positive_inputs_24_31_port, shift_in(30) => 
                           positive_inputs_24_30_port, shift_in(29) => 
                           positive_inputs_24_29_port, shift_in(28) => 
                           positive_inputs_24_28_port, shift_in(27) => 
                           positive_inputs_24_27_port, shift_in(26) => 
                           positive_inputs_24_26_port, shift_in(25) => 
                           positive_inputs_24_25_port, shift_in(24) => 
                           positive_inputs_24_24_port, shift_in(23) => 
                           positive_inputs_24_23_port, shift_in(22) => 
                           positive_inputs_24_22_port, shift_in(21) => 
                           positive_inputs_24_21_port, shift_in(20) => 
                           positive_inputs_24_20_port, shift_in(19) => 
                           positive_inputs_24_19_port, shift_in(18) => 
                           positive_inputs_24_18_port, shift_in(17) => 
                           positive_inputs_24_17_port, shift_in(16) => 
                           positive_inputs_24_16_port, shift_in(15) => 
                           positive_inputs_24_15_port, shift_in(14) => 
                           positive_inputs_24_14_port, shift_in(13) => 
                           positive_inputs_24_13_port, shift_in(12) => 
                           positive_inputs_24_12_port, shift_in(11) => 
                           positive_inputs_24_11_port, shift_in(10) => 
                           positive_inputs_24_10_port, shift_in(9) => 
                           positive_inputs_24_9_port, shift_in(8) => 
                           positive_inputs_24_8_port, shift_in(7) => 
                           positive_inputs_24_7_port, shift_in(6) => 
                           positive_inputs_24_6_port, shift_in(5) => 
                           positive_inputs_24_5_port, shift_in(4) => 
                           positive_inputs_24_4_port, shift_in(3) => 
                           positive_inputs_24_3_port, shift_in(2) => 
                           positive_inputs_24_2_port, shift_in(1) => 
                           positive_inputs_24_1_port, shift_in(0) => n8, 
                           shift_out(63) => positive_inputs_25_63_port, 
                           shift_out(62) => positive_inputs_25_62_port, 
                           shift_out(61) => positive_inputs_25_61_port, 
                           shift_out(60) => positive_inputs_25_60_port, 
                           shift_out(59) => positive_inputs_25_59_port, 
                           shift_out(58) => positive_inputs_25_58_port, 
                           shift_out(57) => positive_inputs_25_57_port, 
                           shift_out(56) => positive_inputs_25_56_port, 
                           shift_out(55) => positive_inputs_25_55_port, 
                           shift_out(54) => positive_inputs_25_54_port, 
                           shift_out(53) => positive_inputs_25_53_port, 
                           shift_out(52) => positive_inputs_25_52_port, 
                           shift_out(51) => positive_inputs_25_51_port, 
                           shift_out(50) => positive_inputs_25_50_port, 
                           shift_out(49) => positive_inputs_25_49_port, 
                           shift_out(48) => positive_inputs_25_48_port, 
                           shift_out(47) => positive_inputs_25_47_port, 
                           shift_out(46) => positive_inputs_25_46_port, 
                           shift_out(45) => positive_inputs_25_45_port, 
                           shift_out(44) => positive_inputs_25_44_port, 
                           shift_out(43) => positive_inputs_25_43_port, 
                           shift_out(42) => positive_inputs_25_42_port, 
                           shift_out(41) => positive_inputs_25_41_port, 
                           shift_out(40) => positive_inputs_25_40_port, 
                           shift_out(39) => positive_inputs_25_39_port, 
                           shift_out(38) => positive_inputs_25_38_port, 
                           shift_out(37) => positive_inputs_25_37_port, 
                           shift_out(36) => positive_inputs_25_36_port, 
                           shift_out(35) => positive_inputs_25_35_port, 
                           shift_out(34) => positive_inputs_25_34_port, 
                           shift_out(33) => positive_inputs_25_33_port, 
                           shift_out(32) => positive_inputs_25_32_port, 
                           shift_out(31) => positive_inputs_25_31_port, 
                           shift_out(30) => positive_inputs_25_30_port, 
                           shift_out(29) => positive_inputs_25_29_port, 
                           shift_out(28) => positive_inputs_25_28_port, 
                           shift_out(27) => positive_inputs_25_27_port, 
                           shift_out(26) => positive_inputs_25_26_port, 
                           shift_out(25) => positive_inputs_25_25_port, 
                           shift_out(24) => positive_inputs_25_24_port, 
                           shift_out(23) => positive_inputs_25_23_port, 
                           shift_out(22) => positive_inputs_25_22_port, 
                           shift_out(21) => positive_inputs_25_21_port, 
                           shift_out(20) => positive_inputs_25_20_port, 
                           shift_out(19) => positive_inputs_25_19_port, 
                           shift_out(18) => positive_inputs_25_18_port, 
                           shift_out(17) => positive_inputs_25_17_port, 
                           shift_out(16) => positive_inputs_25_16_port, 
                           shift_out(15) => positive_inputs_25_15_port, 
                           shift_out(14) => positive_inputs_25_14_port, 
                           shift_out(13) => positive_inputs_25_13_port, 
                           shift_out(12) => positive_inputs_25_12_port, 
                           shift_out(11) => positive_inputs_25_11_port, 
                           shift_out(10) => positive_inputs_25_10_port, 
                           shift_out(9) => positive_inputs_25_9_port, 
                           shift_out(8) => positive_inputs_25_8_port, 
                           shift_out(7) => positive_inputs_25_7_port, 
                           shift_out(6) => positive_inputs_25_6_port, 
                           shift_out(5) => positive_inputs_25_5_port, 
                           shift_out(4) => positive_inputs_25_4_port, 
                           shift_out(3) => positive_inputs_25_3_port, 
                           shift_out(2) => positive_inputs_25_2_port, 
                           shift_out(1) => positive_inputs_25_1_port, 
                           shift_out(0) => n_1025);
   shifted_pos_26 : leftshifter_NbitShifter64_101 port map( shift_in(63) => 
                           positive_inputs_25_63_port, shift_in(62) => 
                           positive_inputs_25_62_port, shift_in(61) => 
                           positive_inputs_25_61_port, shift_in(60) => 
                           positive_inputs_25_60_port, shift_in(59) => 
                           positive_inputs_25_59_port, shift_in(58) => 
                           positive_inputs_25_58_port, shift_in(57) => 
                           positive_inputs_25_57_port, shift_in(56) => 
                           positive_inputs_25_56_port, shift_in(55) => 
                           positive_inputs_25_55_port, shift_in(54) => 
                           positive_inputs_25_54_port, shift_in(53) => 
                           positive_inputs_25_53_port, shift_in(52) => 
                           positive_inputs_25_52_port, shift_in(51) => 
                           positive_inputs_25_51_port, shift_in(50) => 
                           positive_inputs_25_50_port, shift_in(49) => 
                           positive_inputs_25_49_port, shift_in(48) => 
                           positive_inputs_25_48_port, shift_in(47) => 
                           positive_inputs_25_47_port, shift_in(46) => 
                           positive_inputs_25_46_port, shift_in(45) => 
                           positive_inputs_25_45_port, shift_in(44) => 
                           positive_inputs_25_44_port, shift_in(43) => 
                           positive_inputs_25_43_port, shift_in(42) => 
                           positive_inputs_25_42_port, shift_in(41) => 
                           positive_inputs_25_41_port, shift_in(40) => 
                           positive_inputs_25_40_port, shift_in(39) => 
                           positive_inputs_25_39_port, shift_in(38) => 
                           positive_inputs_25_38_port, shift_in(37) => 
                           positive_inputs_25_37_port, shift_in(36) => 
                           positive_inputs_25_36_port, shift_in(35) => 
                           positive_inputs_25_35_port, shift_in(34) => 
                           positive_inputs_25_34_port, shift_in(33) => 
                           positive_inputs_25_33_port, shift_in(32) => 
                           positive_inputs_25_32_port, shift_in(31) => 
                           positive_inputs_25_31_port, shift_in(30) => 
                           positive_inputs_25_30_port, shift_in(29) => 
                           positive_inputs_25_29_port, shift_in(28) => 
                           positive_inputs_25_28_port, shift_in(27) => 
                           positive_inputs_25_27_port, shift_in(26) => 
                           positive_inputs_25_26_port, shift_in(25) => 
                           positive_inputs_25_25_port, shift_in(24) => 
                           positive_inputs_25_24_port, shift_in(23) => 
                           positive_inputs_25_23_port, shift_in(22) => 
                           positive_inputs_25_22_port, shift_in(21) => 
                           positive_inputs_25_21_port, shift_in(20) => 
                           positive_inputs_25_20_port, shift_in(19) => 
                           positive_inputs_25_19_port, shift_in(18) => 
                           positive_inputs_25_18_port, shift_in(17) => 
                           positive_inputs_25_17_port, shift_in(16) => 
                           positive_inputs_25_16_port, shift_in(15) => 
                           positive_inputs_25_15_port, shift_in(14) => 
                           positive_inputs_25_14_port, shift_in(13) => 
                           positive_inputs_25_13_port, shift_in(12) => 
                           positive_inputs_25_12_port, shift_in(11) => 
                           positive_inputs_25_11_port, shift_in(10) => 
                           positive_inputs_25_10_port, shift_in(9) => 
                           positive_inputs_25_9_port, shift_in(8) => 
                           positive_inputs_25_8_port, shift_in(7) => 
                           positive_inputs_25_7_port, shift_in(6) => 
                           positive_inputs_25_6_port, shift_in(5) => 
                           positive_inputs_25_5_port, shift_in(4) => 
                           positive_inputs_25_4_port, shift_in(3) => 
                           positive_inputs_25_3_port, shift_in(2) => 
                           positive_inputs_25_2_port, shift_in(1) => 
                           positive_inputs_25_1_port, shift_in(0) => n8, 
                           shift_out(63) => positive_inputs_26_63_port, 
                           shift_out(62) => positive_inputs_26_62_port, 
                           shift_out(61) => positive_inputs_26_61_port, 
                           shift_out(60) => positive_inputs_26_60_port, 
                           shift_out(59) => positive_inputs_26_59_port, 
                           shift_out(58) => positive_inputs_26_58_port, 
                           shift_out(57) => positive_inputs_26_57_port, 
                           shift_out(56) => positive_inputs_26_56_port, 
                           shift_out(55) => positive_inputs_26_55_port, 
                           shift_out(54) => positive_inputs_26_54_port, 
                           shift_out(53) => positive_inputs_26_53_port, 
                           shift_out(52) => positive_inputs_26_52_port, 
                           shift_out(51) => positive_inputs_26_51_port, 
                           shift_out(50) => positive_inputs_26_50_port, 
                           shift_out(49) => positive_inputs_26_49_port, 
                           shift_out(48) => positive_inputs_26_48_port, 
                           shift_out(47) => positive_inputs_26_47_port, 
                           shift_out(46) => positive_inputs_26_46_port, 
                           shift_out(45) => positive_inputs_26_45_port, 
                           shift_out(44) => positive_inputs_26_44_port, 
                           shift_out(43) => positive_inputs_26_43_port, 
                           shift_out(42) => positive_inputs_26_42_port, 
                           shift_out(41) => positive_inputs_26_41_port, 
                           shift_out(40) => positive_inputs_26_40_port, 
                           shift_out(39) => positive_inputs_26_39_port, 
                           shift_out(38) => positive_inputs_26_38_port, 
                           shift_out(37) => positive_inputs_26_37_port, 
                           shift_out(36) => positive_inputs_26_36_port, 
                           shift_out(35) => positive_inputs_26_35_port, 
                           shift_out(34) => positive_inputs_26_34_port, 
                           shift_out(33) => positive_inputs_26_33_port, 
                           shift_out(32) => positive_inputs_26_32_port, 
                           shift_out(31) => positive_inputs_26_31_port, 
                           shift_out(30) => positive_inputs_26_30_port, 
                           shift_out(29) => positive_inputs_26_29_port, 
                           shift_out(28) => positive_inputs_26_28_port, 
                           shift_out(27) => positive_inputs_26_27_port, 
                           shift_out(26) => positive_inputs_26_26_port, 
                           shift_out(25) => positive_inputs_26_25_port, 
                           shift_out(24) => positive_inputs_26_24_port, 
                           shift_out(23) => positive_inputs_26_23_port, 
                           shift_out(22) => positive_inputs_26_22_port, 
                           shift_out(21) => positive_inputs_26_21_port, 
                           shift_out(20) => positive_inputs_26_20_port, 
                           shift_out(19) => positive_inputs_26_19_port, 
                           shift_out(18) => positive_inputs_26_18_port, 
                           shift_out(17) => positive_inputs_26_17_port, 
                           shift_out(16) => positive_inputs_26_16_port, 
                           shift_out(15) => positive_inputs_26_15_port, 
                           shift_out(14) => positive_inputs_26_14_port, 
                           shift_out(13) => positive_inputs_26_13_port, 
                           shift_out(12) => positive_inputs_26_12_port, 
                           shift_out(11) => positive_inputs_26_11_port, 
                           shift_out(10) => positive_inputs_26_10_port, 
                           shift_out(9) => positive_inputs_26_9_port, 
                           shift_out(8) => positive_inputs_26_8_port, 
                           shift_out(7) => positive_inputs_26_7_port, 
                           shift_out(6) => positive_inputs_26_6_port, 
                           shift_out(5) => positive_inputs_26_5_port, 
                           shift_out(4) => positive_inputs_26_4_port, 
                           shift_out(3) => positive_inputs_26_3_port, 
                           shift_out(2) => positive_inputs_26_2_port, 
                           shift_out(1) => positive_inputs_26_1_port, 
                           shift_out(0) => n_1026);
   shifted_pos_27 : leftshifter_NbitShifter64_100 port map( shift_in(63) => 
                           positive_inputs_26_63_port, shift_in(62) => 
                           positive_inputs_26_62_port, shift_in(61) => 
                           positive_inputs_26_61_port, shift_in(60) => 
                           positive_inputs_26_60_port, shift_in(59) => 
                           positive_inputs_26_59_port, shift_in(58) => 
                           positive_inputs_26_58_port, shift_in(57) => 
                           positive_inputs_26_57_port, shift_in(56) => 
                           positive_inputs_26_56_port, shift_in(55) => 
                           positive_inputs_26_55_port, shift_in(54) => 
                           positive_inputs_26_54_port, shift_in(53) => 
                           positive_inputs_26_53_port, shift_in(52) => 
                           positive_inputs_26_52_port, shift_in(51) => 
                           positive_inputs_26_51_port, shift_in(50) => 
                           positive_inputs_26_50_port, shift_in(49) => 
                           positive_inputs_26_49_port, shift_in(48) => 
                           positive_inputs_26_48_port, shift_in(47) => 
                           positive_inputs_26_47_port, shift_in(46) => 
                           positive_inputs_26_46_port, shift_in(45) => 
                           positive_inputs_26_45_port, shift_in(44) => 
                           positive_inputs_26_44_port, shift_in(43) => 
                           positive_inputs_26_43_port, shift_in(42) => 
                           positive_inputs_26_42_port, shift_in(41) => 
                           positive_inputs_26_41_port, shift_in(40) => 
                           positive_inputs_26_40_port, shift_in(39) => 
                           positive_inputs_26_39_port, shift_in(38) => 
                           positive_inputs_26_38_port, shift_in(37) => 
                           positive_inputs_26_37_port, shift_in(36) => 
                           positive_inputs_26_36_port, shift_in(35) => 
                           positive_inputs_26_35_port, shift_in(34) => 
                           positive_inputs_26_34_port, shift_in(33) => 
                           positive_inputs_26_33_port, shift_in(32) => 
                           positive_inputs_26_32_port, shift_in(31) => 
                           positive_inputs_26_31_port, shift_in(30) => 
                           positive_inputs_26_30_port, shift_in(29) => 
                           positive_inputs_26_29_port, shift_in(28) => 
                           positive_inputs_26_28_port, shift_in(27) => 
                           positive_inputs_26_27_port, shift_in(26) => 
                           positive_inputs_26_26_port, shift_in(25) => 
                           positive_inputs_26_25_port, shift_in(24) => 
                           positive_inputs_26_24_port, shift_in(23) => 
                           positive_inputs_26_23_port, shift_in(22) => 
                           positive_inputs_26_22_port, shift_in(21) => 
                           positive_inputs_26_21_port, shift_in(20) => 
                           positive_inputs_26_20_port, shift_in(19) => 
                           positive_inputs_26_19_port, shift_in(18) => 
                           positive_inputs_26_18_port, shift_in(17) => 
                           positive_inputs_26_17_port, shift_in(16) => 
                           positive_inputs_26_16_port, shift_in(15) => 
                           positive_inputs_26_15_port, shift_in(14) => 
                           positive_inputs_26_14_port, shift_in(13) => 
                           positive_inputs_26_13_port, shift_in(12) => 
                           positive_inputs_26_12_port, shift_in(11) => 
                           positive_inputs_26_11_port, shift_in(10) => 
                           positive_inputs_26_10_port, shift_in(9) => 
                           positive_inputs_26_9_port, shift_in(8) => 
                           positive_inputs_26_8_port, shift_in(7) => 
                           positive_inputs_26_7_port, shift_in(6) => 
                           positive_inputs_26_6_port, shift_in(5) => 
                           positive_inputs_26_5_port, shift_in(4) => 
                           positive_inputs_26_4_port, shift_in(3) => 
                           positive_inputs_26_3_port, shift_in(2) => 
                           positive_inputs_26_2_port, shift_in(1) => 
                           positive_inputs_26_1_port, shift_in(0) => n8, 
                           shift_out(63) => positive_inputs_27_63_port, 
                           shift_out(62) => positive_inputs_27_62_port, 
                           shift_out(61) => positive_inputs_27_61_port, 
                           shift_out(60) => positive_inputs_27_60_port, 
                           shift_out(59) => positive_inputs_27_59_port, 
                           shift_out(58) => positive_inputs_27_58_port, 
                           shift_out(57) => positive_inputs_27_57_port, 
                           shift_out(56) => positive_inputs_27_56_port, 
                           shift_out(55) => positive_inputs_27_55_port, 
                           shift_out(54) => positive_inputs_27_54_port, 
                           shift_out(53) => positive_inputs_27_53_port, 
                           shift_out(52) => positive_inputs_27_52_port, 
                           shift_out(51) => positive_inputs_27_51_port, 
                           shift_out(50) => positive_inputs_27_50_port, 
                           shift_out(49) => positive_inputs_27_49_port, 
                           shift_out(48) => positive_inputs_27_48_port, 
                           shift_out(47) => positive_inputs_27_47_port, 
                           shift_out(46) => positive_inputs_27_46_port, 
                           shift_out(45) => positive_inputs_27_45_port, 
                           shift_out(44) => positive_inputs_27_44_port, 
                           shift_out(43) => positive_inputs_27_43_port, 
                           shift_out(42) => positive_inputs_27_42_port, 
                           shift_out(41) => positive_inputs_27_41_port, 
                           shift_out(40) => positive_inputs_27_40_port, 
                           shift_out(39) => positive_inputs_27_39_port, 
                           shift_out(38) => positive_inputs_27_38_port, 
                           shift_out(37) => positive_inputs_27_37_port, 
                           shift_out(36) => positive_inputs_27_36_port, 
                           shift_out(35) => positive_inputs_27_35_port, 
                           shift_out(34) => positive_inputs_27_34_port, 
                           shift_out(33) => positive_inputs_27_33_port, 
                           shift_out(32) => positive_inputs_27_32_port, 
                           shift_out(31) => positive_inputs_27_31_port, 
                           shift_out(30) => positive_inputs_27_30_port, 
                           shift_out(29) => positive_inputs_27_29_port, 
                           shift_out(28) => positive_inputs_27_28_port, 
                           shift_out(27) => positive_inputs_27_27_port, 
                           shift_out(26) => positive_inputs_27_26_port, 
                           shift_out(25) => positive_inputs_27_25_port, 
                           shift_out(24) => positive_inputs_27_24_port, 
                           shift_out(23) => positive_inputs_27_23_port, 
                           shift_out(22) => positive_inputs_27_22_port, 
                           shift_out(21) => positive_inputs_27_21_port, 
                           shift_out(20) => positive_inputs_27_20_port, 
                           shift_out(19) => positive_inputs_27_19_port, 
                           shift_out(18) => positive_inputs_27_18_port, 
                           shift_out(17) => positive_inputs_27_17_port, 
                           shift_out(16) => positive_inputs_27_16_port, 
                           shift_out(15) => positive_inputs_27_15_port, 
                           shift_out(14) => positive_inputs_27_14_port, 
                           shift_out(13) => positive_inputs_27_13_port, 
                           shift_out(12) => positive_inputs_27_12_port, 
                           shift_out(11) => positive_inputs_27_11_port, 
                           shift_out(10) => positive_inputs_27_10_port, 
                           shift_out(9) => positive_inputs_27_9_port, 
                           shift_out(8) => positive_inputs_27_8_port, 
                           shift_out(7) => positive_inputs_27_7_port, 
                           shift_out(6) => positive_inputs_27_6_port, 
                           shift_out(5) => positive_inputs_27_5_port, 
                           shift_out(4) => positive_inputs_27_4_port, 
                           shift_out(3) => positive_inputs_27_3_port, 
                           shift_out(2) => positive_inputs_27_2_port, 
                           shift_out(1) => positive_inputs_27_1_port, 
                           shift_out(0) => n_1027);
   shifted_pos_28 : leftshifter_NbitShifter64_99 port map( shift_in(63) => 
                           positive_inputs_27_63_port, shift_in(62) => 
                           positive_inputs_27_62_port, shift_in(61) => 
                           positive_inputs_27_61_port, shift_in(60) => 
                           positive_inputs_27_60_port, shift_in(59) => 
                           positive_inputs_27_59_port, shift_in(58) => 
                           positive_inputs_27_58_port, shift_in(57) => 
                           positive_inputs_27_57_port, shift_in(56) => 
                           positive_inputs_27_56_port, shift_in(55) => 
                           positive_inputs_27_55_port, shift_in(54) => 
                           positive_inputs_27_54_port, shift_in(53) => 
                           positive_inputs_27_53_port, shift_in(52) => 
                           positive_inputs_27_52_port, shift_in(51) => 
                           positive_inputs_27_51_port, shift_in(50) => 
                           positive_inputs_27_50_port, shift_in(49) => 
                           positive_inputs_27_49_port, shift_in(48) => 
                           positive_inputs_27_48_port, shift_in(47) => 
                           positive_inputs_27_47_port, shift_in(46) => 
                           positive_inputs_27_46_port, shift_in(45) => 
                           positive_inputs_27_45_port, shift_in(44) => 
                           positive_inputs_27_44_port, shift_in(43) => 
                           positive_inputs_27_43_port, shift_in(42) => 
                           positive_inputs_27_42_port, shift_in(41) => 
                           positive_inputs_27_41_port, shift_in(40) => 
                           positive_inputs_27_40_port, shift_in(39) => 
                           positive_inputs_27_39_port, shift_in(38) => 
                           positive_inputs_27_38_port, shift_in(37) => 
                           positive_inputs_27_37_port, shift_in(36) => 
                           positive_inputs_27_36_port, shift_in(35) => 
                           positive_inputs_27_35_port, shift_in(34) => 
                           positive_inputs_27_34_port, shift_in(33) => 
                           positive_inputs_27_33_port, shift_in(32) => 
                           positive_inputs_27_32_port, shift_in(31) => 
                           positive_inputs_27_31_port, shift_in(30) => 
                           positive_inputs_27_30_port, shift_in(29) => 
                           positive_inputs_27_29_port, shift_in(28) => 
                           positive_inputs_27_28_port, shift_in(27) => 
                           positive_inputs_27_27_port, shift_in(26) => 
                           positive_inputs_27_26_port, shift_in(25) => 
                           positive_inputs_27_25_port, shift_in(24) => 
                           positive_inputs_27_24_port, shift_in(23) => 
                           positive_inputs_27_23_port, shift_in(22) => 
                           positive_inputs_27_22_port, shift_in(21) => 
                           positive_inputs_27_21_port, shift_in(20) => 
                           positive_inputs_27_20_port, shift_in(19) => 
                           positive_inputs_27_19_port, shift_in(18) => 
                           positive_inputs_27_18_port, shift_in(17) => 
                           positive_inputs_27_17_port, shift_in(16) => 
                           positive_inputs_27_16_port, shift_in(15) => 
                           positive_inputs_27_15_port, shift_in(14) => 
                           positive_inputs_27_14_port, shift_in(13) => 
                           positive_inputs_27_13_port, shift_in(12) => 
                           positive_inputs_27_12_port, shift_in(11) => 
                           positive_inputs_27_11_port, shift_in(10) => 
                           positive_inputs_27_10_port, shift_in(9) => 
                           positive_inputs_27_9_port, shift_in(8) => 
                           positive_inputs_27_8_port, shift_in(7) => 
                           positive_inputs_27_7_port, shift_in(6) => 
                           positive_inputs_27_6_port, shift_in(5) => 
                           positive_inputs_27_5_port, shift_in(4) => 
                           positive_inputs_27_4_port, shift_in(3) => 
                           positive_inputs_27_3_port, shift_in(2) => 
                           positive_inputs_27_2_port, shift_in(1) => 
                           positive_inputs_27_1_port, shift_in(0) => n8, 
                           shift_out(63) => positive_inputs_28_63_port, 
                           shift_out(62) => positive_inputs_28_62_port, 
                           shift_out(61) => positive_inputs_28_61_port, 
                           shift_out(60) => positive_inputs_28_60_port, 
                           shift_out(59) => positive_inputs_28_59_port, 
                           shift_out(58) => positive_inputs_28_58_port, 
                           shift_out(57) => positive_inputs_28_57_port, 
                           shift_out(56) => positive_inputs_28_56_port, 
                           shift_out(55) => positive_inputs_28_55_port, 
                           shift_out(54) => positive_inputs_28_54_port, 
                           shift_out(53) => positive_inputs_28_53_port, 
                           shift_out(52) => positive_inputs_28_52_port, 
                           shift_out(51) => positive_inputs_28_51_port, 
                           shift_out(50) => positive_inputs_28_50_port, 
                           shift_out(49) => positive_inputs_28_49_port, 
                           shift_out(48) => positive_inputs_28_48_port, 
                           shift_out(47) => positive_inputs_28_47_port, 
                           shift_out(46) => positive_inputs_28_46_port, 
                           shift_out(45) => positive_inputs_28_45_port, 
                           shift_out(44) => positive_inputs_28_44_port, 
                           shift_out(43) => positive_inputs_28_43_port, 
                           shift_out(42) => positive_inputs_28_42_port, 
                           shift_out(41) => positive_inputs_28_41_port, 
                           shift_out(40) => positive_inputs_28_40_port, 
                           shift_out(39) => positive_inputs_28_39_port, 
                           shift_out(38) => positive_inputs_28_38_port, 
                           shift_out(37) => positive_inputs_28_37_port, 
                           shift_out(36) => positive_inputs_28_36_port, 
                           shift_out(35) => positive_inputs_28_35_port, 
                           shift_out(34) => positive_inputs_28_34_port, 
                           shift_out(33) => positive_inputs_28_33_port, 
                           shift_out(32) => positive_inputs_28_32_port, 
                           shift_out(31) => positive_inputs_28_31_port, 
                           shift_out(30) => positive_inputs_28_30_port, 
                           shift_out(29) => positive_inputs_28_29_port, 
                           shift_out(28) => positive_inputs_28_28_port, 
                           shift_out(27) => positive_inputs_28_27_port, 
                           shift_out(26) => positive_inputs_28_26_port, 
                           shift_out(25) => positive_inputs_28_25_port, 
                           shift_out(24) => positive_inputs_28_24_port, 
                           shift_out(23) => positive_inputs_28_23_port, 
                           shift_out(22) => positive_inputs_28_22_port, 
                           shift_out(21) => positive_inputs_28_21_port, 
                           shift_out(20) => positive_inputs_28_20_port, 
                           shift_out(19) => positive_inputs_28_19_port, 
                           shift_out(18) => positive_inputs_28_18_port, 
                           shift_out(17) => positive_inputs_28_17_port, 
                           shift_out(16) => positive_inputs_28_16_port, 
                           shift_out(15) => positive_inputs_28_15_port, 
                           shift_out(14) => positive_inputs_28_14_port, 
                           shift_out(13) => positive_inputs_28_13_port, 
                           shift_out(12) => positive_inputs_28_12_port, 
                           shift_out(11) => positive_inputs_28_11_port, 
                           shift_out(10) => positive_inputs_28_10_port, 
                           shift_out(9) => positive_inputs_28_9_port, 
                           shift_out(8) => positive_inputs_28_8_port, 
                           shift_out(7) => positive_inputs_28_7_port, 
                           shift_out(6) => positive_inputs_28_6_port, 
                           shift_out(5) => positive_inputs_28_5_port, 
                           shift_out(4) => positive_inputs_28_4_port, 
                           shift_out(3) => positive_inputs_28_3_port, 
                           shift_out(2) => positive_inputs_28_2_port, 
                           shift_out(1) => positive_inputs_28_1_port, 
                           shift_out(0) => n_1028);
   shifted_pos_29 : leftshifter_NbitShifter64_98 port map( shift_in(63) => 
                           positive_inputs_28_63_port, shift_in(62) => 
                           positive_inputs_28_62_port, shift_in(61) => 
                           positive_inputs_28_61_port, shift_in(60) => 
                           positive_inputs_28_60_port, shift_in(59) => 
                           positive_inputs_28_59_port, shift_in(58) => 
                           positive_inputs_28_58_port, shift_in(57) => 
                           positive_inputs_28_57_port, shift_in(56) => 
                           positive_inputs_28_56_port, shift_in(55) => 
                           positive_inputs_28_55_port, shift_in(54) => 
                           positive_inputs_28_54_port, shift_in(53) => 
                           positive_inputs_28_53_port, shift_in(52) => 
                           positive_inputs_28_52_port, shift_in(51) => 
                           positive_inputs_28_51_port, shift_in(50) => 
                           positive_inputs_28_50_port, shift_in(49) => 
                           positive_inputs_28_49_port, shift_in(48) => 
                           positive_inputs_28_48_port, shift_in(47) => 
                           positive_inputs_28_47_port, shift_in(46) => 
                           positive_inputs_28_46_port, shift_in(45) => 
                           positive_inputs_28_45_port, shift_in(44) => 
                           positive_inputs_28_44_port, shift_in(43) => 
                           positive_inputs_28_43_port, shift_in(42) => 
                           positive_inputs_28_42_port, shift_in(41) => 
                           positive_inputs_28_41_port, shift_in(40) => 
                           positive_inputs_28_40_port, shift_in(39) => 
                           positive_inputs_28_39_port, shift_in(38) => 
                           positive_inputs_28_38_port, shift_in(37) => 
                           positive_inputs_28_37_port, shift_in(36) => 
                           positive_inputs_28_36_port, shift_in(35) => 
                           positive_inputs_28_35_port, shift_in(34) => 
                           positive_inputs_28_34_port, shift_in(33) => 
                           positive_inputs_28_33_port, shift_in(32) => 
                           positive_inputs_28_32_port, shift_in(31) => 
                           positive_inputs_28_31_port, shift_in(30) => 
                           positive_inputs_28_30_port, shift_in(29) => 
                           positive_inputs_28_29_port, shift_in(28) => 
                           positive_inputs_28_28_port, shift_in(27) => 
                           positive_inputs_28_27_port, shift_in(26) => 
                           positive_inputs_28_26_port, shift_in(25) => 
                           positive_inputs_28_25_port, shift_in(24) => 
                           positive_inputs_28_24_port, shift_in(23) => 
                           positive_inputs_28_23_port, shift_in(22) => 
                           positive_inputs_28_22_port, shift_in(21) => 
                           positive_inputs_28_21_port, shift_in(20) => 
                           positive_inputs_28_20_port, shift_in(19) => 
                           positive_inputs_28_19_port, shift_in(18) => 
                           positive_inputs_28_18_port, shift_in(17) => 
                           positive_inputs_28_17_port, shift_in(16) => 
                           positive_inputs_28_16_port, shift_in(15) => 
                           positive_inputs_28_15_port, shift_in(14) => 
                           positive_inputs_28_14_port, shift_in(13) => 
                           positive_inputs_28_13_port, shift_in(12) => 
                           positive_inputs_28_12_port, shift_in(11) => 
                           positive_inputs_28_11_port, shift_in(10) => 
                           positive_inputs_28_10_port, shift_in(9) => 
                           positive_inputs_28_9_port, shift_in(8) => 
                           positive_inputs_28_8_port, shift_in(7) => 
                           positive_inputs_28_7_port, shift_in(6) => 
                           positive_inputs_28_6_port, shift_in(5) => 
                           positive_inputs_28_5_port, shift_in(4) => 
                           positive_inputs_28_4_port, shift_in(3) => 
                           positive_inputs_28_3_port, shift_in(2) => 
                           positive_inputs_28_2_port, shift_in(1) => 
                           positive_inputs_28_1_port, shift_in(0) => n8, 
                           shift_out(63) => positive_inputs_29_63_port, 
                           shift_out(62) => positive_inputs_29_62_port, 
                           shift_out(61) => positive_inputs_29_61_port, 
                           shift_out(60) => positive_inputs_29_60_port, 
                           shift_out(59) => positive_inputs_29_59_port, 
                           shift_out(58) => positive_inputs_29_58_port, 
                           shift_out(57) => positive_inputs_29_57_port, 
                           shift_out(56) => positive_inputs_29_56_port, 
                           shift_out(55) => positive_inputs_29_55_port, 
                           shift_out(54) => positive_inputs_29_54_port, 
                           shift_out(53) => positive_inputs_29_53_port, 
                           shift_out(52) => positive_inputs_29_52_port, 
                           shift_out(51) => positive_inputs_29_51_port, 
                           shift_out(50) => positive_inputs_29_50_port, 
                           shift_out(49) => positive_inputs_29_49_port, 
                           shift_out(48) => positive_inputs_29_48_port, 
                           shift_out(47) => positive_inputs_29_47_port, 
                           shift_out(46) => positive_inputs_29_46_port, 
                           shift_out(45) => positive_inputs_29_45_port, 
                           shift_out(44) => positive_inputs_29_44_port, 
                           shift_out(43) => positive_inputs_29_43_port, 
                           shift_out(42) => positive_inputs_29_42_port, 
                           shift_out(41) => positive_inputs_29_41_port, 
                           shift_out(40) => positive_inputs_29_40_port, 
                           shift_out(39) => positive_inputs_29_39_port, 
                           shift_out(38) => positive_inputs_29_38_port, 
                           shift_out(37) => positive_inputs_29_37_port, 
                           shift_out(36) => positive_inputs_29_36_port, 
                           shift_out(35) => positive_inputs_29_35_port, 
                           shift_out(34) => positive_inputs_29_34_port, 
                           shift_out(33) => positive_inputs_29_33_port, 
                           shift_out(32) => positive_inputs_29_32_port, 
                           shift_out(31) => positive_inputs_29_31_port, 
                           shift_out(30) => positive_inputs_29_30_port, 
                           shift_out(29) => positive_inputs_29_29_port, 
                           shift_out(28) => positive_inputs_29_28_port, 
                           shift_out(27) => positive_inputs_29_27_port, 
                           shift_out(26) => positive_inputs_29_26_port, 
                           shift_out(25) => positive_inputs_29_25_port, 
                           shift_out(24) => positive_inputs_29_24_port, 
                           shift_out(23) => positive_inputs_29_23_port, 
                           shift_out(22) => positive_inputs_29_22_port, 
                           shift_out(21) => positive_inputs_29_21_port, 
                           shift_out(20) => positive_inputs_29_20_port, 
                           shift_out(19) => positive_inputs_29_19_port, 
                           shift_out(18) => positive_inputs_29_18_port, 
                           shift_out(17) => positive_inputs_29_17_port, 
                           shift_out(16) => positive_inputs_29_16_port, 
                           shift_out(15) => positive_inputs_29_15_port, 
                           shift_out(14) => positive_inputs_29_14_port, 
                           shift_out(13) => positive_inputs_29_13_port, 
                           shift_out(12) => positive_inputs_29_12_port, 
                           shift_out(11) => positive_inputs_29_11_port, 
                           shift_out(10) => positive_inputs_29_10_port, 
                           shift_out(9) => positive_inputs_29_9_port, 
                           shift_out(8) => positive_inputs_29_8_port, 
                           shift_out(7) => positive_inputs_29_7_port, 
                           shift_out(6) => positive_inputs_29_6_port, 
                           shift_out(5) => positive_inputs_29_5_port, 
                           shift_out(4) => positive_inputs_29_4_port, 
                           shift_out(3) => positive_inputs_29_3_port, 
                           shift_out(2) => positive_inputs_29_2_port, 
                           shift_out(1) => positive_inputs_29_1_port, 
                           shift_out(0) => n_1029);
   shifted_pos_30 : leftshifter_NbitShifter64_97 port map( shift_in(63) => 
                           positive_inputs_29_63_port, shift_in(62) => 
                           positive_inputs_29_62_port, shift_in(61) => 
                           positive_inputs_29_61_port, shift_in(60) => 
                           positive_inputs_29_60_port, shift_in(59) => 
                           positive_inputs_29_59_port, shift_in(58) => 
                           positive_inputs_29_58_port, shift_in(57) => 
                           positive_inputs_29_57_port, shift_in(56) => 
                           positive_inputs_29_56_port, shift_in(55) => 
                           positive_inputs_29_55_port, shift_in(54) => 
                           positive_inputs_29_54_port, shift_in(53) => 
                           positive_inputs_29_53_port, shift_in(52) => 
                           positive_inputs_29_52_port, shift_in(51) => 
                           positive_inputs_29_51_port, shift_in(50) => 
                           positive_inputs_29_50_port, shift_in(49) => 
                           positive_inputs_29_49_port, shift_in(48) => 
                           positive_inputs_29_48_port, shift_in(47) => 
                           positive_inputs_29_47_port, shift_in(46) => 
                           positive_inputs_29_46_port, shift_in(45) => 
                           positive_inputs_29_45_port, shift_in(44) => 
                           positive_inputs_29_44_port, shift_in(43) => 
                           positive_inputs_29_43_port, shift_in(42) => 
                           positive_inputs_29_42_port, shift_in(41) => 
                           positive_inputs_29_41_port, shift_in(40) => 
                           positive_inputs_29_40_port, shift_in(39) => 
                           positive_inputs_29_39_port, shift_in(38) => 
                           positive_inputs_29_38_port, shift_in(37) => 
                           positive_inputs_29_37_port, shift_in(36) => 
                           positive_inputs_29_36_port, shift_in(35) => 
                           positive_inputs_29_35_port, shift_in(34) => 
                           positive_inputs_29_34_port, shift_in(33) => 
                           positive_inputs_29_33_port, shift_in(32) => 
                           positive_inputs_29_32_port, shift_in(31) => 
                           positive_inputs_29_31_port, shift_in(30) => 
                           positive_inputs_29_30_port, shift_in(29) => 
                           positive_inputs_29_29_port, shift_in(28) => 
                           positive_inputs_29_28_port, shift_in(27) => 
                           positive_inputs_29_27_port, shift_in(26) => 
                           positive_inputs_29_26_port, shift_in(25) => 
                           positive_inputs_29_25_port, shift_in(24) => 
                           positive_inputs_29_24_port, shift_in(23) => 
                           positive_inputs_29_23_port, shift_in(22) => 
                           positive_inputs_29_22_port, shift_in(21) => 
                           positive_inputs_29_21_port, shift_in(20) => 
                           positive_inputs_29_20_port, shift_in(19) => 
                           positive_inputs_29_19_port, shift_in(18) => 
                           positive_inputs_29_18_port, shift_in(17) => 
                           positive_inputs_29_17_port, shift_in(16) => 
                           positive_inputs_29_16_port, shift_in(15) => 
                           positive_inputs_29_15_port, shift_in(14) => 
                           positive_inputs_29_14_port, shift_in(13) => 
                           positive_inputs_29_13_port, shift_in(12) => 
                           positive_inputs_29_12_port, shift_in(11) => 
                           positive_inputs_29_11_port, shift_in(10) => 
                           positive_inputs_29_10_port, shift_in(9) => 
                           positive_inputs_29_9_port, shift_in(8) => 
                           positive_inputs_29_8_port, shift_in(7) => 
                           positive_inputs_29_7_port, shift_in(6) => 
                           positive_inputs_29_6_port, shift_in(5) => 
                           positive_inputs_29_5_port, shift_in(4) => 
                           positive_inputs_29_4_port, shift_in(3) => 
                           positive_inputs_29_3_port, shift_in(2) => 
                           positive_inputs_29_2_port, shift_in(1) => 
                           positive_inputs_29_1_port, shift_in(0) => n8, 
                           shift_out(63) => positive_inputs_30_63_port, 
                           shift_out(62) => positive_inputs_30_62_port, 
                           shift_out(61) => positive_inputs_30_61_port, 
                           shift_out(60) => positive_inputs_30_60_port, 
                           shift_out(59) => positive_inputs_30_59_port, 
                           shift_out(58) => positive_inputs_30_58_port, 
                           shift_out(57) => positive_inputs_30_57_port, 
                           shift_out(56) => positive_inputs_30_56_port, 
                           shift_out(55) => positive_inputs_30_55_port, 
                           shift_out(54) => positive_inputs_30_54_port, 
                           shift_out(53) => positive_inputs_30_53_port, 
                           shift_out(52) => positive_inputs_30_52_port, 
                           shift_out(51) => positive_inputs_30_51_port, 
                           shift_out(50) => positive_inputs_30_50_port, 
                           shift_out(49) => positive_inputs_30_49_port, 
                           shift_out(48) => positive_inputs_30_48_port, 
                           shift_out(47) => positive_inputs_30_47_port, 
                           shift_out(46) => positive_inputs_30_46_port, 
                           shift_out(45) => positive_inputs_30_45_port, 
                           shift_out(44) => positive_inputs_30_44_port, 
                           shift_out(43) => positive_inputs_30_43_port, 
                           shift_out(42) => positive_inputs_30_42_port, 
                           shift_out(41) => positive_inputs_30_41_port, 
                           shift_out(40) => positive_inputs_30_40_port, 
                           shift_out(39) => positive_inputs_30_39_port, 
                           shift_out(38) => positive_inputs_30_38_port, 
                           shift_out(37) => positive_inputs_30_37_port, 
                           shift_out(36) => positive_inputs_30_36_port, 
                           shift_out(35) => positive_inputs_30_35_port, 
                           shift_out(34) => positive_inputs_30_34_port, 
                           shift_out(33) => positive_inputs_30_33_port, 
                           shift_out(32) => positive_inputs_30_32_port, 
                           shift_out(31) => positive_inputs_30_31_port, 
                           shift_out(30) => positive_inputs_30_30_port, 
                           shift_out(29) => positive_inputs_30_29_port, 
                           shift_out(28) => positive_inputs_30_28_port, 
                           shift_out(27) => positive_inputs_30_27_port, 
                           shift_out(26) => positive_inputs_30_26_port, 
                           shift_out(25) => positive_inputs_30_25_port, 
                           shift_out(24) => positive_inputs_30_24_port, 
                           shift_out(23) => positive_inputs_30_23_port, 
                           shift_out(22) => positive_inputs_30_22_port, 
                           shift_out(21) => positive_inputs_30_21_port, 
                           shift_out(20) => positive_inputs_30_20_port, 
                           shift_out(19) => positive_inputs_30_19_port, 
                           shift_out(18) => positive_inputs_30_18_port, 
                           shift_out(17) => positive_inputs_30_17_port, 
                           shift_out(16) => positive_inputs_30_16_port, 
                           shift_out(15) => positive_inputs_30_15_port, 
                           shift_out(14) => positive_inputs_30_14_port, 
                           shift_out(13) => positive_inputs_30_13_port, 
                           shift_out(12) => positive_inputs_30_12_port, 
                           shift_out(11) => positive_inputs_30_11_port, 
                           shift_out(10) => positive_inputs_30_10_port, 
                           shift_out(9) => positive_inputs_30_9_port, 
                           shift_out(8) => positive_inputs_30_8_port, 
                           shift_out(7) => positive_inputs_30_7_port, 
                           shift_out(6) => positive_inputs_30_6_port, 
                           shift_out(5) => positive_inputs_30_5_port, 
                           shift_out(4) => positive_inputs_30_4_port, 
                           shift_out(3) => positive_inputs_30_3_port, 
                           shift_out(2) => positive_inputs_30_2_port, 
                           shift_out(1) => positive_inputs_30_1_port, 
                           shift_out(0) => n_1030);
   shifted_pos_31 : leftshifter_NbitShifter64_96 port map( shift_in(63) => 
                           positive_inputs_30_63_port, shift_in(62) => 
                           positive_inputs_30_62_port, shift_in(61) => 
                           positive_inputs_30_61_port, shift_in(60) => 
                           positive_inputs_30_60_port, shift_in(59) => 
                           positive_inputs_30_59_port, shift_in(58) => 
                           positive_inputs_30_58_port, shift_in(57) => 
                           positive_inputs_30_57_port, shift_in(56) => 
                           positive_inputs_30_56_port, shift_in(55) => 
                           positive_inputs_30_55_port, shift_in(54) => 
                           positive_inputs_30_54_port, shift_in(53) => 
                           positive_inputs_30_53_port, shift_in(52) => 
                           positive_inputs_30_52_port, shift_in(51) => 
                           positive_inputs_30_51_port, shift_in(50) => 
                           positive_inputs_30_50_port, shift_in(49) => 
                           positive_inputs_30_49_port, shift_in(48) => 
                           positive_inputs_30_48_port, shift_in(47) => 
                           positive_inputs_30_47_port, shift_in(46) => 
                           positive_inputs_30_46_port, shift_in(45) => 
                           positive_inputs_30_45_port, shift_in(44) => 
                           positive_inputs_30_44_port, shift_in(43) => 
                           positive_inputs_30_43_port, shift_in(42) => 
                           positive_inputs_30_42_port, shift_in(41) => 
                           positive_inputs_30_41_port, shift_in(40) => 
                           positive_inputs_30_40_port, shift_in(39) => 
                           positive_inputs_30_39_port, shift_in(38) => 
                           positive_inputs_30_38_port, shift_in(37) => 
                           positive_inputs_30_37_port, shift_in(36) => 
                           positive_inputs_30_36_port, shift_in(35) => 
                           positive_inputs_30_35_port, shift_in(34) => 
                           positive_inputs_30_34_port, shift_in(33) => 
                           positive_inputs_30_33_port, shift_in(32) => 
                           positive_inputs_30_32_port, shift_in(31) => 
                           positive_inputs_30_31_port, shift_in(30) => 
                           positive_inputs_30_30_port, shift_in(29) => 
                           positive_inputs_30_29_port, shift_in(28) => 
                           positive_inputs_30_28_port, shift_in(27) => 
                           positive_inputs_30_27_port, shift_in(26) => 
                           positive_inputs_30_26_port, shift_in(25) => 
                           positive_inputs_30_25_port, shift_in(24) => 
                           positive_inputs_30_24_port, shift_in(23) => 
                           positive_inputs_30_23_port, shift_in(22) => 
                           positive_inputs_30_22_port, shift_in(21) => 
                           positive_inputs_30_21_port, shift_in(20) => 
                           positive_inputs_30_20_port, shift_in(19) => 
                           positive_inputs_30_19_port, shift_in(18) => 
                           positive_inputs_30_18_port, shift_in(17) => 
                           positive_inputs_30_17_port, shift_in(16) => 
                           positive_inputs_30_16_port, shift_in(15) => 
                           positive_inputs_30_15_port, shift_in(14) => 
                           positive_inputs_30_14_port, shift_in(13) => 
                           positive_inputs_30_13_port, shift_in(12) => 
                           positive_inputs_30_12_port, shift_in(11) => 
                           positive_inputs_30_11_port, shift_in(10) => 
                           positive_inputs_30_10_port, shift_in(9) => 
                           positive_inputs_30_9_port, shift_in(8) => 
                           positive_inputs_30_8_port, shift_in(7) => 
                           positive_inputs_30_7_port, shift_in(6) => 
                           positive_inputs_30_6_port, shift_in(5) => 
                           positive_inputs_30_5_port, shift_in(4) => 
                           positive_inputs_30_4_port, shift_in(3) => 
                           positive_inputs_30_3_port, shift_in(2) => 
                           positive_inputs_30_2_port, shift_in(1) => 
                           positive_inputs_30_1_port, shift_in(0) => n8, 
                           shift_out(63) => positive_inputs_31_63_port, 
                           shift_out(62) => positive_inputs_31_62_port, 
                           shift_out(61) => positive_inputs_31_61_port, 
                           shift_out(60) => positive_inputs_31_60_port, 
                           shift_out(59) => positive_inputs_31_59_port, 
                           shift_out(58) => positive_inputs_31_58_port, 
                           shift_out(57) => positive_inputs_31_57_port, 
                           shift_out(56) => positive_inputs_31_56_port, 
                           shift_out(55) => positive_inputs_31_55_port, 
                           shift_out(54) => positive_inputs_31_54_port, 
                           shift_out(53) => positive_inputs_31_53_port, 
                           shift_out(52) => positive_inputs_31_52_port, 
                           shift_out(51) => positive_inputs_31_51_port, 
                           shift_out(50) => positive_inputs_31_50_port, 
                           shift_out(49) => positive_inputs_31_49_port, 
                           shift_out(48) => positive_inputs_31_48_port, 
                           shift_out(47) => positive_inputs_31_47_port, 
                           shift_out(46) => positive_inputs_31_46_port, 
                           shift_out(45) => positive_inputs_31_45_port, 
                           shift_out(44) => positive_inputs_31_44_port, 
                           shift_out(43) => positive_inputs_31_43_port, 
                           shift_out(42) => positive_inputs_31_42_port, 
                           shift_out(41) => positive_inputs_31_41_port, 
                           shift_out(40) => positive_inputs_31_40_port, 
                           shift_out(39) => positive_inputs_31_39_port, 
                           shift_out(38) => positive_inputs_31_38_port, 
                           shift_out(37) => positive_inputs_31_37_port, 
                           shift_out(36) => positive_inputs_31_36_port, 
                           shift_out(35) => positive_inputs_31_35_port, 
                           shift_out(34) => positive_inputs_31_34_port, 
                           shift_out(33) => positive_inputs_31_33_port, 
                           shift_out(32) => positive_inputs_31_32_port, 
                           shift_out(31) => positive_inputs_31_31_port, 
                           shift_out(30) => positive_inputs_31_30_port, 
                           shift_out(29) => positive_inputs_31_29_port, 
                           shift_out(28) => positive_inputs_31_28_port, 
                           shift_out(27) => positive_inputs_31_27_port, 
                           shift_out(26) => positive_inputs_31_26_port, 
                           shift_out(25) => positive_inputs_31_25_port, 
                           shift_out(24) => positive_inputs_31_24_port, 
                           shift_out(23) => positive_inputs_31_23_port, 
                           shift_out(22) => positive_inputs_31_22_port, 
                           shift_out(21) => positive_inputs_31_21_port, 
                           shift_out(20) => positive_inputs_31_20_port, 
                           shift_out(19) => positive_inputs_31_19_port, 
                           shift_out(18) => positive_inputs_31_18_port, 
                           shift_out(17) => positive_inputs_31_17_port, 
                           shift_out(16) => positive_inputs_31_16_port, 
                           shift_out(15) => positive_inputs_31_15_port, 
                           shift_out(14) => positive_inputs_31_14_port, 
                           shift_out(13) => positive_inputs_31_13_port, 
                           shift_out(12) => positive_inputs_31_12_port, 
                           shift_out(11) => positive_inputs_31_11_port, 
                           shift_out(10) => positive_inputs_31_10_port, 
                           shift_out(9) => positive_inputs_31_9_port, 
                           shift_out(8) => positive_inputs_31_8_port, 
                           shift_out(7) => positive_inputs_31_7_port, 
                           shift_out(6) => positive_inputs_31_6_port, 
                           shift_out(5) => positive_inputs_31_5_port, 
                           shift_out(4) => positive_inputs_31_4_port, 
                           shift_out(3) => positive_inputs_31_3_port, 
                           shift_out(2) => positive_inputs_31_2_port, 
                           shift_out(1) => positive_inputs_31_1_port, 
                           shift_out(0) => n_1031);
   shifted_pos_32 : leftshifter_NbitShifter64_95 port map( shift_in(63) => 
                           positive_inputs_31_63_port, shift_in(62) => 
                           positive_inputs_31_62_port, shift_in(61) => 
                           positive_inputs_31_61_port, shift_in(60) => 
                           positive_inputs_31_60_port, shift_in(59) => 
                           positive_inputs_31_59_port, shift_in(58) => 
                           positive_inputs_31_58_port, shift_in(57) => 
                           positive_inputs_31_57_port, shift_in(56) => 
                           positive_inputs_31_56_port, shift_in(55) => 
                           positive_inputs_31_55_port, shift_in(54) => 
                           positive_inputs_31_54_port, shift_in(53) => 
                           positive_inputs_31_53_port, shift_in(52) => 
                           positive_inputs_31_52_port, shift_in(51) => 
                           positive_inputs_31_51_port, shift_in(50) => 
                           positive_inputs_31_50_port, shift_in(49) => 
                           positive_inputs_31_49_port, shift_in(48) => 
                           positive_inputs_31_48_port, shift_in(47) => 
                           positive_inputs_31_47_port, shift_in(46) => 
                           positive_inputs_31_46_port, shift_in(45) => 
                           positive_inputs_31_45_port, shift_in(44) => 
                           positive_inputs_31_44_port, shift_in(43) => 
                           positive_inputs_31_43_port, shift_in(42) => 
                           positive_inputs_31_42_port, shift_in(41) => 
                           positive_inputs_31_41_port, shift_in(40) => 
                           positive_inputs_31_40_port, shift_in(39) => 
                           positive_inputs_31_39_port, shift_in(38) => 
                           positive_inputs_31_38_port, shift_in(37) => 
                           positive_inputs_31_37_port, shift_in(36) => 
                           positive_inputs_31_36_port, shift_in(35) => 
                           positive_inputs_31_35_port, shift_in(34) => 
                           positive_inputs_31_34_port, shift_in(33) => 
                           positive_inputs_31_33_port, shift_in(32) => 
                           positive_inputs_31_32_port, shift_in(31) => 
                           positive_inputs_31_31_port, shift_in(30) => 
                           positive_inputs_31_30_port, shift_in(29) => 
                           positive_inputs_31_29_port, shift_in(28) => 
                           positive_inputs_31_28_port, shift_in(27) => 
                           positive_inputs_31_27_port, shift_in(26) => 
                           positive_inputs_31_26_port, shift_in(25) => 
                           positive_inputs_31_25_port, shift_in(24) => 
                           positive_inputs_31_24_port, shift_in(23) => 
                           positive_inputs_31_23_port, shift_in(22) => 
                           positive_inputs_31_22_port, shift_in(21) => 
                           positive_inputs_31_21_port, shift_in(20) => 
                           positive_inputs_31_20_port, shift_in(19) => 
                           positive_inputs_31_19_port, shift_in(18) => 
                           positive_inputs_31_18_port, shift_in(17) => 
                           positive_inputs_31_17_port, shift_in(16) => 
                           positive_inputs_31_16_port, shift_in(15) => 
                           positive_inputs_31_15_port, shift_in(14) => 
                           positive_inputs_31_14_port, shift_in(13) => 
                           positive_inputs_31_13_port, shift_in(12) => 
                           positive_inputs_31_12_port, shift_in(11) => 
                           positive_inputs_31_11_port, shift_in(10) => 
                           positive_inputs_31_10_port, shift_in(9) => 
                           positive_inputs_31_9_port, shift_in(8) => 
                           positive_inputs_31_8_port, shift_in(7) => 
                           positive_inputs_31_7_port, shift_in(6) => 
                           positive_inputs_31_6_port, shift_in(5) => 
                           positive_inputs_31_5_port, shift_in(4) => 
                           positive_inputs_31_4_port, shift_in(3) => 
                           positive_inputs_31_3_port, shift_in(2) => 
                           positive_inputs_31_2_port, shift_in(1) => 
                           positive_inputs_31_1_port, shift_in(0) => n8, 
                           shift_out(63) => n_1032, shift_out(62) => n_1033, 
                           shift_out(61) => n_1034, shift_out(60) => n_1035, 
                           shift_out(59) => n_1036, shift_out(58) => n_1037, 
                           shift_out(57) => n_1038, shift_out(56) => n_1039, 
                           shift_out(55) => n_1040, shift_out(54) => n_1041, 
                           shift_out(53) => n_1042, shift_out(52) => n_1043, 
                           shift_out(51) => n_1044, shift_out(50) => n_1045, 
                           shift_out(49) => n_1046, shift_out(48) => n_1047, 
                           shift_out(47) => n_1048, shift_out(46) => n_1049, 
                           shift_out(45) => n_1050, shift_out(44) => n_1051, 
                           shift_out(43) => n_1052, shift_out(42) => n_1053, 
                           shift_out(41) => n_1054, shift_out(40) => n_1055, 
                           shift_out(39) => n_1056, shift_out(38) => n_1057, 
                           shift_out(37) => n_1058, shift_out(36) => n_1059, 
                           shift_out(35) => n_1060, shift_out(34) => n_1061, 
                           shift_out(33) => n_1062, shift_out(32) => n_1063, 
                           shift_out(31) => n_1064, shift_out(30) => n_1065, 
                           shift_out(29) => n_1066, shift_out(28) => n_1067, 
                           shift_out(27) => n_1068, shift_out(26) => n_1069, 
                           shift_out(25) => n_1070, shift_out(24) => n_1071, 
                           shift_out(23) => n_1072, shift_out(22) => n_1073, 
                           shift_out(21) => n_1074, shift_out(20) => n_1075, 
                           shift_out(19) => n_1076, shift_out(18) => n_1077, 
                           shift_out(17) => n_1078, shift_out(16) => n_1079, 
                           shift_out(15) => n_1080, shift_out(14) => n_1081, 
                           shift_out(13) => n_1082, shift_out(12) => n_1083, 
                           shift_out(11) => n_1084, shift_out(10) => n_1085, 
                           shift_out(9) => n_1086, shift_out(8) => n_1087, 
                           shift_out(7) => n_1088, shift_out(6) => n_1089, 
                           shift_out(5) => n_1090, shift_out(4) => n_1091, 
                           shift_out(3) => n_1092, shift_out(2) => n_1093, 
                           shift_out(1) => n_1094, shift_out(0) => n_1095);
   shifted_neg_1 : leftshifter_NbitShifter64_94 port map( shift_in(63) => 
                           negative_inputs_0_63_port, shift_in(62) => 
                           negative_inputs_0_62_port, shift_in(61) => 
                           negative_inputs_0_61_port, shift_in(60) => 
                           negative_inputs_0_60_port, shift_in(59) => 
                           negative_inputs_0_59_port, shift_in(58) => 
                           negative_inputs_0_58_port, shift_in(57) => 
                           negative_inputs_0_57_port, shift_in(56) => 
                           negative_inputs_0_56_port, shift_in(55) => 
                           negative_inputs_0_55_port, shift_in(54) => 
                           negative_inputs_0_54_port, shift_in(53) => 
                           negative_inputs_0_53_port, shift_in(52) => n40, 
                           shift_in(51) => n39, shift_in(50) => 
                           negative_inputs_0_50_port, shift_in(49) => n41, 
                           shift_in(48) => negative_inputs_0_48_port, 
                           shift_in(47) => negative_inputs_0_47_port, 
                           shift_in(46) => negative_inputs_0_46_port, 
                           shift_in(45) => negative_inputs_0_45_port, 
                           shift_in(44) => negative_inputs_0_44_port, 
                           shift_in(43) => negative_inputs_0_43_port, 
                           shift_in(42) => negative_inputs_0_42_port, 
                           shift_in(41) => negative_inputs_0_41_port, 
                           shift_in(40) => negative_inputs_0_40_port, 
                           shift_in(39) => negative_inputs_0_39_port, 
                           shift_in(38) => negative_inputs_0_38_port, 
                           shift_in(37) => negative_inputs_0_37_port, 
                           shift_in(36) => negative_inputs_0_36_port, 
                           shift_in(35) => negative_inputs_0_35_port, 
                           shift_in(34) => negative_inputs_0_34_port, 
                           shift_in(33) => negative_inputs_0_33_port, 
                           shift_in(32) => negative_inputs_0_32_port, 
                           shift_in(31) => negative_inputs_0_31_port, 
                           shift_in(30) => negative_inputs_0_30_port, 
                           shift_in(29) => negative_inputs_0_29_port, 
                           shift_in(28) => negative_inputs_0_28_port, 
                           shift_in(27) => negative_inputs_0_27_port, 
                           shift_in(26) => negative_inputs_0_26_port, 
                           shift_in(25) => negative_inputs_0_25_port, 
                           shift_in(24) => negative_inputs_0_24_port, 
                           shift_in(23) => negative_inputs_0_23_port, 
                           shift_in(22) => negative_inputs_0_22_port, 
                           shift_in(21) => negative_inputs_0_21_port, 
                           shift_in(20) => negative_inputs_0_20_port, 
                           shift_in(19) => negative_inputs_0_19_port, 
                           shift_in(18) => negative_inputs_0_18_port, 
                           shift_in(17) => n10, shift_in(16) => 
                           negative_inputs_0_16_port, shift_in(15) => 
                           negative_inputs_0_15_port, shift_in(14) => n9, 
                           shift_in(13) => negative_inputs_0_13_port, 
                           shift_in(12) => negative_inputs_0_12_port, 
                           shift_in(11) => negative_inputs_0_11_port, 
                           shift_in(10) => negative_inputs_0_10_port, 
                           shift_in(9) => negative_inputs_0_9_port, shift_in(8)
                           => negative_inputs_0_8_port, shift_in(7) => 
                           negative_inputs_0_7_port, shift_in(6) => 
                           negative_inputs_0_6_port, shift_in(5) => n11, 
                           shift_in(4) => n12, shift_in(3) => n14, shift_in(2) 
                           => negative_inputs_0_2_port, shift_in(1) => 
                           negative_inputs_0_1_port, shift_in(0) => 
                           negative_inputs_0_0_port, shift_out(63) => 
                           negative_inputs_1_63_port, shift_out(62) => 
                           negative_inputs_1_62_port, shift_out(61) => 
                           negative_inputs_1_61_port, shift_out(60) => 
                           negative_inputs_1_60_port, shift_out(59) => 
                           negative_inputs_1_59_port, shift_out(58) => 
                           negative_inputs_1_58_port, shift_out(57) => 
                           negative_inputs_1_57_port, shift_out(56) => 
                           negative_inputs_1_56_port, shift_out(55) => 
                           negative_inputs_1_55_port, shift_out(54) => 
                           negative_inputs_1_54_port, shift_out(53) => 
                           negative_inputs_1_53_port, shift_out(52) => 
                           negative_inputs_1_52_port, shift_out(51) => 
                           negative_inputs_1_51_port, shift_out(50) => 
                           negative_inputs_1_50_port, shift_out(49) => 
                           negative_inputs_1_49_port, shift_out(48) => 
                           negative_inputs_1_48_port, shift_out(47) => 
                           negative_inputs_1_47_port, shift_out(46) => 
                           negative_inputs_1_46_port, shift_out(45) => 
                           negative_inputs_1_45_port, shift_out(44) => 
                           negative_inputs_1_44_port, shift_out(43) => 
                           negative_inputs_1_43_port, shift_out(42) => 
                           negative_inputs_1_42_port, shift_out(41) => 
                           negative_inputs_1_41_port, shift_out(40) => 
                           negative_inputs_1_40_port, shift_out(39) => 
                           negative_inputs_1_39_port, shift_out(38) => 
                           negative_inputs_1_38_port, shift_out(37) => 
                           negative_inputs_1_37_port, shift_out(36) => 
                           negative_inputs_1_36_port, shift_out(35) => 
                           negative_inputs_1_35_port, shift_out(34) => 
                           negative_inputs_1_34_port, shift_out(33) => 
                           negative_inputs_1_33_port, shift_out(32) => 
                           negative_inputs_1_32_port, shift_out(31) => 
                           negative_inputs_1_31_port, shift_out(30) => 
                           negative_inputs_1_30_port, shift_out(29) => 
                           negative_inputs_1_29_port, shift_out(28) => 
                           negative_inputs_1_28_port, shift_out(27) => 
                           negative_inputs_1_27_port, shift_out(26) => 
                           negative_inputs_1_26_port, shift_out(25) => 
                           negative_inputs_1_25_port, shift_out(24) => 
                           negative_inputs_1_24_port, shift_out(23) => 
                           negative_inputs_1_23_port, shift_out(22) => 
                           negative_inputs_1_22_port, shift_out(21) => 
                           negative_inputs_1_21_port, shift_out(20) => 
                           negative_inputs_1_20_port, shift_out(19) => 
                           negative_inputs_1_19_port, shift_out(18) => 
                           negative_inputs_1_18_port, shift_out(17) => 
                           negative_inputs_1_17_port, shift_out(16) => 
                           negative_inputs_1_16_port, shift_out(15) => 
                           negative_inputs_1_15_port, shift_out(14) => 
                           negative_inputs_1_14_port, shift_out(13) => 
                           negative_inputs_1_13_port, shift_out(12) => 
                           negative_inputs_1_12_port, shift_out(11) => 
                           negative_inputs_1_11_port, shift_out(10) => 
                           negative_inputs_1_10_port, shift_out(9) => 
                           negative_inputs_1_9_port, shift_out(8) => 
                           negative_inputs_1_8_port, shift_out(7) => 
                           negative_inputs_1_7_port, shift_out(6) => 
                           negative_inputs_1_6_port, shift_out(5) => 
                           negative_inputs_1_5_port, shift_out(4) => 
                           negative_inputs_1_4_port, shift_out(3) => 
                           negative_inputs_1_3_port, shift_out(2) => 
                           negative_inputs_1_2_port, shift_out(1) => 
                           negative_inputs_1_1_port, shift_out(0) => n_1096);
   shifted_neg_2 : leftshifter_NbitShifter64_93 port map( shift_in(63) => 
                           negative_inputs_1_63_port, shift_in(62) => 
                           negative_inputs_1_62_port, shift_in(61) => 
                           negative_inputs_1_61_port, shift_in(60) => 
                           negative_inputs_1_60_port, shift_in(59) => 
                           negative_inputs_1_59_port, shift_in(58) => 
                           negative_inputs_1_58_port, shift_in(57) => 
                           negative_inputs_1_57_port, shift_in(56) => 
                           negative_inputs_1_56_port, shift_in(55) => 
                           negative_inputs_1_55_port, shift_in(54) => 
                           negative_inputs_1_54_port, shift_in(53) => 
                           negative_inputs_1_53_port, shift_in(52) => 
                           negative_inputs_1_52_port, shift_in(51) => 
                           negative_inputs_1_51_port, shift_in(50) => 
                           negative_inputs_1_50_port, shift_in(49) => 
                           negative_inputs_1_49_port, shift_in(48) => 
                           negative_inputs_1_48_port, shift_in(47) => 
                           negative_inputs_1_47_port, shift_in(46) => 
                           negative_inputs_1_46_port, shift_in(45) => 
                           negative_inputs_1_45_port, shift_in(44) => 
                           negative_inputs_1_44_port, shift_in(43) => 
                           negative_inputs_1_43_port, shift_in(42) => n17, 
                           shift_in(41) => negative_inputs_1_41_port, 
                           shift_in(40) => negative_inputs_1_40_port, 
                           shift_in(39) => negative_inputs_1_39_port, 
                           shift_in(38) => negative_inputs_1_38_port, 
                           shift_in(37) => n114, shift_in(36) => 
                           negative_inputs_1_36_port, shift_in(35) => 
                           negative_inputs_1_35_port, shift_in(34) => 
                           negative_inputs_1_34_port, shift_in(33) => 
                           negative_inputs_1_33_port, shift_in(32) => 
                           negative_inputs_1_32_port, shift_in(31) => 
                           negative_inputs_1_31_port, shift_in(30) => 
                           negative_inputs_1_30_port, shift_in(29) => 
                           negative_inputs_1_29_port, shift_in(28) => 
                           negative_inputs_1_28_port, shift_in(27) => 
                           negative_inputs_1_27_port, shift_in(26) => 
                           negative_inputs_1_26_port, shift_in(25) => 
                           negative_inputs_1_25_port, shift_in(24) => 
                           negative_inputs_1_24_port, shift_in(23) => 
                           negative_inputs_1_23_port, shift_in(22) => 
                           negative_inputs_1_22_port, shift_in(21) => 
                           negative_inputs_1_21_port, shift_in(20) => 
                           negative_inputs_1_20_port, shift_in(19) => 
                           negative_inputs_1_19_port, shift_in(18) => 
                           negative_inputs_1_18_port, shift_in(17) => 
                           negative_inputs_1_17_port, shift_in(16) => 
                           negative_inputs_1_16_port, shift_in(15) => 
                           negative_inputs_1_15_port, shift_in(14) => 
                           negative_inputs_1_14_port, shift_in(13) => 
                           negative_inputs_1_13_port, shift_in(12) => 
                           negative_inputs_1_12_port, shift_in(11) => 
                           negative_inputs_1_11_port, shift_in(10) => 
                           negative_inputs_1_10_port, shift_in(9) => 
                           negative_inputs_1_9_port, shift_in(8) => 
                           negative_inputs_1_8_port, shift_in(7) => 
                           negative_inputs_1_7_port, shift_in(6) => 
                           negative_inputs_1_6_port, shift_in(5) => 
                           negative_inputs_1_5_port, shift_in(4) => 
                           negative_inputs_1_4_port, shift_in(3) => n13, 
                           shift_in(2) => negative_inputs_1_2_port, shift_in(1)
                           => negative_inputs_1_1_port, shift_in(0) => n8, 
                           shift_out(63) => negative_inputs_2_63_port, 
                           shift_out(62) => negative_inputs_2_62_port, 
                           shift_out(61) => negative_inputs_2_61_port, 
                           shift_out(60) => negative_inputs_2_60_port, 
                           shift_out(59) => negative_inputs_2_59_port, 
                           shift_out(58) => negative_inputs_2_58_port, 
                           shift_out(57) => negative_inputs_2_57_port, 
                           shift_out(56) => negative_inputs_2_56_port, 
                           shift_out(55) => negative_inputs_2_55_port, 
                           shift_out(54) => negative_inputs_2_54_port, 
                           shift_out(53) => negative_inputs_2_53_port, 
                           shift_out(52) => negative_inputs_2_52_port, 
                           shift_out(51) => negative_inputs_2_51_port, 
                           shift_out(50) => negative_inputs_2_50_port, 
                           shift_out(49) => negative_inputs_2_49_port, 
                           shift_out(48) => negative_inputs_2_48_port, 
                           shift_out(47) => negative_inputs_2_47_port, 
                           shift_out(46) => negative_inputs_2_46_port, 
                           shift_out(45) => negative_inputs_2_45_port, 
                           shift_out(44) => negative_inputs_2_44_port, 
                           shift_out(43) => negative_inputs_2_43_port, 
                           shift_out(42) => negative_inputs_2_42_port, 
                           shift_out(41) => negative_inputs_2_41_port, 
                           shift_out(40) => negative_inputs_2_40_port, 
                           shift_out(39) => negative_inputs_2_39_port, 
                           shift_out(38) => negative_inputs_2_38_port, 
                           shift_out(37) => negative_inputs_2_37_port, 
                           shift_out(36) => negative_inputs_2_36_port, 
                           shift_out(35) => negative_inputs_2_35_port, 
                           shift_out(34) => negative_inputs_2_34_port, 
                           shift_out(33) => negative_inputs_2_33_port, 
                           shift_out(32) => negative_inputs_2_32_port, 
                           shift_out(31) => negative_inputs_2_31_port, 
                           shift_out(30) => negative_inputs_2_30_port, 
                           shift_out(29) => negative_inputs_2_29_port, 
                           shift_out(28) => negative_inputs_2_28_port, 
                           shift_out(27) => negative_inputs_2_27_port, 
                           shift_out(26) => negative_inputs_2_26_port, 
                           shift_out(25) => negative_inputs_2_25_port, 
                           shift_out(24) => negative_inputs_2_24_port, 
                           shift_out(23) => negative_inputs_2_23_port, 
                           shift_out(22) => negative_inputs_2_22_port, 
                           shift_out(21) => negative_inputs_2_21_port, 
                           shift_out(20) => negative_inputs_2_20_port, 
                           shift_out(19) => negative_inputs_2_19_port, 
                           shift_out(18) => negative_inputs_2_18_port, 
                           shift_out(17) => negative_inputs_2_17_port, 
                           shift_out(16) => negative_inputs_2_16_port, 
                           shift_out(15) => negative_inputs_2_15_port, 
                           shift_out(14) => negative_inputs_2_14_port, 
                           shift_out(13) => negative_inputs_2_13_port, 
                           shift_out(12) => negative_inputs_2_12_port, 
                           shift_out(11) => negative_inputs_2_11_port, 
                           shift_out(10) => negative_inputs_2_10_port, 
                           shift_out(9) => negative_inputs_2_9_port, 
                           shift_out(8) => negative_inputs_2_8_port, 
                           shift_out(7) => negative_inputs_2_7_port, 
                           shift_out(6) => negative_inputs_2_6_port, 
                           shift_out(5) => negative_inputs_2_5_port, 
                           shift_out(4) => negative_inputs_2_4_port, 
                           shift_out(3) => negative_inputs_2_3_port, 
                           shift_out(2) => negative_inputs_2_2_port, 
                           shift_out(1) => negative_inputs_2_1_port, 
                           shift_out(0) => n_1097);
   shifted_neg_3 : leftshifter_NbitShifter64_92 port map( shift_in(63) => 
                           negative_inputs_2_63_port, shift_in(62) => 
                           negative_inputs_2_62_port, shift_in(61) => 
                           negative_inputs_2_61_port, shift_in(60) => 
                           negative_inputs_2_60_port, shift_in(59) => 
                           negative_inputs_2_59_port, shift_in(58) => 
                           negative_inputs_2_58_port, shift_in(57) => 
                           negative_inputs_2_57_port, shift_in(56) => 
                           negative_inputs_2_56_port, shift_in(55) => 
                           negative_inputs_2_55_port, shift_in(54) => 
                           negative_inputs_2_54_port, shift_in(53) => 
                           negative_inputs_2_53_port, shift_in(52) => 
                           negative_inputs_2_52_port, shift_in(51) => 
                           negative_inputs_2_51_port, shift_in(50) => 
                           negative_inputs_2_50_port, shift_in(49) => 
                           negative_inputs_2_49_port, shift_in(48) => 
                           negative_inputs_2_48_port, shift_in(47) => 
                           negative_inputs_2_47_port, shift_in(46) => 
                           negative_inputs_2_46_port, shift_in(45) => 
                           negative_inputs_2_45_port, shift_in(44) => 
                           negative_inputs_2_44_port, shift_in(43) => 
                           negative_inputs_2_43_port, shift_in(42) => 
                           negative_inputs_2_42_port, shift_in(41) => 
                           negative_inputs_2_41_port, shift_in(40) => 
                           negative_inputs_2_40_port, shift_in(39) => 
                           negative_inputs_2_39_port, shift_in(38) => 
                           negative_inputs_2_38_port, shift_in(37) => n112, 
                           shift_in(36) => negative_inputs_2_36_port, 
                           shift_in(35) => negative_inputs_2_35_port, 
                           shift_in(34) => negative_inputs_2_34_port, 
                           shift_in(33) => negative_inputs_2_33_port, 
                           shift_in(32) => negative_inputs_2_32_port, 
                           shift_in(31) => negative_inputs_2_31_port, 
                           shift_in(30) => negative_inputs_2_30_port, 
                           shift_in(29) => negative_inputs_2_29_port, 
                           shift_in(28) => negative_inputs_2_28_port, 
                           shift_in(27) => negative_inputs_2_27_port, 
                           shift_in(26) => negative_inputs_2_26_port, 
                           shift_in(25) => negative_inputs_2_25_port, 
                           shift_in(24) => negative_inputs_2_24_port, 
                           shift_in(23) => negative_inputs_2_23_port, 
                           shift_in(22) => negative_inputs_2_22_port, 
                           shift_in(21) => negative_inputs_2_21_port, 
                           shift_in(20) => negative_inputs_2_20_port, 
                           shift_in(19) => negative_inputs_2_19_port, 
                           shift_in(18) => negative_inputs_2_18_port, 
                           shift_in(17) => negative_inputs_2_17_port, 
                           shift_in(16) => negative_inputs_2_16_port, 
                           shift_in(15) => negative_inputs_2_15_port, 
                           shift_in(14) => negative_inputs_2_14_port, 
                           shift_in(13) => negative_inputs_2_13_port, 
                           shift_in(12) => negative_inputs_2_12_port, 
                           shift_in(11) => negative_inputs_2_11_port, 
                           shift_in(10) => negative_inputs_2_10_port, 
                           shift_in(9) => negative_inputs_2_9_port, shift_in(8)
                           => negative_inputs_2_8_port, shift_in(7) => 
                           negative_inputs_2_7_port, shift_in(6) => 
                           negative_inputs_2_6_port, shift_in(5) => 
                           negative_inputs_2_5_port, shift_in(4) => 
                           negative_inputs_2_4_port, shift_in(3) => 
                           negative_inputs_2_3_port, shift_in(2) => 
                           negative_inputs_2_2_port, shift_in(1) => 
                           negative_inputs_2_1_port, shift_in(0) => n8, 
                           shift_out(63) => negative_inputs_3_63_port, 
                           shift_out(62) => negative_inputs_3_62_port, 
                           shift_out(61) => negative_inputs_3_61_port, 
                           shift_out(60) => negative_inputs_3_60_port, 
                           shift_out(59) => negative_inputs_3_59_port, 
                           shift_out(58) => negative_inputs_3_58_port, 
                           shift_out(57) => negative_inputs_3_57_port, 
                           shift_out(56) => negative_inputs_3_56_port, 
                           shift_out(55) => negative_inputs_3_55_port, 
                           shift_out(54) => negative_inputs_3_54_port, 
                           shift_out(53) => negative_inputs_3_53_port, 
                           shift_out(52) => negative_inputs_3_52_port, 
                           shift_out(51) => negative_inputs_3_51_port, 
                           shift_out(50) => negative_inputs_3_50_port, 
                           shift_out(49) => negative_inputs_3_49_port, 
                           shift_out(48) => negative_inputs_3_48_port, 
                           shift_out(47) => negative_inputs_3_47_port, 
                           shift_out(46) => negative_inputs_3_46_port, 
                           shift_out(45) => negative_inputs_3_45_port, 
                           shift_out(44) => negative_inputs_3_44_port, 
                           shift_out(43) => negative_inputs_3_43_port, 
                           shift_out(42) => negative_inputs_3_42_port, 
                           shift_out(41) => negative_inputs_3_41_port, 
                           shift_out(40) => negative_inputs_3_40_port, 
                           shift_out(39) => negative_inputs_3_39_port, 
                           shift_out(38) => negative_inputs_3_38_port, 
                           shift_out(37) => negative_inputs_3_37_port, 
                           shift_out(36) => negative_inputs_3_36_port, 
                           shift_out(35) => negative_inputs_3_35_port, 
                           shift_out(34) => negative_inputs_3_34_port, 
                           shift_out(33) => negative_inputs_3_33_port, 
                           shift_out(32) => negative_inputs_3_32_port, 
                           shift_out(31) => negative_inputs_3_31_port, 
                           shift_out(30) => negative_inputs_3_30_port, 
                           shift_out(29) => negative_inputs_3_29_port, 
                           shift_out(28) => negative_inputs_3_28_port, 
                           shift_out(27) => negative_inputs_3_27_port, 
                           shift_out(26) => negative_inputs_3_26_port, 
                           shift_out(25) => negative_inputs_3_25_port, 
                           shift_out(24) => negative_inputs_3_24_port, 
                           shift_out(23) => negative_inputs_3_23_port, 
                           shift_out(22) => negative_inputs_3_22_port, 
                           shift_out(21) => negative_inputs_3_21_port, 
                           shift_out(20) => negative_inputs_3_20_port, 
                           shift_out(19) => negative_inputs_3_19_port, 
                           shift_out(18) => negative_inputs_3_18_port, 
                           shift_out(17) => negative_inputs_3_17_port, 
                           shift_out(16) => negative_inputs_3_16_port, 
                           shift_out(15) => negative_inputs_3_15_port, 
                           shift_out(14) => negative_inputs_3_14_port, 
                           shift_out(13) => negative_inputs_3_13_port, 
                           shift_out(12) => negative_inputs_3_12_port, 
                           shift_out(11) => negative_inputs_3_11_port, 
                           shift_out(10) => negative_inputs_3_10_port, 
                           shift_out(9) => negative_inputs_3_9_port, 
                           shift_out(8) => negative_inputs_3_8_port, 
                           shift_out(7) => negative_inputs_3_7_port, 
                           shift_out(6) => negative_inputs_3_6_port, 
                           shift_out(5) => negative_inputs_3_5_port, 
                           shift_out(4) => negative_inputs_3_4_port, 
                           shift_out(3) => negative_inputs_3_3_port, 
                           shift_out(2) => negative_inputs_3_2_port, 
                           shift_out(1) => negative_inputs_3_1_port, 
                           shift_out(0) => n_1098);
   shifted_neg_4 : leftshifter_NbitShifter64_91 port map( shift_in(63) => 
                           negative_inputs_3_63_port, shift_in(62) => 
                           negative_inputs_3_62_port, shift_in(61) => 
                           negative_inputs_3_61_port, shift_in(60) => 
                           negative_inputs_3_60_port, shift_in(59) => 
                           negative_inputs_3_59_port, shift_in(58) => 
                           negative_inputs_3_58_port, shift_in(57) => 
                           negative_inputs_3_57_port, shift_in(56) => 
                           negative_inputs_3_56_port, shift_in(55) => 
                           negative_inputs_3_55_port, shift_in(54) => 
                           negative_inputs_3_54_port, shift_in(53) => 
                           negative_inputs_3_53_port, shift_in(52) => 
                           negative_inputs_3_52_port, shift_in(51) => 
                           negative_inputs_3_51_port, shift_in(50) => 
                           negative_inputs_3_50_port, shift_in(49) => 
                           negative_inputs_3_49_port, shift_in(48) => 
                           negative_inputs_3_48_port, shift_in(47) => 
                           negative_inputs_3_47_port, shift_in(46) => 
                           negative_inputs_3_46_port, shift_in(45) => 
                           negative_inputs_3_45_port, shift_in(44) => 
                           negative_inputs_3_44_port, shift_in(43) => 
                           negative_inputs_3_43_port, shift_in(42) => 
                           negative_inputs_3_42_port, shift_in(41) => 
                           negative_inputs_3_41_port, shift_in(40) => 
                           negative_inputs_3_40_port, shift_in(39) => 
                           negative_inputs_3_39_port, shift_in(38) => 
                           negative_inputs_3_38_port, shift_in(37) => n110, 
                           shift_in(36) => negative_inputs_3_36_port, 
                           shift_in(35) => negative_inputs_3_35_port, 
                           shift_in(34) => negative_inputs_3_34_port, 
                           shift_in(33) => negative_inputs_3_33_port, 
                           shift_in(32) => negative_inputs_3_32_port, 
                           shift_in(31) => negative_inputs_3_31_port, 
                           shift_in(30) => negative_inputs_3_30_port, 
                           shift_in(29) => negative_inputs_3_29_port, 
                           shift_in(28) => negative_inputs_3_28_port, 
                           shift_in(27) => negative_inputs_3_27_port, 
                           shift_in(26) => negative_inputs_3_26_port, 
                           shift_in(25) => negative_inputs_3_25_port, 
                           shift_in(24) => negative_inputs_3_24_port, 
                           shift_in(23) => negative_inputs_3_23_port, 
                           shift_in(22) => negative_inputs_3_22_port, 
                           shift_in(21) => negative_inputs_3_21_port, 
                           shift_in(20) => negative_inputs_3_20_port, 
                           shift_in(19) => negative_inputs_3_19_port, 
                           shift_in(18) => negative_inputs_3_18_port, 
                           shift_in(17) => negative_inputs_3_17_port, 
                           shift_in(16) => negative_inputs_3_16_port, 
                           shift_in(15) => negative_inputs_3_15_port, 
                           shift_in(14) => negative_inputs_3_14_port, 
                           shift_in(13) => negative_inputs_3_13_port, 
                           shift_in(12) => negative_inputs_3_12_port, 
                           shift_in(11) => negative_inputs_3_11_port, 
                           shift_in(10) => negative_inputs_3_10_port, 
                           shift_in(9) => negative_inputs_3_9_port, shift_in(8)
                           => negative_inputs_3_8_port, shift_in(7) => 
                           negative_inputs_3_7_port, shift_in(6) => 
                           negative_inputs_3_6_port, shift_in(5) => 
                           negative_inputs_3_5_port, shift_in(4) => 
                           negative_inputs_3_4_port, shift_in(3) => 
                           negative_inputs_3_3_port, shift_in(2) => 
                           negative_inputs_3_2_port, shift_in(1) => 
                           negative_inputs_3_1_port, shift_in(0) => n8, 
                           shift_out(63) => negative_inputs_4_63_port, 
                           shift_out(62) => negative_inputs_4_62_port, 
                           shift_out(61) => negative_inputs_4_61_port, 
                           shift_out(60) => negative_inputs_4_60_port, 
                           shift_out(59) => negative_inputs_4_59_port, 
                           shift_out(58) => negative_inputs_4_58_port, 
                           shift_out(57) => negative_inputs_4_57_port, 
                           shift_out(56) => negative_inputs_4_56_port, 
                           shift_out(55) => negative_inputs_4_55_port, 
                           shift_out(54) => negative_inputs_4_54_port, 
                           shift_out(53) => negative_inputs_4_53_port, 
                           shift_out(52) => negative_inputs_4_52_port, 
                           shift_out(51) => negative_inputs_4_51_port, 
                           shift_out(50) => negative_inputs_4_50_port, 
                           shift_out(49) => negative_inputs_4_49_port, 
                           shift_out(48) => negative_inputs_4_48_port, 
                           shift_out(47) => negative_inputs_4_47_port, 
                           shift_out(46) => negative_inputs_4_46_port, 
                           shift_out(45) => negative_inputs_4_45_port, 
                           shift_out(44) => negative_inputs_4_44_port, 
                           shift_out(43) => negative_inputs_4_43_port, 
                           shift_out(42) => negative_inputs_4_42_port, 
                           shift_out(41) => negative_inputs_4_41_port, 
                           shift_out(40) => negative_inputs_4_40_port, 
                           shift_out(39) => negative_inputs_4_39_port, 
                           shift_out(38) => negative_inputs_4_38_port, 
                           shift_out(37) => negative_inputs_4_37_port, 
                           shift_out(36) => negative_inputs_4_36_port, 
                           shift_out(35) => negative_inputs_4_35_port, 
                           shift_out(34) => negative_inputs_4_34_port, 
                           shift_out(33) => negative_inputs_4_33_port, 
                           shift_out(32) => negative_inputs_4_32_port, 
                           shift_out(31) => negative_inputs_4_31_port, 
                           shift_out(30) => negative_inputs_4_30_port, 
                           shift_out(29) => negative_inputs_4_29_port, 
                           shift_out(28) => negative_inputs_4_28_port, 
                           shift_out(27) => negative_inputs_4_27_port, 
                           shift_out(26) => negative_inputs_4_26_port, 
                           shift_out(25) => negative_inputs_4_25_port, 
                           shift_out(24) => negative_inputs_4_24_port, 
                           shift_out(23) => negative_inputs_4_23_port, 
                           shift_out(22) => negative_inputs_4_22_port, 
                           shift_out(21) => negative_inputs_4_21_port, 
                           shift_out(20) => negative_inputs_4_20_port, 
                           shift_out(19) => negative_inputs_4_19_port, 
                           shift_out(18) => negative_inputs_4_18_port, 
                           shift_out(17) => negative_inputs_4_17_port, 
                           shift_out(16) => negative_inputs_4_16_port, 
                           shift_out(15) => negative_inputs_4_15_port, 
                           shift_out(14) => negative_inputs_4_14_port, 
                           shift_out(13) => negative_inputs_4_13_port, 
                           shift_out(12) => negative_inputs_4_12_port, 
                           shift_out(11) => negative_inputs_4_11_port, 
                           shift_out(10) => negative_inputs_4_10_port, 
                           shift_out(9) => negative_inputs_4_9_port, 
                           shift_out(8) => negative_inputs_4_8_port, 
                           shift_out(7) => negative_inputs_4_7_port, 
                           shift_out(6) => negative_inputs_4_6_port, 
                           shift_out(5) => negative_inputs_4_5_port, 
                           shift_out(4) => negative_inputs_4_4_port, 
                           shift_out(3) => negative_inputs_4_3_port, 
                           shift_out(2) => negative_inputs_4_2_port, 
                           shift_out(1) => negative_inputs_4_1_port, 
                           shift_out(0) => n_1099);
   shifted_neg_5 : leftshifter_NbitShifter64_90 port map( shift_in(63) => 
                           negative_inputs_4_63_port, shift_in(62) => 
                           negative_inputs_4_62_port, shift_in(61) => 
                           negative_inputs_4_61_port, shift_in(60) => 
                           negative_inputs_4_60_port, shift_in(59) => 
                           negative_inputs_4_59_port, shift_in(58) => 
                           negative_inputs_4_58_port, shift_in(57) => 
                           negative_inputs_4_57_port, shift_in(56) => 
                           negative_inputs_4_56_port, shift_in(55) => 
                           negative_inputs_4_55_port, shift_in(54) => 
                           negative_inputs_4_54_port, shift_in(53) => 
                           negative_inputs_4_53_port, shift_in(52) => 
                           negative_inputs_4_52_port, shift_in(51) => 
                           negative_inputs_4_51_port, shift_in(50) => 
                           negative_inputs_4_50_port, shift_in(49) => 
                           negative_inputs_4_49_port, shift_in(48) => 
                           negative_inputs_4_48_port, shift_in(47) => 
                           negative_inputs_4_47_port, shift_in(46) => 
                           negative_inputs_4_46_port, shift_in(45) => 
                           negative_inputs_4_45_port, shift_in(44) => 
                           negative_inputs_4_44_port, shift_in(43) => 
                           negative_inputs_4_43_port, shift_in(42) => 
                           negative_inputs_4_42_port, shift_in(41) => 
                           negative_inputs_4_41_port, shift_in(40) => 
                           negative_inputs_4_40_port, shift_in(39) => 
                           negative_inputs_4_39_port, shift_in(38) => 
                           negative_inputs_4_38_port, shift_in(37) => n108, 
                           shift_in(36) => negative_inputs_4_36_port, 
                           shift_in(35) => negative_inputs_4_35_port, 
                           shift_in(34) => negative_inputs_4_34_port, 
                           shift_in(33) => negative_inputs_4_33_port, 
                           shift_in(32) => negative_inputs_4_32_port, 
                           shift_in(31) => negative_inputs_4_31_port, 
                           shift_in(30) => negative_inputs_4_30_port, 
                           shift_in(29) => negative_inputs_4_29_port, 
                           shift_in(28) => negative_inputs_4_28_port, 
                           shift_in(27) => negative_inputs_4_27_port, 
                           shift_in(26) => negative_inputs_4_26_port, 
                           shift_in(25) => negative_inputs_4_25_port, 
                           shift_in(24) => negative_inputs_4_24_port, 
                           shift_in(23) => negative_inputs_4_23_port, 
                           shift_in(22) => negative_inputs_4_22_port, 
                           shift_in(21) => negative_inputs_4_21_port, 
                           shift_in(20) => negative_inputs_4_20_port, 
                           shift_in(19) => negative_inputs_4_19_port, 
                           shift_in(18) => negative_inputs_4_18_port, 
                           shift_in(17) => negative_inputs_4_17_port, 
                           shift_in(16) => negative_inputs_4_16_port, 
                           shift_in(15) => negative_inputs_4_15_port, 
                           shift_in(14) => negative_inputs_4_14_port, 
                           shift_in(13) => negative_inputs_4_13_port, 
                           shift_in(12) => negative_inputs_4_12_port, 
                           shift_in(11) => negative_inputs_4_11_port, 
                           shift_in(10) => negative_inputs_4_10_port, 
                           shift_in(9) => negative_inputs_4_9_port, shift_in(8)
                           => negative_inputs_4_8_port, shift_in(7) => 
                           negative_inputs_4_7_port, shift_in(6) => 
                           negative_inputs_4_6_port, shift_in(5) => 
                           negative_inputs_4_5_port, shift_in(4) => 
                           negative_inputs_4_4_port, shift_in(3) => 
                           negative_inputs_4_3_port, shift_in(2) => 
                           negative_inputs_4_2_port, shift_in(1) => 
                           negative_inputs_4_1_port, shift_in(0) => n8, 
                           shift_out(63) => negative_inputs_5_63_port, 
                           shift_out(62) => negative_inputs_5_62_port, 
                           shift_out(61) => negative_inputs_5_61_port, 
                           shift_out(60) => negative_inputs_5_60_port, 
                           shift_out(59) => negative_inputs_5_59_port, 
                           shift_out(58) => negative_inputs_5_58_port, 
                           shift_out(57) => negative_inputs_5_57_port, 
                           shift_out(56) => negative_inputs_5_56_port, 
                           shift_out(55) => negative_inputs_5_55_port, 
                           shift_out(54) => negative_inputs_5_54_port, 
                           shift_out(53) => negative_inputs_5_53_port, 
                           shift_out(52) => negative_inputs_5_52_port, 
                           shift_out(51) => negative_inputs_5_51_port, 
                           shift_out(50) => negative_inputs_5_50_port, 
                           shift_out(49) => negative_inputs_5_49_port, 
                           shift_out(48) => negative_inputs_5_48_port, 
                           shift_out(47) => negative_inputs_5_47_port, 
                           shift_out(46) => negative_inputs_5_46_port, 
                           shift_out(45) => negative_inputs_5_45_port, 
                           shift_out(44) => negative_inputs_5_44_port, 
                           shift_out(43) => negative_inputs_5_43_port, 
                           shift_out(42) => negative_inputs_5_42_port, 
                           shift_out(41) => negative_inputs_5_41_port, 
                           shift_out(40) => negative_inputs_5_40_port, 
                           shift_out(39) => negative_inputs_5_39_port, 
                           shift_out(38) => negative_inputs_5_38_port, 
                           shift_out(37) => negative_inputs_5_37_port, 
                           shift_out(36) => negative_inputs_5_36_port, 
                           shift_out(35) => negative_inputs_5_35_port, 
                           shift_out(34) => negative_inputs_5_34_port, 
                           shift_out(33) => negative_inputs_5_33_port, 
                           shift_out(32) => negative_inputs_5_32_port, 
                           shift_out(31) => negative_inputs_5_31_port, 
                           shift_out(30) => negative_inputs_5_30_port, 
                           shift_out(29) => negative_inputs_5_29_port, 
                           shift_out(28) => negative_inputs_5_28_port, 
                           shift_out(27) => negative_inputs_5_27_port, 
                           shift_out(26) => negative_inputs_5_26_port, 
                           shift_out(25) => negative_inputs_5_25_port, 
                           shift_out(24) => negative_inputs_5_24_port, 
                           shift_out(23) => negative_inputs_5_23_port, 
                           shift_out(22) => negative_inputs_5_22_port, 
                           shift_out(21) => negative_inputs_5_21_port, 
                           shift_out(20) => negative_inputs_5_20_port, 
                           shift_out(19) => negative_inputs_5_19_port, 
                           shift_out(18) => negative_inputs_5_18_port, 
                           shift_out(17) => negative_inputs_5_17_port, 
                           shift_out(16) => negative_inputs_5_16_port, 
                           shift_out(15) => negative_inputs_5_15_port, 
                           shift_out(14) => negative_inputs_5_14_port, 
                           shift_out(13) => negative_inputs_5_13_port, 
                           shift_out(12) => negative_inputs_5_12_port, 
                           shift_out(11) => negative_inputs_5_11_port, 
                           shift_out(10) => negative_inputs_5_10_port, 
                           shift_out(9) => negative_inputs_5_9_port, 
                           shift_out(8) => negative_inputs_5_8_port, 
                           shift_out(7) => negative_inputs_5_7_port, 
                           shift_out(6) => negative_inputs_5_6_port, 
                           shift_out(5) => negative_inputs_5_5_port, 
                           shift_out(4) => negative_inputs_5_4_port, 
                           shift_out(3) => negative_inputs_5_3_port, 
                           shift_out(2) => negative_inputs_5_2_port, 
                           shift_out(1) => negative_inputs_5_1_port, 
                           shift_out(0) => n_1100);
   shifted_neg_6 : leftshifter_NbitShifter64_89 port map( shift_in(63) => 
                           negative_inputs_5_63_port, shift_in(62) => 
                           negative_inputs_5_62_port, shift_in(61) => 
                           negative_inputs_5_61_port, shift_in(60) => 
                           negative_inputs_5_60_port, shift_in(59) => 
                           negative_inputs_5_59_port, shift_in(58) => 
                           negative_inputs_5_58_port, shift_in(57) => 
                           negative_inputs_5_57_port, shift_in(56) => 
                           negative_inputs_5_56_port, shift_in(55) => 
                           negative_inputs_5_55_port, shift_in(54) => 
                           negative_inputs_5_54_port, shift_in(53) => 
                           negative_inputs_5_53_port, shift_in(52) => 
                           negative_inputs_5_52_port, shift_in(51) => 
                           negative_inputs_5_51_port, shift_in(50) => 
                           negative_inputs_5_50_port, shift_in(49) => 
                           negative_inputs_5_49_port, shift_in(48) => 
                           negative_inputs_5_48_port, shift_in(47) => 
                           negative_inputs_5_47_port, shift_in(46) => 
                           negative_inputs_5_46_port, shift_in(45) => 
                           negative_inputs_5_45_port, shift_in(44) => 
                           negative_inputs_5_44_port, shift_in(43) => 
                           negative_inputs_5_43_port, shift_in(42) => 
                           negative_inputs_5_42_port, shift_in(41) => 
                           negative_inputs_5_41_port, shift_in(40) => 
                           negative_inputs_5_40_port, shift_in(39) => 
                           negative_inputs_5_39_port, shift_in(38) => 
                           negative_inputs_5_38_port, shift_in(37) => n106, 
                           shift_in(36) => n104, shift_in(35) => n102, 
                           shift_in(34) => n100, shift_in(33) => n98, 
                           shift_in(32) => n96, shift_in(31) => n94, 
                           shift_in(30) => n92, shift_in(29) => n90, 
                           shift_in(28) => n88, shift_in(27) => n86, 
                           shift_in(26) => n84, shift_in(25) => n82, 
                           shift_in(24) => n80, shift_in(23) => n78, 
                           shift_in(22) => n76, shift_in(21) => n74, 
                           shift_in(20) => n72, shift_in(19) => n70, 
                           shift_in(18) => n68, shift_in(17) => n66, 
                           shift_in(16) => n64, shift_in(15) => n62, 
                           shift_in(14) => n60, shift_in(13) => n58, 
                           shift_in(12) => n56, shift_in(11) => n54, 
                           shift_in(10) => n52, shift_in(9) => n50, shift_in(8)
                           => n48, shift_in(7) => n46, shift_in(6) => n44, 
                           shift_in(5) => n42, shift_in(4) => 
                           negative_inputs_5_4_port, shift_in(3) => 
                           negative_inputs_5_3_port, shift_in(2) => 
                           negative_inputs_5_2_port, shift_in(1) => 
                           negative_inputs_5_1_port, shift_in(0) => n8, 
                           shift_out(63) => negative_inputs_6_63_port, 
                           shift_out(62) => negative_inputs_6_62_port, 
                           shift_out(61) => negative_inputs_6_61_port, 
                           shift_out(60) => negative_inputs_6_60_port, 
                           shift_out(59) => negative_inputs_6_59_port, 
                           shift_out(58) => negative_inputs_6_58_port, 
                           shift_out(57) => negative_inputs_6_57_port, 
                           shift_out(56) => negative_inputs_6_56_port, 
                           shift_out(55) => negative_inputs_6_55_port, 
                           shift_out(54) => negative_inputs_6_54_port, 
                           shift_out(53) => negative_inputs_6_53_port, 
                           shift_out(52) => negative_inputs_6_52_port, 
                           shift_out(51) => negative_inputs_6_51_port, 
                           shift_out(50) => negative_inputs_6_50_port, 
                           shift_out(49) => negative_inputs_6_49_port, 
                           shift_out(48) => negative_inputs_6_48_port, 
                           shift_out(47) => negative_inputs_6_47_port, 
                           shift_out(46) => negative_inputs_6_46_port, 
                           shift_out(45) => negative_inputs_6_45_port, 
                           shift_out(44) => negative_inputs_6_44_port, 
                           shift_out(43) => negative_inputs_6_43_port, 
                           shift_out(42) => negative_inputs_6_42_port, 
                           shift_out(41) => negative_inputs_6_41_port, 
                           shift_out(40) => negative_inputs_6_40_port, 
                           shift_out(39) => negative_inputs_6_39_port, 
                           shift_out(38) => negative_inputs_6_38_port, 
                           shift_out(37) => negative_inputs_6_37_port, 
                           shift_out(36) => negative_inputs_6_36_port, 
                           shift_out(35) => negative_inputs_6_35_port, 
                           shift_out(34) => negative_inputs_6_34_port, 
                           shift_out(33) => negative_inputs_6_33_port, 
                           shift_out(32) => negative_inputs_6_32_port, 
                           shift_out(31) => negative_inputs_6_31_port, 
                           shift_out(30) => negative_inputs_6_30_port, 
                           shift_out(29) => negative_inputs_6_29_port, 
                           shift_out(28) => negative_inputs_6_28_port, 
                           shift_out(27) => negative_inputs_6_27_port, 
                           shift_out(26) => negative_inputs_6_26_port, 
                           shift_out(25) => negative_inputs_6_25_port, 
                           shift_out(24) => negative_inputs_6_24_port, 
                           shift_out(23) => negative_inputs_6_23_port, 
                           shift_out(22) => negative_inputs_6_22_port, 
                           shift_out(21) => negative_inputs_6_21_port, 
                           shift_out(20) => negative_inputs_6_20_port, 
                           shift_out(19) => negative_inputs_6_19_port, 
                           shift_out(18) => negative_inputs_6_18_port, 
                           shift_out(17) => negative_inputs_6_17_port, 
                           shift_out(16) => negative_inputs_6_16_port, 
                           shift_out(15) => negative_inputs_6_15_port, 
                           shift_out(14) => negative_inputs_6_14_port, 
                           shift_out(13) => negative_inputs_6_13_port, 
                           shift_out(12) => negative_inputs_6_12_port, 
                           shift_out(11) => negative_inputs_6_11_port, 
                           shift_out(10) => negative_inputs_6_10_port, 
                           shift_out(9) => negative_inputs_6_9_port, 
                           shift_out(8) => negative_inputs_6_8_port, 
                           shift_out(7) => negative_inputs_6_7_port, 
                           shift_out(6) => negative_inputs_6_6_port, 
                           shift_out(5) => negative_inputs_6_5_port, 
                           shift_out(4) => negative_inputs_6_4_port, 
                           shift_out(3) => negative_inputs_6_3_port, 
                           shift_out(2) => negative_inputs_6_2_port, 
                           shift_out(1) => negative_inputs_6_1_port, 
                           shift_out(0) => n_1101);
   shifted_neg_7 : leftshifter_NbitShifter64_88 port map( shift_in(63) => 
                           negative_inputs_6_63_port, shift_in(62) => 
                           negative_inputs_6_62_port, shift_in(61) => 
                           negative_inputs_6_61_port, shift_in(60) => 
                           negative_inputs_6_60_port, shift_in(59) => 
                           negative_inputs_6_59_port, shift_in(58) => 
                           negative_inputs_6_58_port, shift_in(57) => 
                           negative_inputs_6_57_port, shift_in(56) => 
                           negative_inputs_6_56_port, shift_in(55) => 
                           negative_inputs_6_55_port, shift_in(54) => 
                           negative_inputs_6_54_port, shift_in(53) => 
                           negative_inputs_6_53_port, shift_in(52) => 
                           negative_inputs_6_52_port, shift_in(51) => 
                           negative_inputs_6_51_port, shift_in(50) => 
                           negative_inputs_6_50_port, shift_in(49) => 
                           negative_inputs_6_49_port, shift_in(48) => 
                           negative_inputs_6_48_port, shift_in(47) => 
                           negative_inputs_6_47_port, shift_in(46) => 
                           negative_inputs_6_46_port, shift_in(45) => 
                           negative_inputs_6_45_port, shift_in(44) => 
                           negative_inputs_6_44_port, shift_in(43) => 
                           negative_inputs_6_43_port, shift_in(42) => 
                           negative_inputs_6_42_port, shift_in(41) => 
                           negative_inputs_6_41_port, shift_in(40) => 
                           negative_inputs_6_40_port, shift_in(39) => 
                           negative_inputs_6_39_port, shift_in(38) => 
                           negative_inputs_6_38_port, shift_in(37) => 
                           negative_inputs_6_37_port, shift_in(36) => 
                           negative_inputs_6_36_port, shift_in(35) => 
                           negative_inputs_6_35_port, shift_in(34) => 
                           negative_inputs_6_34_port, shift_in(33) => 
                           negative_inputs_6_33_port, shift_in(32) => 
                           negative_inputs_6_32_port, shift_in(31) => 
                           negative_inputs_6_31_port, shift_in(30) => 
                           negative_inputs_6_30_port, shift_in(29) => 
                           negative_inputs_6_29_port, shift_in(28) => 
                           negative_inputs_6_28_port, shift_in(27) => 
                           negative_inputs_6_27_port, shift_in(26) => 
                           negative_inputs_6_26_port, shift_in(25) => 
                           negative_inputs_6_25_port, shift_in(24) => 
                           negative_inputs_6_24_port, shift_in(23) => 
                           negative_inputs_6_23_port, shift_in(22) => 
                           negative_inputs_6_22_port, shift_in(21) => 
                           negative_inputs_6_21_port, shift_in(20) => 
                           negative_inputs_6_20_port, shift_in(19) => 
                           negative_inputs_6_19_port, shift_in(18) => 
                           negative_inputs_6_18_port, shift_in(17) => 
                           negative_inputs_6_17_port, shift_in(16) => 
                           negative_inputs_6_16_port, shift_in(15) => 
                           negative_inputs_6_15_port, shift_in(14) => 
                           negative_inputs_6_14_port, shift_in(13) => 
                           negative_inputs_6_13_port, shift_in(12) => 
                           negative_inputs_6_12_port, shift_in(11) => 
                           negative_inputs_6_11_port, shift_in(10) => 
                           negative_inputs_6_10_port, shift_in(9) => 
                           negative_inputs_6_9_port, shift_in(8) => 
                           negative_inputs_6_8_port, shift_in(7) => 
                           negative_inputs_6_7_port, shift_in(6) => 
                           negative_inputs_6_6_port, shift_in(5) => 
                           negative_inputs_6_5_port, shift_in(4) => 
                           negative_inputs_6_4_port, shift_in(3) => 
                           negative_inputs_6_3_port, shift_in(2) => 
                           negative_inputs_6_2_port, shift_in(1) => 
                           negative_inputs_6_1_port, shift_in(0) => n8, 
                           shift_out(63) => negative_inputs_7_63_port, 
                           shift_out(62) => negative_inputs_7_62_port, 
                           shift_out(61) => negative_inputs_7_61_port, 
                           shift_out(60) => negative_inputs_7_60_port, 
                           shift_out(59) => negative_inputs_7_59_port, 
                           shift_out(58) => negative_inputs_7_58_port, 
                           shift_out(57) => negative_inputs_7_57_port, 
                           shift_out(56) => negative_inputs_7_56_port, 
                           shift_out(55) => negative_inputs_7_55_port, 
                           shift_out(54) => negative_inputs_7_54_port, 
                           shift_out(53) => negative_inputs_7_53_port, 
                           shift_out(52) => negative_inputs_7_52_port, 
                           shift_out(51) => negative_inputs_7_51_port, 
                           shift_out(50) => negative_inputs_7_50_port, 
                           shift_out(49) => negative_inputs_7_49_port, 
                           shift_out(48) => negative_inputs_7_48_port, 
                           shift_out(47) => negative_inputs_7_47_port, 
                           shift_out(46) => negative_inputs_7_46_port, 
                           shift_out(45) => negative_inputs_7_45_port, 
                           shift_out(44) => negative_inputs_7_44_port, 
                           shift_out(43) => negative_inputs_7_43_port, 
                           shift_out(42) => negative_inputs_7_42_port, 
                           shift_out(41) => negative_inputs_7_41_port, 
                           shift_out(40) => negative_inputs_7_40_port, 
                           shift_out(39) => negative_inputs_7_39_port, 
                           shift_out(38) => negative_inputs_7_38_port, 
                           shift_out(37) => negative_inputs_7_37_port, 
                           shift_out(36) => negative_inputs_7_36_port, 
                           shift_out(35) => negative_inputs_7_35_port, 
                           shift_out(34) => negative_inputs_7_34_port, 
                           shift_out(33) => negative_inputs_7_33_port, 
                           shift_out(32) => negative_inputs_7_32_port, 
                           shift_out(31) => negative_inputs_7_31_port, 
                           shift_out(30) => negative_inputs_7_30_port, 
                           shift_out(29) => negative_inputs_7_29_port, 
                           shift_out(28) => negative_inputs_7_28_port, 
                           shift_out(27) => negative_inputs_7_27_port, 
                           shift_out(26) => negative_inputs_7_26_port, 
                           shift_out(25) => negative_inputs_7_25_port, 
                           shift_out(24) => negative_inputs_7_24_port, 
                           shift_out(23) => negative_inputs_7_23_port, 
                           shift_out(22) => negative_inputs_7_22_port, 
                           shift_out(21) => negative_inputs_7_21_port, 
                           shift_out(20) => negative_inputs_7_20_port, 
                           shift_out(19) => negative_inputs_7_19_port, 
                           shift_out(18) => negative_inputs_7_18_port, 
                           shift_out(17) => negative_inputs_7_17_port, 
                           shift_out(16) => negative_inputs_7_16_port, 
                           shift_out(15) => negative_inputs_7_15_port, 
                           shift_out(14) => negative_inputs_7_14_port, 
                           shift_out(13) => negative_inputs_7_13_port, 
                           shift_out(12) => negative_inputs_7_12_port, 
                           shift_out(11) => negative_inputs_7_11_port, 
                           shift_out(10) => negative_inputs_7_10_port, 
                           shift_out(9) => negative_inputs_7_9_port, 
                           shift_out(8) => negative_inputs_7_8_port, 
                           shift_out(7) => negative_inputs_7_7_port, 
                           shift_out(6) => negative_inputs_7_6_port, 
                           shift_out(5) => negative_inputs_7_5_port, 
                           shift_out(4) => negative_inputs_7_4_port, 
                           shift_out(3) => negative_inputs_7_3_port, 
                           shift_out(2) => negative_inputs_7_2_port, 
                           shift_out(1) => negative_inputs_7_1_port, 
                           shift_out(0) => n_1102);
   shifted_neg_8 : leftshifter_NbitShifter64_87 port map( shift_in(63) => 
                           negative_inputs_7_63_port, shift_in(62) => 
                           negative_inputs_7_62_port, shift_in(61) => 
                           negative_inputs_7_61_port, shift_in(60) => 
                           negative_inputs_7_60_port, shift_in(59) => 
                           negative_inputs_7_59_port, shift_in(58) => 
                           negative_inputs_7_58_port, shift_in(57) => 
                           negative_inputs_7_57_port, shift_in(56) => 
                           negative_inputs_7_56_port, shift_in(55) => 
                           negative_inputs_7_55_port, shift_in(54) => 
                           negative_inputs_7_54_port, shift_in(53) => 
                           negative_inputs_7_53_port, shift_in(52) => 
                           negative_inputs_7_52_port, shift_in(51) => 
                           negative_inputs_7_51_port, shift_in(50) => 
                           negative_inputs_7_50_port, shift_in(49) => 
                           negative_inputs_7_49_port, shift_in(48) => 
                           negative_inputs_7_48_port, shift_in(47) => n119, 
                           shift_in(46) => negative_inputs_7_46_port, 
                           shift_in(45) => negative_inputs_7_45_port, 
                           shift_in(44) => negative_inputs_7_44_port, 
                           shift_in(43) => negative_inputs_7_43_port, 
                           shift_in(42) => negative_inputs_7_42_port, 
                           shift_in(41) => negative_inputs_7_41_port, 
                           shift_in(40) => negative_inputs_7_40_port, 
                           shift_in(39) => negative_inputs_7_39_port, 
                           shift_in(38) => negative_inputs_7_38_port, 
                           shift_in(37) => negative_inputs_7_37_port, 
                           shift_in(36) => negative_inputs_7_36_port, 
                           shift_in(35) => negative_inputs_7_35_port, 
                           shift_in(34) => negative_inputs_7_34_port, 
                           shift_in(33) => negative_inputs_7_33_port, 
                           shift_in(32) => negative_inputs_7_32_port, 
                           shift_in(31) => negative_inputs_7_31_port, 
                           shift_in(30) => negative_inputs_7_30_port, 
                           shift_in(29) => negative_inputs_7_29_port, 
                           shift_in(28) => negative_inputs_7_28_port, 
                           shift_in(27) => negative_inputs_7_27_port, 
                           shift_in(26) => negative_inputs_7_26_port, 
                           shift_in(25) => negative_inputs_7_25_port, 
                           shift_in(24) => negative_inputs_7_24_port, 
                           shift_in(23) => negative_inputs_7_23_port, 
                           shift_in(22) => negative_inputs_7_22_port, 
                           shift_in(21) => negative_inputs_7_21_port, 
                           shift_in(20) => negative_inputs_7_20_port, 
                           shift_in(19) => negative_inputs_7_19_port, 
                           shift_in(18) => negative_inputs_7_18_port, 
                           shift_in(17) => negative_inputs_7_17_port, 
                           shift_in(16) => negative_inputs_7_16_port, 
                           shift_in(15) => negative_inputs_7_15_port, 
                           shift_in(14) => negative_inputs_7_14_port, 
                           shift_in(13) => negative_inputs_7_13_port, 
                           shift_in(12) => negative_inputs_7_12_port, 
                           shift_in(11) => negative_inputs_7_11_port, 
                           shift_in(10) => negative_inputs_7_10_port, 
                           shift_in(9) => negative_inputs_7_9_port, shift_in(8)
                           => negative_inputs_7_8_port, shift_in(7) => 
                           negative_inputs_7_7_port, shift_in(6) => 
                           negative_inputs_7_6_port, shift_in(5) => 
                           negative_inputs_7_5_port, shift_in(4) => 
                           negative_inputs_7_4_port, shift_in(3) => 
                           negative_inputs_7_3_port, shift_in(2) => 
                           negative_inputs_7_2_port, shift_in(1) => 
                           negative_inputs_7_1_port, shift_in(0) => n8, 
                           shift_out(63) => negative_inputs_8_63_port, 
                           shift_out(62) => negative_inputs_8_62_port, 
                           shift_out(61) => negative_inputs_8_61_port, 
                           shift_out(60) => negative_inputs_8_60_port, 
                           shift_out(59) => negative_inputs_8_59_port, 
                           shift_out(58) => negative_inputs_8_58_port, 
                           shift_out(57) => negative_inputs_8_57_port, 
                           shift_out(56) => negative_inputs_8_56_port, 
                           shift_out(55) => negative_inputs_8_55_port, 
                           shift_out(54) => negative_inputs_8_54_port, 
                           shift_out(53) => negative_inputs_8_53_port, 
                           shift_out(52) => negative_inputs_8_52_port, 
                           shift_out(51) => negative_inputs_8_51_port, 
                           shift_out(50) => negative_inputs_8_50_port, 
                           shift_out(49) => negative_inputs_8_49_port, 
                           shift_out(48) => negative_inputs_8_48_port, 
                           shift_out(47) => negative_inputs_8_47_port, 
                           shift_out(46) => negative_inputs_8_46_port, 
                           shift_out(45) => negative_inputs_8_45_port, 
                           shift_out(44) => negative_inputs_8_44_port, 
                           shift_out(43) => negative_inputs_8_43_port, 
                           shift_out(42) => negative_inputs_8_42_port, 
                           shift_out(41) => negative_inputs_8_41_port, 
                           shift_out(40) => negative_inputs_8_40_port, 
                           shift_out(39) => negative_inputs_8_39_port, 
                           shift_out(38) => negative_inputs_8_38_port, 
                           shift_out(37) => negative_inputs_8_37_port, 
                           shift_out(36) => negative_inputs_8_36_port, 
                           shift_out(35) => negative_inputs_8_35_port, 
                           shift_out(34) => negative_inputs_8_34_port, 
                           shift_out(33) => negative_inputs_8_33_port, 
                           shift_out(32) => negative_inputs_8_32_port, 
                           shift_out(31) => negative_inputs_8_31_port, 
                           shift_out(30) => negative_inputs_8_30_port, 
                           shift_out(29) => negative_inputs_8_29_port, 
                           shift_out(28) => negative_inputs_8_28_port, 
                           shift_out(27) => negative_inputs_8_27_port, 
                           shift_out(26) => negative_inputs_8_26_port, 
                           shift_out(25) => negative_inputs_8_25_port, 
                           shift_out(24) => negative_inputs_8_24_port, 
                           shift_out(23) => negative_inputs_8_23_port, 
                           shift_out(22) => negative_inputs_8_22_port, 
                           shift_out(21) => negative_inputs_8_21_port, 
                           shift_out(20) => negative_inputs_8_20_port, 
                           shift_out(19) => negative_inputs_8_19_port, 
                           shift_out(18) => negative_inputs_8_18_port, 
                           shift_out(17) => negative_inputs_8_17_port, 
                           shift_out(16) => negative_inputs_8_16_port, 
                           shift_out(15) => negative_inputs_8_15_port, 
                           shift_out(14) => negative_inputs_8_14_port, 
                           shift_out(13) => negative_inputs_8_13_port, 
                           shift_out(12) => negative_inputs_8_12_port, 
                           shift_out(11) => negative_inputs_8_11_port, 
                           shift_out(10) => negative_inputs_8_10_port, 
                           shift_out(9) => negative_inputs_8_9_port, 
                           shift_out(8) => negative_inputs_8_8_port, 
                           shift_out(7) => negative_inputs_8_7_port, 
                           shift_out(6) => negative_inputs_8_6_port, 
                           shift_out(5) => negative_inputs_8_5_port, 
                           shift_out(4) => negative_inputs_8_4_port, 
                           shift_out(3) => negative_inputs_8_3_port, 
                           shift_out(2) => negative_inputs_8_2_port, 
                           shift_out(1) => negative_inputs_8_1_port, 
                           shift_out(0) => n_1103);
   shifted_neg_9 : leftshifter_NbitShifter64_86 port map( shift_in(63) => 
                           negative_inputs_8_63_port, shift_in(62) => 
                           negative_inputs_8_62_port, shift_in(61) => 
                           negative_inputs_8_61_port, shift_in(60) => 
                           negative_inputs_8_60_port, shift_in(59) => 
                           negative_inputs_8_59_port, shift_in(58) => 
                           negative_inputs_8_58_port, shift_in(57) => 
                           negative_inputs_8_57_port, shift_in(56) => 
                           negative_inputs_8_56_port, shift_in(55) => 
                           negative_inputs_8_55_port, shift_in(54) => 
                           negative_inputs_8_54_port, shift_in(53) => 
                           negative_inputs_8_53_port, shift_in(52) => 
                           negative_inputs_8_52_port, shift_in(51) => 
                           negative_inputs_8_51_port, shift_in(50) => 
                           negative_inputs_8_50_port, shift_in(49) => 
                           negative_inputs_8_49_port, shift_in(48) => 
                           negative_inputs_8_48_port, shift_in(47) => n118, 
                           shift_in(46) => negative_inputs_8_46_port, 
                           shift_in(45) => negative_inputs_8_45_port, 
                           shift_in(44) => negative_inputs_8_44_port, 
                           shift_in(43) => negative_inputs_8_43_port, 
                           shift_in(42) => negative_inputs_8_42_port, 
                           shift_in(41) => negative_inputs_8_41_port, 
                           shift_in(40) => negative_inputs_8_40_port, 
                           shift_in(39) => negative_inputs_8_39_port, 
                           shift_in(38) => negative_inputs_8_38_port, 
                           shift_in(37) => negative_inputs_8_37_port, 
                           shift_in(36) => negative_inputs_8_36_port, 
                           shift_in(35) => negative_inputs_8_35_port, 
                           shift_in(34) => negative_inputs_8_34_port, 
                           shift_in(33) => negative_inputs_8_33_port, 
                           shift_in(32) => negative_inputs_8_32_port, 
                           shift_in(31) => negative_inputs_8_31_port, 
                           shift_in(30) => negative_inputs_8_30_port, 
                           shift_in(29) => negative_inputs_8_29_port, 
                           shift_in(28) => negative_inputs_8_28_port, 
                           shift_in(27) => negative_inputs_8_27_port, 
                           shift_in(26) => negative_inputs_8_26_port, 
                           shift_in(25) => negative_inputs_8_25_port, 
                           shift_in(24) => negative_inputs_8_24_port, 
                           shift_in(23) => negative_inputs_8_23_port, 
                           shift_in(22) => negative_inputs_8_22_port, 
                           shift_in(21) => negative_inputs_8_21_port, 
                           shift_in(20) => negative_inputs_8_20_port, 
                           shift_in(19) => negative_inputs_8_19_port, 
                           shift_in(18) => negative_inputs_8_18_port, 
                           shift_in(17) => negative_inputs_8_17_port, 
                           shift_in(16) => negative_inputs_8_16_port, 
                           shift_in(15) => negative_inputs_8_15_port, 
                           shift_in(14) => negative_inputs_8_14_port, 
                           shift_in(13) => negative_inputs_8_13_port, 
                           shift_in(12) => negative_inputs_8_12_port, 
                           shift_in(11) => negative_inputs_8_11_port, 
                           shift_in(10) => negative_inputs_8_10_port, 
                           shift_in(9) => negative_inputs_8_9_port, shift_in(8)
                           => negative_inputs_8_8_port, shift_in(7) => 
                           negative_inputs_8_7_port, shift_in(6) => 
                           negative_inputs_8_6_port, shift_in(5) => 
                           negative_inputs_8_5_port, shift_in(4) => 
                           negative_inputs_8_4_port, shift_in(3) => 
                           negative_inputs_8_3_port, shift_in(2) => 
                           negative_inputs_8_2_port, shift_in(1) => 
                           negative_inputs_8_1_port, shift_in(0) => n8, 
                           shift_out(63) => negative_inputs_9_63_port, 
                           shift_out(62) => negative_inputs_9_62_port, 
                           shift_out(61) => negative_inputs_9_61_port, 
                           shift_out(60) => negative_inputs_9_60_port, 
                           shift_out(59) => negative_inputs_9_59_port, 
                           shift_out(58) => negative_inputs_9_58_port, 
                           shift_out(57) => negative_inputs_9_57_port, 
                           shift_out(56) => negative_inputs_9_56_port, 
                           shift_out(55) => negative_inputs_9_55_port, 
                           shift_out(54) => negative_inputs_9_54_port, 
                           shift_out(53) => negative_inputs_9_53_port, 
                           shift_out(52) => negative_inputs_9_52_port, 
                           shift_out(51) => negative_inputs_9_51_port, 
                           shift_out(50) => negative_inputs_9_50_port, 
                           shift_out(49) => negative_inputs_9_49_port, 
                           shift_out(48) => negative_inputs_9_48_port, 
                           shift_out(47) => negative_inputs_9_47_port, 
                           shift_out(46) => negative_inputs_9_46_port, 
                           shift_out(45) => negative_inputs_9_45_port, 
                           shift_out(44) => negative_inputs_9_44_port, 
                           shift_out(43) => negative_inputs_9_43_port, 
                           shift_out(42) => negative_inputs_9_42_port, 
                           shift_out(41) => negative_inputs_9_41_port, 
                           shift_out(40) => negative_inputs_9_40_port, 
                           shift_out(39) => negative_inputs_9_39_port, 
                           shift_out(38) => negative_inputs_9_38_port, 
                           shift_out(37) => negative_inputs_9_37_port, 
                           shift_out(36) => negative_inputs_9_36_port, 
                           shift_out(35) => negative_inputs_9_35_port, 
                           shift_out(34) => negative_inputs_9_34_port, 
                           shift_out(33) => negative_inputs_9_33_port, 
                           shift_out(32) => negative_inputs_9_32_port, 
                           shift_out(31) => negative_inputs_9_31_port, 
                           shift_out(30) => negative_inputs_9_30_port, 
                           shift_out(29) => negative_inputs_9_29_port, 
                           shift_out(28) => negative_inputs_9_28_port, 
                           shift_out(27) => negative_inputs_9_27_port, 
                           shift_out(26) => negative_inputs_9_26_port, 
                           shift_out(25) => negative_inputs_9_25_port, 
                           shift_out(24) => negative_inputs_9_24_port, 
                           shift_out(23) => negative_inputs_9_23_port, 
                           shift_out(22) => negative_inputs_9_22_port, 
                           shift_out(21) => negative_inputs_9_21_port, 
                           shift_out(20) => negative_inputs_9_20_port, 
                           shift_out(19) => negative_inputs_9_19_port, 
                           shift_out(18) => negative_inputs_9_18_port, 
                           shift_out(17) => negative_inputs_9_17_port, 
                           shift_out(16) => negative_inputs_9_16_port, 
                           shift_out(15) => negative_inputs_9_15_port, 
                           shift_out(14) => negative_inputs_9_14_port, 
                           shift_out(13) => negative_inputs_9_13_port, 
                           shift_out(12) => negative_inputs_9_12_port, 
                           shift_out(11) => negative_inputs_9_11_port, 
                           shift_out(10) => negative_inputs_9_10_port, 
                           shift_out(9) => negative_inputs_9_9_port, 
                           shift_out(8) => negative_inputs_9_8_port, 
                           shift_out(7) => negative_inputs_9_7_port, 
                           shift_out(6) => negative_inputs_9_6_port, 
                           shift_out(5) => negative_inputs_9_5_port, 
                           shift_out(4) => negative_inputs_9_4_port, 
                           shift_out(3) => negative_inputs_9_3_port, 
                           shift_out(2) => negative_inputs_9_2_port, 
                           shift_out(1) => negative_inputs_9_1_port, 
                           shift_out(0) => n_1104);
   shifted_neg_10 : leftshifter_NbitShifter64_85 port map( shift_in(63) => 
                           negative_inputs_9_63_port, shift_in(62) => 
                           negative_inputs_9_62_port, shift_in(61) => 
                           negative_inputs_9_61_port, shift_in(60) => 
                           negative_inputs_9_60_port, shift_in(59) => 
                           negative_inputs_9_59_port, shift_in(58) => 
                           negative_inputs_9_58_port, shift_in(57) => 
                           negative_inputs_9_57_port, shift_in(56) => 
                           negative_inputs_9_56_port, shift_in(55) => 
                           negative_inputs_9_55_port, shift_in(54) => 
                           negative_inputs_9_54_port, shift_in(53) => 
                           negative_inputs_9_53_port, shift_in(52) => 
                           negative_inputs_9_52_port, shift_in(51) => 
                           negative_inputs_9_51_port, shift_in(50) => 
                           negative_inputs_9_50_port, shift_in(49) => 
                           negative_inputs_9_49_port, shift_in(48) => 
                           negative_inputs_9_48_port, shift_in(47) => n117, 
                           shift_in(46) => negative_inputs_9_46_port, 
                           shift_in(45) => negative_inputs_9_45_port, 
                           shift_in(44) => negative_inputs_9_44_port, 
                           shift_in(43) => negative_inputs_9_43_port, 
                           shift_in(42) => negative_inputs_9_42_port, 
                           shift_in(41) => negative_inputs_9_41_port, 
                           shift_in(40) => negative_inputs_9_40_port, 
                           shift_in(39) => negative_inputs_9_39_port, 
                           shift_in(38) => negative_inputs_9_38_port, 
                           shift_in(37) => negative_inputs_9_37_port, 
                           shift_in(36) => negative_inputs_9_36_port, 
                           shift_in(35) => negative_inputs_9_35_port, 
                           shift_in(34) => negative_inputs_9_34_port, 
                           shift_in(33) => negative_inputs_9_33_port, 
                           shift_in(32) => negative_inputs_9_32_port, 
                           shift_in(31) => negative_inputs_9_31_port, 
                           shift_in(30) => negative_inputs_9_30_port, 
                           shift_in(29) => negative_inputs_9_29_port, 
                           shift_in(28) => negative_inputs_9_28_port, 
                           shift_in(27) => negative_inputs_9_27_port, 
                           shift_in(26) => negative_inputs_9_26_port, 
                           shift_in(25) => negative_inputs_9_25_port, 
                           shift_in(24) => negative_inputs_9_24_port, 
                           shift_in(23) => negative_inputs_9_23_port, 
                           shift_in(22) => negative_inputs_9_22_port, 
                           shift_in(21) => negative_inputs_9_21_port, 
                           shift_in(20) => negative_inputs_9_20_port, 
                           shift_in(19) => negative_inputs_9_19_port, 
                           shift_in(18) => negative_inputs_9_18_port, 
                           shift_in(17) => negative_inputs_9_17_port, 
                           shift_in(16) => negative_inputs_9_16_port, 
                           shift_in(15) => negative_inputs_9_15_port, 
                           shift_in(14) => negative_inputs_9_14_port, 
                           shift_in(13) => negative_inputs_9_13_port, 
                           shift_in(12) => negative_inputs_9_12_port, 
                           shift_in(11) => negative_inputs_9_11_port, 
                           shift_in(10) => negative_inputs_9_10_port, 
                           shift_in(9) => negative_inputs_9_9_port, shift_in(8)
                           => negative_inputs_9_8_port, shift_in(7) => 
                           negative_inputs_9_7_port, shift_in(6) => 
                           negative_inputs_9_6_port, shift_in(5) => 
                           negative_inputs_9_5_port, shift_in(4) => 
                           negative_inputs_9_4_port, shift_in(3) => 
                           negative_inputs_9_3_port, shift_in(2) => 
                           negative_inputs_9_2_port, shift_in(1) => 
                           negative_inputs_9_1_port, shift_in(0) => n8, 
                           shift_out(63) => negative_inputs_10_63_port, 
                           shift_out(62) => negative_inputs_10_62_port, 
                           shift_out(61) => negative_inputs_10_61_port, 
                           shift_out(60) => negative_inputs_10_60_port, 
                           shift_out(59) => negative_inputs_10_59_port, 
                           shift_out(58) => negative_inputs_10_58_port, 
                           shift_out(57) => negative_inputs_10_57_port, 
                           shift_out(56) => negative_inputs_10_56_port, 
                           shift_out(55) => negative_inputs_10_55_port, 
                           shift_out(54) => negative_inputs_10_54_port, 
                           shift_out(53) => negative_inputs_10_53_port, 
                           shift_out(52) => negative_inputs_10_52_port, 
                           shift_out(51) => negative_inputs_10_51_port, 
                           shift_out(50) => negative_inputs_10_50_port, 
                           shift_out(49) => negative_inputs_10_49_port, 
                           shift_out(48) => negative_inputs_10_48_port, 
                           shift_out(47) => negative_inputs_10_47_port, 
                           shift_out(46) => negative_inputs_10_46_port, 
                           shift_out(45) => negative_inputs_10_45_port, 
                           shift_out(44) => negative_inputs_10_44_port, 
                           shift_out(43) => negative_inputs_10_43_port, 
                           shift_out(42) => negative_inputs_10_42_port, 
                           shift_out(41) => negative_inputs_10_41_port, 
                           shift_out(40) => negative_inputs_10_40_port, 
                           shift_out(39) => negative_inputs_10_39_port, 
                           shift_out(38) => negative_inputs_10_38_port, 
                           shift_out(37) => negative_inputs_10_37_port, 
                           shift_out(36) => negative_inputs_10_36_port, 
                           shift_out(35) => negative_inputs_10_35_port, 
                           shift_out(34) => negative_inputs_10_34_port, 
                           shift_out(33) => negative_inputs_10_33_port, 
                           shift_out(32) => negative_inputs_10_32_port, 
                           shift_out(31) => negative_inputs_10_31_port, 
                           shift_out(30) => negative_inputs_10_30_port, 
                           shift_out(29) => negative_inputs_10_29_port, 
                           shift_out(28) => negative_inputs_10_28_port, 
                           shift_out(27) => negative_inputs_10_27_port, 
                           shift_out(26) => negative_inputs_10_26_port, 
                           shift_out(25) => negative_inputs_10_25_port, 
                           shift_out(24) => negative_inputs_10_24_port, 
                           shift_out(23) => negative_inputs_10_23_port, 
                           shift_out(22) => negative_inputs_10_22_port, 
                           shift_out(21) => negative_inputs_10_21_port, 
                           shift_out(20) => negative_inputs_10_20_port, 
                           shift_out(19) => negative_inputs_10_19_port, 
                           shift_out(18) => negative_inputs_10_18_port, 
                           shift_out(17) => negative_inputs_10_17_port, 
                           shift_out(16) => negative_inputs_10_16_port, 
                           shift_out(15) => negative_inputs_10_15_port, 
                           shift_out(14) => negative_inputs_10_14_port, 
                           shift_out(13) => negative_inputs_10_13_port, 
                           shift_out(12) => negative_inputs_10_12_port, 
                           shift_out(11) => negative_inputs_10_11_port, 
                           shift_out(10) => negative_inputs_10_10_port, 
                           shift_out(9) => negative_inputs_10_9_port, 
                           shift_out(8) => negative_inputs_10_8_port, 
                           shift_out(7) => negative_inputs_10_7_port, 
                           shift_out(6) => negative_inputs_10_6_port, 
                           shift_out(5) => negative_inputs_10_5_port, 
                           shift_out(4) => negative_inputs_10_4_port, 
                           shift_out(3) => negative_inputs_10_3_port, 
                           shift_out(2) => negative_inputs_10_2_port, 
                           shift_out(1) => negative_inputs_10_1_port, 
                           shift_out(0) => n_1105);
   shifted_neg_11 : leftshifter_NbitShifter64_84 port map( shift_in(63) => 
                           negative_inputs_10_63_port, shift_in(62) => 
                           negative_inputs_10_62_port, shift_in(61) => 
                           negative_inputs_10_61_port, shift_in(60) => 
                           negative_inputs_10_60_port, shift_in(59) => 
                           negative_inputs_10_59_port, shift_in(58) => 
                           negative_inputs_10_58_port, shift_in(57) => 
                           negative_inputs_10_57_port, shift_in(56) => 
                           negative_inputs_10_56_port, shift_in(55) => 
                           negative_inputs_10_55_port, shift_in(54) => 
                           negative_inputs_10_54_port, shift_in(53) => 
                           negative_inputs_10_53_port, shift_in(52) => 
                           negative_inputs_10_52_port, shift_in(51) => 
                           negative_inputs_10_51_port, shift_in(50) => 
                           negative_inputs_10_50_port, shift_in(49) => 
                           negative_inputs_10_49_port, shift_in(48) => 
                           negative_inputs_10_48_port, shift_in(47) => n116, 
                           shift_in(46) => negative_inputs_10_46_port, 
                           shift_in(45) => negative_inputs_10_45_port, 
                           shift_in(44) => negative_inputs_10_44_port, 
                           shift_in(43) => negative_inputs_10_43_port, 
                           shift_in(42) => negative_inputs_10_42_port, 
                           shift_in(41) => negative_inputs_10_41_port, 
                           shift_in(40) => negative_inputs_10_40_port, 
                           shift_in(39) => negative_inputs_10_39_port, 
                           shift_in(38) => negative_inputs_10_38_port, 
                           shift_in(37) => negative_inputs_10_37_port, 
                           shift_in(36) => negative_inputs_10_36_port, 
                           shift_in(35) => negative_inputs_10_35_port, 
                           shift_in(34) => negative_inputs_10_34_port, 
                           shift_in(33) => negative_inputs_10_33_port, 
                           shift_in(32) => negative_inputs_10_32_port, 
                           shift_in(31) => negative_inputs_10_31_port, 
                           shift_in(30) => negative_inputs_10_30_port, 
                           shift_in(29) => negative_inputs_10_29_port, 
                           shift_in(28) => negative_inputs_10_28_port, 
                           shift_in(27) => negative_inputs_10_27_port, 
                           shift_in(26) => negative_inputs_10_26_port, 
                           shift_in(25) => negative_inputs_10_25_port, 
                           shift_in(24) => negative_inputs_10_24_port, 
                           shift_in(23) => negative_inputs_10_23_port, 
                           shift_in(22) => negative_inputs_10_22_port, 
                           shift_in(21) => negative_inputs_10_21_port, 
                           shift_in(20) => negative_inputs_10_20_port, 
                           shift_in(19) => negative_inputs_10_19_port, 
                           shift_in(18) => negative_inputs_10_18_port, 
                           shift_in(17) => negative_inputs_10_17_port, 
                           shift_in(16) => negative_inputs_10_16_port, 
                           shift_in(15) => negative_inputs_10_15_port, 
                           shift_in(14) => negative_inputs_10_14_port, 
                           shift_in(13) => negative_inputs_10_13_port, 
                           shift_in(12) => negative_inputs_10_12_port, 
                           shift_in(11) => negative_inputs_10_11_port, 
                           shift_in(10) => negative_inputs_10_10_port, 
                           shift_in(9) => negative_inputs_10_9_port, 
                           shift_in(8) => negative_inputs_10_8_port, 
                           shift_in(7) => negative_inputs_10_7_port, 
                           shift_in(6) => negative_inputs_10_6_port, 
                           shift_in(5) => negative_inputs_10_5_port, 
                           shift_in(4) => negative_inputs_10_4_port, 
                           shift_in(3) => negative_inputs_10_3_port, 
                           shift_in(2) => negative_inputs_10_2_port, 
                           shift_in(1) => negative_inputs_10_1_port, 
                           shift_in(0) => n8, shift_out(63) => 
                           negative_inputs_11_63_port, shift_out(62) => 
                           negative_inputs_11_62_port, shift_out(61) => 
                           negative_inputs_11_61_port, shift_out(60) => 
                           negative_inputs_11_60_port, shift_out(59) => 
                           negative_inputs_11_59_port, shift_out(58) => 
                           negative_inputs_11_58_port, shift_out(57) => 
                           negative_inputs_11_57_port, shift_out(56) => 
                           negative_inputs_11_56_port, shift_out(55) => 
                           negative_inputs_11_55_port, shift_out(54) => 
                           negative_inputs_11_54_port, shift_out(53) => 
                           negative_inputs_11_53_port, shift_out(52) => 
                           negative_inputs_11_52_port, shift_out(51) => 
                           negative_inputs_11_51_port, shift_out(50) => 
                           negative_inputs_11_50_port, shift_out(49) => 
                           negative_inputs_11_49_port, shift_out(48) => 
                           negative_inputs_11_48_port, shift_out(47) => 
                           negative_inputs_11_47_port, shift_out(46) => 
                           negative_inputs_11_46_port, shift_out(45) => 
                           negative_inputs_11_45_port, shift_out(44) => 
                           negative_inputs_11_44_port, shift_out(43) => 
                           negative_inputs_11_43_port, shift_out(42) => 
                           negative_inputs_11_42_port, shift_out(41) => 
                           negative_inputs_11_41_port, shift_out(40) => 
                           negative_inputs_11_40_port, shift_out(39) => 
                           negative_inputs_11_39_port, shift_out(38) => 
                           negative_inputs_11_38_port, shift_out(37) => 
                           negative_inputs_11_37_port, shift_out(36) => 
                           negative_inputs_11_36_port, shift_out(35) => 
                           negative_inputs_11_35_port, shift_out(34) => 
                           negative_inputs_11_34_port, shift_out(33) => 
                           negative_inputs_11_33_port, shift_out(32) => 
                           negative_inputs_11_32_port, shift_out(31) => 
                           negative_inputs_11_31_port, shift_out(30) => 
                           negative_inputs_11_30_port, shift_out(29) => 
                           negative_inputs_11_29_port, shift_out(28) => 
                           negative_inputs_11_28_port, shift_out(27) => 
                           negative_inputs_11_27_port, shift_out(26) => 
                           negative_inputs_11_26_port, shift_out(25) => 
                           negative_inputs_11_25_port, shift_out(24) => 
                           negative_inputs_11_24_port, shift_out(23) => 
                           negative_inputs_11_23_port, shift_out(22) => 
                           negative_inputs_11_22_port, shift_out(21) => 
                           negative_inputs_11_21_port, shift_out(20) => 
                           negative_inputs_11_20_port, shift_out(19) => 
                           negative_inputs_11_19_port, shift_out(18) => 
                           negative_inputs_11_18_port, shift_out(17) => 
                           negative_inputs_11_17_port, shift_out(16) => 
                           negative_inputs_11_16_port, shift_out(15) => 
                           negative_inputs_11_15_port, shift_out(14) => 
                           negative_inputs_11_14_port, shift_out(13) => 
                           negative_inputs_11_13_port, shift_out(12) => 
                           negative_inputs_11_12_port, shift_out(11) => 
                           negative_inputs_11_11_port, shift_out(10) => 
                           negative_inputs_11_10_port, shift_out(9) => 
                           negative_inputs_11_9_port, shift_out(8) => 
                           negative_inputs_11_8_port, shift_out(7) => 
                           negative_inputs_11_7_port, shift_out(6) => 
                           negative_inputs_11_6_port, shift_out(5) => 
                           negative_inputs_11_5_port, shift_out(4) => 
                           negative_inputs_11_4_port, shift_out(3) => 
                           negative_inputs_11_3_port, shift_out(2) => 
                           negative_inputs_11_2_port, shift_out(1) => 
                           negative_inputs_11_1_port, shift_out(0) => n_1106);
   shifted_neg_12 : leftshifter_NbitShifter64_83 port map( shift_in(63) => 
                           negative_inputs_11_63_port, shift_in(62) => 
                           negative_inputs_11_62_port, shift_in(61) => 
                           negative_inputs_11_61_port, shift_in(60) => 
                           negative_inputs_11_60_port, shift_in(59) => 
                           negative_inputs_11_59_port, shift_in(58) => 
                           negative_inputs_11_58_port, shift_in(57) => 
                           negative_inputs_11_57_port, shift_in(56) => 
                           negative_inputs_11_56_port, shift_in(55) => 
                           negative_inputs_11_55_port, shift_in(54) => 
                           negative_inputs_11_54_port, shift_in(53) => 
                           negative_inputs_11_53_port, shift_in(52) => 
                           negative_inputs_11_52_port, shift_in(51) => 
                           negative_inputs_11_51_port, shift_in(50) => 
                           negative_inputs_11_50_port, shift_in(49) => 
                           negative_inputs_11_49_port, shift_in(48) => 
                           negative_inputs_11_48_port, shift_in(47) => n115, 
                           shift_in(46) => negative_inputs_11_46_port, 
                           shift_in(45) => negative_inputs_11_45_port, 
                           shift_in(44) => negative_inputs_11_44_port, 
                           shift_in(43) => negative_inputs_11_43_port, 
                           shift_in(42) => negative_inputs_11_42_port, 
                           shift_in(41) => negative_inputs_11_41_port, 
                           shift_in(40) => negative_inputs_11_40_port, 
                           shift_in(39) => negative_inputs_11_39_port, 
                           shift_in(38) => negative_inputs_11_38_port, 
                           shift_in(37) => negative_inputs_11_37_port, 
                           shift_in(36) => negative_inputs_11_36_port, 
                           shift_in(35) => negative_inputs_11_35_port, 
                           shift_in(34) => negative_inputs_11_34_port, 
                           shift_in(33) => negative_inputs_11_33_port, 
                           shift_in(32) => negative_inputs_11_32_port, 
                           shift_in(31) => negative_inputs_11_31_port, 
                           shift_in(30) => negative_inputs_11_30_port, 
                           shift_in(29) => negative_inputs_11_29_port, 
                           shift_in(28) => negative_inputs_11_28_port, 
                           shift_in(27) => negative_inputs_11_27_port, 
                           shift_in(26) => negative_inputs_11_26_port, 
                           shift_in(25) => negative_inputs_11_25_port, 
                           shift_in(24) => negative_inputs_11_24_port, 
                           shift_in(23) => negative_inputs_11_23_port, 
                           shift_in(22) => negative_inputs_11_22_port, 
                           shift_in(21) => negative_inputs_11_21_port, 
                           shift_in(20) => negative_inputs_11_20_port, 
                           shift_in(19) => negative_inputs_11_19_port, 
                           shift_in(18) => negative_inputs_11_18_port, 
                           shift_in(17) => negative_inputs_11_17_port, 
                           shift_in(16) => negative_inputs_11_16_port, 
                           shift_in(15) => negative_inputs_11_15_port, 
                           shift_in(14) => negative_inputs_11_14_port, 
                           shift_in(13) => negative_inputs_11_13_port, 
                           shift_in(12) => negative_inputs_11_12_port, 
                           shift_in(11) => negative_inputs_11_11_port, 
                           shift_in(10) => negative_inputs_11_10_port, 
                           shift_in(9) => negative_inputs_11_9_port, 
                           shift_in(8) => negative_inputs_11_8_port, 
                           shift_in(7) => negative_inputs_11_7_port, 
                           shift_in(6) => negative_inputs_11_6_port, 
                           shift_in(5) => negative_inputs_11_5_port, 
                           shift_in(4) => negative_inputs_11_4_port, 
                           shift_in(3) => negative_inputs_11_3_port, 
                           shift_in(2) => negative_inputs_11_2_port, 
                           shift_in(1) => negative_inputs_11_1_port, 
                           shift_in(0) => n8, shift_out(63) => 
                           negative_inputs_12_63_port, shift_out(62) => 
                           negative_inputs_12_62_port, shift_out(61) => 
                           negative_inputs_12_61_port, shift_out(60) => 
                           negative_inputs_12_60_port, shift_out(59) => 
                           negative_inputs_12_59_port, shift_out(58) => 
                           negative_inputs_12_58_port, shift_out(57) => 
                           negative_inputs_12_57_port, shift_out(56) => 
                           negative_inputs_12_56_port, shift_out(55) => 
                           negative_inputs_12_55_port, shift_out(54) => 
                           negative_inputs_12_54_port, shift_out(53) => 
                           negative_inputs_12_53_port, shift_out(52) => 
                           negative_inputs_12_52_port, shift_out(51) => 
                           negative_inputs_12_51_port, shift_out(50) => 
                           negative_inputs_12_50_port, shift_out(49) => 
                           negative_inputs_12_49_port, shift_out(48) => 
                           negative_inputs_12_48_port, shift_out(47) => 
                           negative_inputs_12_47_port, shift_out(46) => 
                           negative_inputs_12_46_port, shift_out(45) => 
                           negative_inputs_12_45_port, shift_out(44) => 
                           negative_inputs_12_44_port, shift_out(43) => 
                           negative_inputs_12_43_port, shift_out(42) => 
                           negative_inputs_12_42_port, shift_out(41) => 
                           negative_inputs_12_41_port, shift_out(40) => 
                           negative_inputs_12_40_port, shift_out(39) => 
                           negative_inputs_12_39_port, shift_out(38) => 
                           negative_inputs_12_38_port, shift_out(37) => 
                           negative_inputs_12_37_port, shift_out(36) => 
                           negative_inputs_12_36_port, shift_out(35) => 
                           negative_inputs_12_35_port, shift_out(34) => 
                           negative_inputs_12_34_port, shift_out(33) => 
                           negative_inputs_12_33_port, shift_out(32) => 
                           negative_inputs_12_32_port, shift_out(31) => 
                           negative_inputs_12_31_port, shift_out(30) => 
                           negative_inputs_12_30_port, shift_out(29) => 
                           negative_inputs_12_29_port, shift_out(28) => 
                           negative_inputs_12_28_port, shift_out(27) => 
                           negative_inputs_12_27_port, shift_out(26) => 
                           negative_inputs_12_26_port, shift_out(25) => 
                           negative_inputs_12_25_port, shift_out(24) => 
                           negative_inputs_12_24_port, shift_out(23) => 
                           negative_inputs_12_23_port, shift_out(22) => 
                           negative_inputs_12_22_port, shift_out(21) => 
                           negative_inputs_12_21_port, shift_out(20) => 
                           negative_inputs_12_20_port, shift_out(19) => 
                           negative_inputs_12_19_port, shift_out(18) => 
                           negative_inputs_12_18_port, shift_out(17) => 
                           negative_inputs_12_17_port, shift_out(16) => 
                           negative_inputs_12_16_port, shift_out(15) => 
                           negative_inputs_12_15_port, shift_out(14) => 
                           negative_inputs_12_14_port, shift_out(13) => 
                           negative_inputs_12_13_port, shift_out(12) => 
                           negative_inputs_12_12_port, shift_out(11) => 
                           negative_inputs_12_11_port, shift_out(10) => 
                           negative_inputs_12_10_port, shift_out(9) => 
                           negative_inputs_12_9_port, shift_out(8) => 
                           negative_inputs_12_8_port, shift_out(7) => 
                           negative_inputs_12_7_port, shift_out(6) => 
                           negative_inputs_12_6_port, shift_out(5) => 
                           negative_inputs_12_5_port, shift_out(4) => 
                           negative_inputs_12_4_port, shift_out(3) => 
                           negative_inputs_12_3_port, shift_out(2) => 
                           negative_inputs_12_2_port, shift_out(1) => 
                           negative_inputs_12_1_port, shift_out(0) => n_1107);
   shifted_neg_13 : leftshifter_NbitShifter64_82 port map( shift_in(63) => 
                           negative_inputs_12_63_port, shift_in(62) => 
                           negative_inputs_12_62_port, shift_in(61) => 
                           negative_inputs_12_61_port, shift_in(60) => 
                           negative_inputs_12_60_port, shift_in(59) => 
                           negative_inputs_12_59_port, shift_in(58) => 
                           negative_inputs_12_58_port, shift_in(57) => 
                           negative_inputs_12_57_port, shift_in(56) => 
                           negative_inputs_12_56_port, shift_in(55) => 
                           negative_inputs_12_55_port, shift_in(54) => 
                           negative_inputs_12_54_port, shift_in(53) => 
                           negative_inputs_12_53_port, shift_in(52) => 
                           negative_inputs_12_52_port, shift_in(51) => 
                           negative_inputs_12_51_port, shift_in(50) => 
                           negative_inputs_12_50_port, shift_in(49) => 
                           negative_inputs_12_49_port, shift_in(48) => 
                           negative_inputs_12_48_port, shift_in(47) => n113, 
                           shift_in(46) => negative_inputs_12_46_port, 
                           shift_in(45) => negative_inputs_12_45_port, 
                           shift_in(44) => negative_inputs_12_44_port, 
                           shift_in(43) => negative_inputs_12_43_port, 
                           shift_in(42) => negative_inputs_12_42_port, 
                           shift_in(41) => negative_inputs_12_41_port, 
                           shift_in(40) => negative_inputs_12_40_port, 
                           shift_in(39) => negative_inputs_12_39_port, 
                           shift_in(38) => negative_inputs_12_38_port, 
                           shift_in(37) => negative_inputs_12_37_port, 
                           shift_in(36) => negative_inputs_12_36_port, 
                           shift_in(35) => negative_inputs_12_35_port, 
                           shift_in(34) => negative_inputs_12_34_port, 
                           shift_in(33) => negative_inputs_12_33_port, 
                           shift_in(32) => negative_inputs_12_32_port, 
                           shift_in(31) => negative_inputs_12_31_port, 
                           shift_in(30) => negative_inputs_12_30_port, 
                           shift_in(29) => negative_inputs_12_29_port, 
                           shift_in(28) => negative_inputs_12_28_port, 
                           shift_in(27) => negative_inputs_12_27_port, 
                           shift_in(26) => negative_inputs_12_26_port, 
                           shift_in(25) => negative_inputs_12_25_port, 
                           shift_in(24) => negative_inputs_12_24_port, 
                           shift_in(23) => negative_inputs_12_23_port, 
                           shift_in(22) => negative_inputs_12_22_port, 
                           shift_in(21) => negative_inputs_12_21_port, 
                           shift_in(20) => negative_inputs_12_20_port, 
                           shift_in(19) => negative_inputs_12_19_port, 
                           shift_in(18) => negative_inputs_12_18_port, 
                           shift_in(17) => negative_inputs_12_17_port, 
                           shift_in(16) => negative_inputs_12_16_port, 
                           shift_in(15) => negative_inputs_12_15_port, 
                           shift_in(14) => negative_inputs_12_14_port, 
                           shift_in(13) => negative_inputs_12_13_port, 
                           shift_in(12) => negative_inputs_12_12_port, 
                           shift_in(11) => negative_inputs_12_11_port, 
                           shift_in(10) => negative_inputs_12_10_port, 
                           shift_in(9) => negative_inputs_12_9_port, 
                           shift_in(8) => negative_inputs_12_8_port, 
                           shift_in(7) => negative_inputs_12_7_port, 
                           shift_in(6) => negative_inputs_12_6_port, 
                           shift_in(5) => negative_inputs_12_5_port, 
                           shift_in(4) => negative_inputs_12_4_port, 
                           shift_in(3) => negative_inputs_12_3_port, 
                           shift_in(2) => negative_inputs_12_2_port, 
                           shift_in(1) => negative_inputs_12_1_port, 
                           shift_in(0) => n8, shift_out(63) => 
                           negative_inputs_13_63_port, shift_out(62) => 
                           negative_inputs_13_62_port, shift_out(61) => 
                           negative_inputs_13_61_port, shift_out(60) => 
                           negative_inputs_13_60_port, shift_out(59) => 
                           negative_inputs_13_59_port, shift_out(58) => 
                           negative_inputs_13_58_port, shift_out(57) => 
                           negative_inputs_13_57_port, shift_out(56) => 
                           negative_inputs_13_56_port, shift_out(55) => 
                           negative_inputs_13_55_port, shift_out(54) => 
                           negative_inputs_13_54_port, shift_out(53) => 
                           negative_inputs_13_53_port, shift_out(52) => 
                           negative_inputs_13_52_port, shift_out(51) => 
                           negative_inputs_13_51_port, shift_out(50) => 
                           negative_inputs_13_50_port, shift_out(49) => 
                           negative_inputs_13_49_port, shift_out(48) => 
                           negative_inputs_13_48_port, shift_out(47) => 
                           negative_inputs_13_47_port, shift_out(46) => 
                           negative_inputs_13_46_port, shift_out(45) => 
                           negative_inputs_13_45_port, shift_out(44) => 
                           negative_inputs_13_44_port, shift_out(43) => 
                           negative_inputs_13_43_port, shift_out(42) => 
                           negative_inputs_13_42_port, shift_out(41) => 
                           negative_inputs_13_41_port, shift_out(40) => 
                           negative_inputs_13_40_port, shift_out(39) => 
                           negative_inputs_13_39_port, shift_out(38) => 
                           negative_inputs_13_38_port, shift_out(37) => 
                           negative_inputs_13_37_port, shift_out(36) => 
                           negative_inputs_13_36_port, shift_out(35) => 
                           negative_inputs_13_35_port, shift_out(34) => 
                           negative_inputs_13_34_port, shift_out(33) => 
                           negative_inputs_13_33_port, shift_out(32) => 
                           negative_inputs_13_32_port, shift_out(31) => 
                           negative_inputs_13_31_port, shift_out(30) => 
                           negative_inputs_13_30_port, shift_out(29) => 
                           negative_inputs_13_29_port, shift_out(28) => 
                           negative_inputs_13_28_port, shift_out(27) => 
                           negative_inputs_13_27_port, shift_out(26) => 
                           negative_inputs_13_26_port, shift_out(25) => 
                           negative_inputs_13_25_port, shift_out(24) => 
                           negative_inputs_13_24_port, shift_out(23) => 
                           negative_inputs_13_23_port, shift_out(22) => 
                           negative_inputs_13_22_port, shift_out(21) => 
                           negative_inputs_13_21_port, shift_out(20) => 
                           negative_inputs_13_20_port, shift_out(19) => 
                           negative_inputs_13_19_port, shift_out(18) => 
                           negative_inputs_13_18_port, shift_out(17) => 
                           negative_inputs_13_17_port, shift_out(16) => 
                           negative_inputs_13_16_port, shift_out(15) => 
                           negative_inputs_13_15_port, shift_out(14) => 
                           negative_inputs_13_14_port, shift_out(13) => 
                           negative_inputs_13_13_port, shift_out(12) => 
                           negative_inputs_13_12_port, shift_out(11) => 
                           negative_inputs_13_11_port, shift_out(10) => 
                           negative_inputs_13_10_port, shift_out(9) => 
                           negative_inputs_13_9_port, shift_out(8) => 
                           negative_inputs_13_8_port, shift_out(7) => 
                           negative_inputs_13_7_port, shift_out(6) => 
                           negative_inputs_13_6_port, shift_out(5) => 
                           negative_inputs_13_5_port, shift_out(4) => 
                           negative_inputs_13_4_port, shift_out(3) => 
                           negative_inputs_13_3_port, shift_out(2) => 
                           negative_inputs_13_2_port, shift_out(1) => 
                           negative_inputs_13_1_port, shift_out(0) => n_1108);
   shifted_neg_14 : leftshifter_NbitShifter64_81 port map( shift_in(63) => 
                           negative_inputs_13_63_port, shift_in(62) => 
                           negative_inputs_13_62_port, shift_in(61) => 
                           negative_inputs_13_61_port, shift_in(60) => 
                           negative_inputs_13_60_port, shift_in(59) => 
                           negative_inputs_13_59_port, shift_in(58) => 
                           negative_inputs_13_58_port, shift_in(57) => 
                           negative_inputs_13_57_port, shift_in(56) => 
                           negative_inputs_13_56_port, shift_in(55) => 
                           negative_inputs_13_55_port, shift_in(54) => 
                           negative_inputs_13_54_port, shift_in(53) => 
                           negative_inputs_13_53_port, shift_in(52) => 
                           negative_inputs_13_52_port, shift_in(51) => 
                           negative_inputs_13_51_port, shift_in(50) => 
                           negative_inputs_13_50_port, shift_in(49) => 
                           negative_inputs_13_49_port, shift_in(48) => 
                           negative_inputs_13_48_port, shift_in(47) => n111, 
                           shift_in(46) => negative_inputs_13_46_port, 
                           shift_in(45) => negative_inputs_13_45_port, 
                           shift_in(44) => negative_inputs_13_44_port, 
                           shift_in(43) => negative_inputs_13_43_port, 
                           shift_in(42) => negative_inputs_13_42_port, 
                           shift_in(41) => negative_inputs_13_41_port, 
                           shift_in(40) => negative_inputs_13_40_port, 
                           shift_in(39) => negative_inputs_13_39_port, 
                           shift_in(38) => negative_inputs_13_38_port, 
                           shift_in(37) => negative_inputs_13_37_port, 
                           shift_in(36) => negative_inputs_13_36_port, 
                           shift_in(35) => negative_inputs_13_35_port, 
                           shift_in(34) => negative_inputs_13_34_port, 
                           shift_in(33) => negative_inputs_13_33_port, 
                           shift_in(32) => negative_inputs_13_32_port, 
                           shift_in(31) => negative_inputs_13_31_port, 
                           shift_in(30) => negative_inputs_13_30_port, 
                           shift_in(29) => negative_inputs_13_29_port, 
                           shift_in(28) => negative_inputs_13_28_port, 
                           shift_in(27) => negative_inputs_13_27_port, 
                           shift_in(26) => negative_inputs_13_26_port, 
                           shift_in(25) => negative_inputs_13_25_port, 
                           shift_in(24) => negative_inputs_13_24_port, 
                           shift_in(23) => negative_inputs_13_23_port, 
                           shift_in(22) => negative_inputs_13_22_port, 
                           shift_in(21) => negative_inputs_13_21_port, 
                           shift_in(20) => negative_inputs_13_20_port, 
                           shift_in(19) => negative_inputs_13_19_port, 
                           shift_in(18) => negative_inputs_13_18_port, 
                           shift_in(17) => negative_inputs_13_17_port, 
                           shift_in(16) => negative_inputs_13_16_port, 
                           shift_in(15) => negative_inputs_13_15_port, 
                           shift_in(14) => negative_inputs_13_14_port, 
                           shift_in(13) => negative_inputs_13_13_port, 
                           shift_in(12) => negative_inputs_13_12_port, 
                           shift_in(11) => negative_inputs_13_11_port, 
                           shift_in(10) => negative_inputs_13_10_port, 
                           shift_in(9) => negative_inputs_13_9_port, 
                           shift_in(8) => negative_inputs_13_8_port, 
                           shift_in(7) => negative_inputs_13_7_port, 
                           shift_in(6) => negative_inputs_13_6_port, 
                           shift_in(5) => negative_inputs_13_5_port, 
                           shift_in(4) => negative_inputs_13_4_port, 
                           shift_in(3) => negative_inputs_13_3_port, 
                           shift_in(2) => negative_inputs_13_2_port, 
                           shift_in(1) => negative_inputs_13_1_port, 
                           shift_in(0) => n8, shift_out(63) => 
                           negative_inputs_14_63_port, shift_out(62) => 
                           negative_inputs_14_62_port, shift_out(61) => 
                           negative_inputs_14_61_port, shift_out(60) => 
                           negative_inputs_14_60_port, shift_out(59) => 
                           negative_inputs_14_59_port, shift_out(58) => 
                           negative_inputs_14_58_port, shift_out(57) => 
                           negative_inputs_14_57_port, shift_out(56) => 
                           negative_inputs_14_56_port, shift_out(55) => 
                           negative_inputs_14_55_port, shift_out(54) => 
                           negative_inputs_14_54_port, shift_out(53) => 
                           negative_inputs_14_53_port, shift_out(52) => 
                           negative_inputs_14_52_port, shift_out(51) => 
                           negative_inputs_14_51_port, shift_out(50) => 
                           negative_inputs_14_50_port, shift_out(49) => 
                           negative_inputs_14_49_port, shift_out(48) => 
                           negative_inputs_14_48_port, shift_out(47) => 
                           negative_inputs_14_47_port, shift_out(46) => 
                           negative_inputs_14_46_port, shift_out(45) => 
                           negative_inputs_14_45_port, shift_out(44) => 
                           negative_inputs_14_44_port, shift_out(43) => 
                           negative_inputs_14_43_port, shift_out(42) => 
                           negative_inputs_14_42_port, shift_out(41) => 
                           negative_inputs_14_41_port, shift_out(40) => 
                           negative_inputs_14_40_port, shift_out(39) => 
                           negative_inputs_14_39_port, shift_out(38) => 
                           negative_inputs_14_38_port, shift_out(37) => 
                           negative_inputs_14_37_port, shift_out(36) => 
                           negative_inputs_14_36_port, shift_out(35) => 
                           negative_inputs_14_35_port, shift_out(34) => 
                           negative_inputs_14_34_port, shift_out(33) => 
                           negative_inputs_14_33_port, shift_out(32) => 
                           negative_inputs_14_32_port, shift_out(31) => 
                           negative_inputs_14_31_port, shift_out(30) => 
                           negative_inputs_14_30_port, shift_out(29) => 
                           negative_inputs_14_29_port, shift_out(28) => 
                           negative_inputs_14_28_port, shift_out(27) => 
                           negative_inputs_14_27_port, shift_out(26) => 
                           negative_inputs_14_26_port, shift_out(25) => 
                           negative_inputs_14_25_port, shift_out(24) => 
                           negative_inputs_14_24_port, shift_out(23) => 
                           negative_inputs_14_23_port, shift_out(22) => 
                           negative_inputs_14_22_port, shift_out(21) => 
                           negative_inputs_14_21_port, shift_out(20) => 
                           negative_inputs_14_20_port, shift_out(19) => 
                           negative_inputs_14_19_port, shift_out(18) => 
                           negative_inputs_14_18_port, shift_out(17) => 
                           negative_inputs_14_17_port, shift_out(16) => 
                           negative_inputs_14_16_port, shift_out(15) => 
                           negative_inputs_14_15_port, shift_out(14) => 
                           negative_inputs_14_14_port, shift_out(13) => 
                           negative_inputs_14_13_port, shift_out(12) => 
                           negative_inputs_14_12_port, shift_out(11) => 
                           negative_inputs_14_11_port, shift_out(10) => 
                           negative_inputs_14_10_port, shift_out(9) => 
                           negative_inputs_14_9_port, shift_out(8) => 
                           negative_inputs_14_8_port, shift_out(7) => 
                           negative_inputs_14_7_port, shift_out(6) => 
                           negative_inputs_14_6_port, shift_out(5) => 
                           negative_inputs_14_5_port, shift_out(4) => 
                           negative_inputs_14_4_port, shift_out(3) => 
                           negative_inputs_14_3_port, shift_out(2) => 
                           negative_inputs_14_2_port, shift_out(1) => 
                           negative_inputs_14_1_port, shift_out(0) => n_1109);
   shifted_neg_15 : leftshifter_NbitShifter64_80 port map( shift_in(63) => 
                           negative_inputs_14_63_port, shift_in(62) => 
                           negative_inputs_14_62_port, shift_in(61) => 
                           negative_inputs_14_61_port, shift_in(60) => 
                           negative_inputs_14_60_port, shift_in(59) => 
                           negative_inputs_14_59_port, shift_in(58) => 
                           negative_inputs_14_58_port, shift_in(57) => 
                           negative_inputs_14_57_port, shift_in(56) => 
                           negative_inputs_14_56_port, shift_in(55) => 
                           negative_inputs_14_55_port, shift_in(54) => 
                           negative_inputs_14_54_port, shift_in(53) => 
                           negative_inputs_14_53_port, shift_in(52) => 
                           negative_inputs_14_52_port, shift_in(51) => 
                           negative_inputs_14_51_port, shift_in(50) => 
                           negative_inputs_14_50_port, shift_in(49) => 
                           negative_inputs_14_49_port, shift_in(48) => 
                           negative_inputs_14_48_port, shift_in(47) => n109, 
                           shift_in(46) => negative_inputs_14_46_port, 
                           shift_in(45) => negative_inputs_14_45_port, 
                           shift_in(44) => negative_inputs_14_44_port, 
                           shift_in(43) => negative_inputs_14_43_port, 
                           shift_in(42) => negative_inputs_14_42_port, 
                           shift_in(41) => negative_inputs_14_41_port, 
                           shift_in(40) => negative_inputs_14_40_port, 
                           shift_in(39) => negative_inputs_14_39_port, 
                           shift_in(38) => negative_inputs_14_38_port, 
                           shift_in(37) => negative_inputs_14_37_port, 
                           shift_in(36) => negative_inputs_14_36_port, 
                           shift_in(35) => negative_inputs_14_35_port, 
                           shift_in(34) => negative_inputs_14_34_port, 
                           shift_in(33) => negative_inputs_14_33_port, 
                           shift_in(32) => negative_inputs_14_32_port, 
                           shift_in(31) => negative_inputs_14_31_port, 
                           shift_in(30) => negative_inputs_14_30_port, 
                           shift_in(29) => negative_inputs_14_29_port, 
                           shift_in(28) => negative_inputs_14_28_port, 
                           shift_in(27) => negative_inputs_14_27_port, 
                           shift_in(26) => negative_inputs_14_26_port, 
                           shift_in(25) => negative_inputs_14_25_port, 
                           shift_in(24) => negative_inputs_14_24_port, 
                           shift_in(23) => negative_inputs_14_23_port, 
                           shift_in(22) => negative_inputs_14_22_port, 
                           shift_in(21) => negative_inputs_14_21_port, 
                           shift_in(20) => negative_inputs_14_20_port, 
                           shift_in(19) => negative_inputs_14_19_port, 
                           shift_in(18) => negative_inputs_14_18_port, 
                           shift_in(17) => negative_inputs_14_17_port, 
                           shift_in(16) => negative_inputs_14_16_port, 
                           shift_in(15) => negative_inputs_14_15_port, 
                           shift_in(14) => negative_inputs_14_14_port, 
                           shift_in(13) => negative_inputs_14_13_port, 
                           shift_in(12) => negative_inputs_14_12_port, 
                           shift_in(11) => negative_inputs_14_11_port, 
                           shift_in(10) => negative_inputs_14_10_port, 
                           shift_in(9) => negative_inputs_14_9_port, 
                           shift_in(8) => negative_inputs_14_8_port, 
                           shift_in(7) => negative_inputs_14_7_port, 
                           shift_in(6) => negative_inputs_14_6_port, 
                           shift_in(5) => negative_inputs_14_5_port, 
                           shift_in(4) => negative_inputs_14_4_port, 
                           shift_in(3) => negative_inputs_14_3_port, 
                           shift_in(2) => negative_inputs_14_2_port, 
                           shift_in(1) => negative_inputs_14_1_port, 
                           shift_in(0) => n8, shift_out(63) => 
                           negative_inputs_15_63_port, shift_out(62) => 
                           negative_inputs_15_62_port, shift_out(61) => 
                           negative_inputs_15_61_port, shift_out(60) => 
                           negative_inputs_15_60_port, shift_out(59) => 
                           negative_inputs_15_59_port, shift_out(58) => 
                           negative_inputs_15_58_port, shift_out(57) => 
                           negative_inputs_15_57_port, shift_out(56) => 
                           negative_inputs_15_56_port, shift_out(55) => 
                           negative_inputs_15_55_port, shift_out(54) => 
                           negative_inputs_15_54_port, shift_out(53) => 
                           negative_inputs_15_53_port, shift_out(52) => 
                           negative_inputs_15_52_port, shift_out(51) => 
                           negative_inputs_15_51_port, shift_out(50) => 
                           negative_inputs_15_50_port, shift_out(49) => 
                           negative_inputs_15_49_port, shift_out(48) => 
                           negative_inputs_15_48_port, shift_out(47) => 
                           negative_inputs_15_47_port, shift_out(46) => 
                           negative_inputs_15_46_port, shift_out(45) => 
                           negative_inputs_15_45_port, shift_out(44) => 
                           negative_inputs_15_44_port, shift_out(43) => 
                           negative_inputs_15_43_port, shift_out(42) => 
                           negative_inputs_15_42_port, shift_out(41) => 
                           negative_inputs_15_41_port, shift_out(40) => 
                           negative_inputs_15_40_port, shift_out(39) => 
                           negative_inputs_15_39_port, shift_out(38) => 
                           negative_inputs_15_38_port, shift_out(37) => 
                           negative_inputs_15_37_port, shift_out(36) => 
                           negative_inputs_15_36_port, shift_out(35) => 
                           negative_inputs_15_35_port, shift_out(34) => 
                           negative_inputs_15_34_port, shift_out(33) => 
                           negative_inputs_15_33_port, shift_out(32) => 
                           negative_inputs_15_32_port, shift_out(31) => 
                           negative_inputs_15_31_port, shift_out(30) => 
                           negative_inputs_15_30_port, shift_out(29) => 
                           negative_inputs_15_29_port, shift_out(28) => 
                           negative_inputs_15_28_port, shift_out(27) => 
                           negative_inputs_15_27_port, shift_out(26) => 
                           negative_inputs_15_26_port, shift_out(25) => 
                           negative_inputs_15_25_port, shift_out(24) => 
                           negative_inputs_15_24_port, shift_out(23) => 
                           negative_inputs_15_23_port, shift_out(22) => 
                           negative_inputs_15_22_port, shift_out(21) => 
                           negative_inputs_15_21_port, shift_out(20) => 
                           negative_inputs_15_20_port, shift_out(19) => 
                           negative_inputs_15_19_port, shift_out(18) => 
                           negative_inputs_15_18_port, shift_out(17) => 
                           negative_inputs_15_17_port, shift_out(16) => 
                           negative_inputs_15_16_port, shift_out(15) => 
                           negative_inputs_15_15_port, shift_out(14) => 
                           negative_inputs_15_14_port, shift_out(13) => 
                           negative_inputs_15_13_port, shift_out(12) => 
                           negative_inputs_15_12_port, shift_out(11) => 
                           negative_inputs_15_11_port, shift_out(10) => 
                           negative_inputs_15_10_port, shift_out(9) => 
                           negative_inputs_15_9_port, shift_out(8) => 
                           negative_inputs_15_8_port, shift_out(7) => 
                           negative_inputs_15_7_port, shift_out(6) => 
                           negative_inputs_15_6_port, shift_out(5) => 
                           negative_inputs_15_5_port, shift_out(4) => 
                           negative_inputs_15_4_port, shift_out(3) => 
                           negative_inputs_15_3_port, shift_out(2) => 
                           negative_inputs_15_2_port, shift_out(1) => 
                           negative_inputs_15_1_port, shift_out(0) => n_1110);
   shifted_neg_16 : leftshifter_NbitShifter64_79 port map( shift_in(63) => 
                           negative_inputs_15_63_port, shift_in(62) => 
                           negative_inputs_15_62_port, shift_in(61) => 
                           negative_inputs_15_61_port, shift_in(60) => 
                           negative_inputs_15_60_port, shift_in(59) => 
                           negative_inputs_15_59_port, shift_in(58) => 
                           negative_inputs_15_58_port, shift_in(57) => 
                           negative_inputs_15_57_port, shift_in(56) => 
                           negative_inputs_15_56_port, shift_in(55) => 
                           negative_inputs_15_55_port, shift_in(54) => 
                           negative_inputs_15_54_port, shift_in(53) => 
                           negative_inputs_15_53_port, shift_in(52) => 
                           negative_inputs_15_52_port, shift_in(51) => 
                           negative_inputs_15_51_port, shift_in(50) => 
                           negative_inputs_15_50_port, shift_in(49) => 
                           negative_inputs_15_49_port, shift_in(48) => 
                           negative_inputs_15_48_port, shift_in(47) => n107, 
                           shift_in(46) => n105, shift_in(45) => n103, 
                           shift_in(44) => n101, shift_in(43) => n99, 
                           shift_in(42) => n97, shift_in(41) => n95, 
                           shift_in(40) => n93, shift_in(39) => n91, 
                           shift_in(38) => n89, shift_in(37) => n87, 
                           shift_in(36) => n85, shift_in(35) => n83, 
                           shift_in(34) => n81, shift_in(33) => n79, 
                           shift_in(32) => n77, shift_in(31) => n75, 
                           shift_in(30) => n73, shift_in(29) => n71, 
                           shift_in(28) => n69, shift_in(27) => n67, 
                           shift_in(26) => n65, shift_in(25) => n63, 
                           shift_in(24) => n61, shift_in(23) => n59, 
                           shift_in(22) => n57, shift_in(21) => n55, 
                           shift_in(20) => n53, shift_in(19) => n51, 
                           shift_in(18) => n49, shift_in(17) => n47, 
                           shift_in(16) => n45, shift_in(15) => n43, 
                           shift_in(14) => negative_inputs_15_14_port, 
                           shift_in(13) => negative_inputs_15_13_port, 
                           shift_in(12) => negative_inputs_15_12_port, 
                           shift_in(11) => negative_inputs_15_11_port, 
                           shift_in(10) => negative_inputs_15_10_port, 
                           shift_in(9) => negative_inputs_15_9_port, 
                           shift_in(8) => negative_inputs_15_8_port, 
                           shift_in(7) => negative_inputs_15_7_port, 
                           shift_in(6) => negative_inputs_15_6_port, 
                           shift_in(5) => negative_inputs_15_5_port, 
                           shift_in(4) => negative_inputs_15_4_port, 
                           shift_in(3) => negative_inputs_15_3_port, 
                           shift_in(2) => negative_inputs_15_2_port, 
                           shift_in(1) => negative_inputs_15_1_port, 
                           shift_in(0) => n8, shift_out(63) => 
                           negative_inputs_16_63_port, shift_out(62) => 
                           negative_inputs_16_62_port, shift_out(61) => 
                           negative_inputs_16_61_port, shift_out(60) => 
                           negative_inputs_16_60_port, shift_out(59) => 
                           negative_inputs_16_59_port, shift_out(58) => 
                           negative_inputs_16_58_port, shift_out(57) => 
                           negative_inputs_16_57_port, shift_out(56) => 
                           negative_inputs_16_56_port, shift_out(55) => 
                           negative_inputs_16_55_port, shift_out(54) => 
                           negative_inputs_16_54_port, shift_out(53) => 
                           negative_inputs_16_53_port, shift_out(52) => 
                           negative_inputs_16_52_port, shift_out(51) => 
                           negative_inputs_16_51_port, shift_out(50) => 
                           negative_inputs_16_50_port, shift_out(49) => 
                           negative_inputs_16_49_port, shift_out(48) => 
                           negative_inputs_16_48_port, shift_out(47) => 
                           negative_inputs_16_47_port, shift_out(46) => 
                           negative_inputs_16_46_port, shift_out(45) => 
                           negative_inputs_16_45_port, shift_out(44) => 
                           negative_inputs_16_44_port, shift_out(43) => 
                           negative_inputs_16_43_port, shift_out(42) => 
                           negative_inputs_16_42_port, shift_out(41) => 
                           negative_inputs_16_41_port, shift_out(40) => 
                           negative_inputs_16_40_port, shift_out(39) => 
                           negative_inputs_16_39_port, shift_out(38) => 
                           negative_inputs_16_38_port, shift_out(37) => 
                           negative_inputs_16_37_port, shift_out(36) => 
                           negative_inputs_16_36_port, shift_out(35) => 
                           negative_inputs_16_35_port, shift_out(34) => 
                           negative_inputs_16_34_port, shift_out(33) => 
                           negative_inputs_16_33_port, shift_out(32) => 
                           negative_inputs_16_32_port, shift_out(31) => 
                           negative_inputs_16_31_port, shift_out(30) => 
                           negative_inputs_16_30_port, shift_out(29) => 
                           negative_inputs_16_29_port, shift_out(28) => 
                           negative_inputs_16_28_port, shift_out(27) => 
                           negative_inputs_16_27_port, shift_out(26) => 
                           negative_inputs_16_26_port, shift_out(25) => 
                           negative_inputs_16_25_port, shift_out(24) => 
                           negative_inputs_16_24_port, shift_out(23) => 
                           negative_inputs_16_23_port, shift_out(22) => 
                           negative_inputs_16_22_port, shift_out(21) => 
                           negative_inputs_16_21_port, shift_out(20) => 
                           negative_inputs_16_20_port, shift_out(19) => 
                           negative_inputs_16_19_port, shift_out(18) => 
                           negative_inputs_16_18_port, shift_out(17) => 
                           negative_inputs_16_17_port, shift_out(16) => 
                           negative_inputs_16_16_port, shift_out(15) => 
                           negative_inputs_16_15_port, shift_out(14) => 
                           negative_inputs_16_14_port, shift_out(13) => 
                           negative_inputs_16_13_port, shift_out(12) => 
                           negative_inputs_16_12_port, shift_out(11) => 
                           negative_inputs_16_11_port, shift_out(10) => 
                           negative_inputs_16_10_port, shift_out(9) => 
                           negative_inputs_16_9_port, shift_out(8) => 
                           negative_inputs_16_8_port, shift_out(7) => 
                           negative_inputs_16_7_port, shift_out(6) => 
                           negative_inputs_16_6_port, shift_out(5) => 
                           negative_inputs_16_5_port, shift_out(4) => 
                           negative_inputs_16_4_port, shift_out(3) => 
                           negative_inputs_16_3_port, shift_out(2) => 
                           negative_inputs_16_2_port, shift_out(1) => 
                           negative_inputs_16_1_port, shift_out(0) => n_1111);
   shifted_neg_17 : leftshifter_NbitShifter64_78 port map( shift_in(63) => 
                           negative_inputs_16_63_port, shift_in(62) => 
                           negative_inputs_16_62_port, shift_in(61) => 
                           negative_inputs_16_61_port, shift_in(60) => 
                           negative_inputs_16_60_port, shift_in(59) => 
                           negative_inputs_16_59_port, shift_in(58) => 
                           negative_inputs_16_58_port, shift_in(57) => 
                           negative_inputs_16_57_port, shift_in(56) => 
                           negative_inputs_16_56_port, shift_in(55) => 
                           negative_inputs_16_55_port, shift_in(54) => 
                           negative_inputs_16_54_port, shift_in(53) => 
                           negative_inputs_16_53_port, shift_in(52) => 
                           negative_inputs_16_52_port, shift_in(51) => 
                           negative_inputs_16_51_port, shift_in(50) => 
                           negative_inputs_16_50_port, shift_in(49) => 
                           negative_inputs_16_49_port, shift_in(48) => 
                           negative_inputs_16_48_port, shift_in(47) => 
                           negative_inputs_16_47_port, shift_in(46) => 
                           negative_inputs_16_46_port, shift_in(45) => 
                           negative_inputs_16_45_port, shift_in(44) => 
                           negative_inputs_16_44_port, shift_in(43) => 
                           negative_inputs_16_43_port, shift_in(42) => 
                           negative_inputs_16_42_port, shift_in(41) => 
                           negative_inputs_16_41_port, shift_in(40) => 
                           negative_inputs_16_40_port, shift_in(39) => 
                           negative_inputs_16_39_port, shift_in(38) => 
                           negative_inputs_16_38_port, shift_in(37) => 
                           negative_inputs_16_37_port, shift_in(36) => 
                           negative_inputs_16_36_port, shift_in(35) => 
                           negative_inputs_16_35_port, shift_in(34) => 
                           negative_inputs_16_34_port, shift_in(33) => 
                           negative_inputs_16_33_port, shift_in(32) => 
                           negative_inputs_16_32_port, shift_in(31) => 
                           negative_inputs_16_31_port, shift_in(30) => 
                           negative_inputs_16_30_port, shift_in(29) => 
                           negative_inputs_16_29_port, shift_in(28) => 
                           negative_inputs_16_28_port, shift_in(27) => 
                           negative_inputs_16_27_port, shift_in(26) => 
                           negative_inputs_16_26_port, shift_in(25) => 
                           negative_inputs_16_25_port, shift_in(24) => 
                           negative_inputs_16_24_port, shift_in(23) => 
                           negative_inputs_16_23_port, shift_in(22) => 
                           negative_inputs_16_22_port, shift_in(21) => 
                           negative_inputs_16_21_port, shift_in(20) => 
                           negative_inputs_16_20_port, shift_in(19) => 
                           negative_inputs_16_19_port, shift_in(18) => 
                           negative_inputs_16_18_port, shift_in(17) => 
                           negative_inputs_16_17_port, shift_in(16) => 
                           negative_inputs_16_16_port, shift_in(15) => 
                           negative_inputs_16_15_port, shift_in(14) => 
                           negative_inputs_16_14_port, shift_in(13) => 
                           negative_inputs_16_13_port, shift_in(12) => 
                           negative_inputs_16_12_port, shift_in(11) => 
                           negative_inputs_16_11_port, shift_in(10) => 
                           negative_inputs_16_10_port, shift_in(9) => 
                           negative_inputs_16_9_port, shift_in(8) => 
                           negative_inputs_16_8_port, shift_in(7) => 
                           negative_inputs_16_7_port, shift_in(6) => 
                           negative_inputs_16_6_port, shift_in(5) => 
                           negative_inputs_16_5_port, shift_in(4) => 
                           negative_inputs_16_4_port, shift_in(3) => 
                           negative_inputs_16_3_port, shift_in(2) => 
                           negative_inputs_16_2_port, shift_in(1) => 
                           negative_inputs_16_1_port, shift_in(0) => n8, 
                           shift_out(63) => negative_inputs_17_63_port, 
                           shift_out(62) => negative_inputs_17_62_port, 
                           shift_out(61) => negative_inputs_17_61_port, 
                           shift_out(60) => negative_inputs_17_60_port, 
                           shift_out(59) => negative_inputs_17_59_port, 
                           shift_out(58) => negative_inputs_17_58_port, 
                           shift_out(57) => negative_inputs_17_57_port, 
                           shift_out(56) => negative_inputs_17_56_port, 
                           shift_out(55) => negative_inputs_17_55_port, 
                           shift_out(54) => negative_inputs_17_54_port, 
                           shift_out(53) => negative_inputs_17_53_port, 
                           shift_out(52) => negative_inputs_17_52_port, 
                           shift_out(51) => negative_inputs_17_51_port, 
                           shift_out(50) => negative_inputs_17_50_port, 
                           shift_out(49) => negative_inputs_17_49_port, 
                           shift_out(48) => negative_inputs_17_48_port, 
                           shift_out(47) => negative_inputs_17_47_port, 
                           shift_out(46) => negative_inputs_17_46_port, 
                           shift_out(45) => negative_inputs_17_45_port, 
                           shift_out(44) => negative_inputs_17_44_port, 
                           shift_out(43) => negative_inputs_17_43_port, 
                           shift_out(42) => negative_inputs_17_42_port, 
                           shift_out(41) => negative_inputs_17_41_port, 
                           shift_out(40) => negative_inputs_17_40_port, 
                           shift_out(39) => negative_inputs_17_39_port, 
                           shift_out(38) => negative_inputs_17_38_port, 
                           shift_out(37) => negative_inputs_17_37_port, 
                           shift_out(36) => negative_inputs_17_36_port, 
                           shift_out(35) => negative_inputs_17_35_port, 
                           shift_out(34) => negative_inputs_17_34_port, 
                           shift_out(33) => negative_inputs_17_33_port, 
                           shift_out(32) => negative_inputs_17_32_port, 
                           shift_out(31) => negative_inputs_17_31_port, 
                           shift_out(30) => negative_inputs_17_30_port, 
                           shift_out(29) => negative_inputs_17_29_port, 
                           shift_out(28) => negative_inputs_17_28_port, 
                           shift_out(27) => negative_inputs_17_27_port, 
                           shift_out(26) => negative_inputs_17_26_port, 
                           shift_out(25) => negative_inputs_17_25_port, 
                           shift_out(24) => negative_inputs_17_24_port, 
                           shift_out(23) => negative_inputs_17_23_port, 
                           shift_out(22) => negative_inputs_17_22_port, 
                           shift_out(21) => negative_inputs_17_21_port, 
                           shift_out(20) => negative_inputs_17_20_port, 
                           shift_out(19) => negative_inputs_17_19_port, 
                           shift_out(18) => negative_inputs_17_18_port, 
                           shift_out(17) => negative_inputs_17_17_port, 
                           shift_out(16) => negative_inputs_17_16_port, 
                           shift_out(15) => negative_inputs_17_15_port, 
                           shift_out(14) => negative_inputs_17_14_port, 
                           shift_out(13) => negative_inputs_17_13_port, 
                           shift_out(12) => negative_inputs_17_12_port, 
                           shift_out(11) => negative_inputs_17_11_port, 
                           shift_out(10) => negative_inputs_17_10_port, 
                           shift_out(9) => negative_inputs_17_9_port, 
                           shift_out(8) => negative_inputs_17_8_port, 
                           shift_out(7) => negative_inputs_17_7_port, 
                           shift_out(6) => negative_inputs_17_6_port, 
                           shift_out(5) => negative_inputs_17_5_port, 
                           shift_out(4) => negative_inputs_17_4_port, 
                           shift_out(3) => negative_inputs_17_3_port, 
                           shift_out(2) => negative_inputs_17_2_port, 
                           shift_out(1) => negative_inputs_17_1_port, 
                           shift_out(0) => n_1112);
   shifted_neg_18 : leftshifter_NbitShifter64_77 port map( shift_in(63) => 
                           negative_inputs_17_63_port, shift_in(62) => 
                           negative_inputs_17_62_port, shift_in(61) => 
                           negative_inputs_17_61_port, shift_in(60) => 
                           negative_inputs_17_60_port, shift_in(59) => 
                           negative_inputs_17_59_port, shift_in(58) => 
                           negative_inputs_17_58_port, shift_in(57) => 
                           negative_inputs_17_57_port, shift_in(56) => 
                           negative_inputs_17_56_port, shift_in(55) => 
                           negative_inputs_17_55_port, shift_in(54) => 
                           negative_inputs_17_54_port, shift_in(53) => 
                           negative_inputs_17_53_port, shift_in(52) => 
                           negative_inputs_17_52_port, shift_in(51) => 
                           negative_inputs_17_51_port, shift_in(50) => 
                           negative_inputs_17_50_port, shift_in(49) => 
                           negative_inputs_17_49_port, shift_in(48) => 
                           negative_inputs_17_48_port, shift_in(47) => 
                           negative_inputs_17_47_port, shift_in(46) => 
                           negative_inputs_17_46_port, shift_in(45) => 
                           negative_inputs_17_45_port, shift_in(44) => 
                           negative_inputs_17_44_port, shift_in(43) => 
                           negative_inputs_17_43_port, shift_in(42) => 
                           negative_inputs_17_42_port, shift_in(41) => 
                           negative_inputs_17_41_port, shift_in(40) => 
                           negative_inputs_17_40_port, shift_in(39) => 
                           negative_inputs_17_39_port, shift_in(38) => 
                           negative_inputs_17_38_port, shift_in(37) => 
                           negative_inputs_17_37_port, shift_in(36) => 
                           negative_inputs_17_36_port, shift_in(35) => 
                           negative_inputs_17_35_port, shift_in(34) => 
                           negative_inputs_17_34_port, shift_in(33) => 
                           negative_inputs_17_33_port, shift_in(32) => 
                           negative_inputs_17_32_port, shift_in(31) => 
                           negative_inputs_17_31_port, shift_in(30) => 
                           negative_inputs_17_30_port, shift_in(29) => 
                           negative_inputs_17_29_port, shift_in(28) => 
                           negative_inputs_17_28_port, shift_in(27) => 
                           negative_inputs_17_27_port, shift_in(26) => 
                           negative_inputs_17_26_port, shift_in(25) => 
                           negative_inputs_17_25_port, shift_in(24) => 
                           negative_inputs_17_24_port, shift_in(23) => 
                           negative_inputs_17_23_port, shift_in(22) => 
                           negative_inputs_17_22_port, shift_in(21) => 
                           negative_inputs_17_21_port, shift_in(20) => 
                           negative_inputs_17_20_port, shift_in(19) => 
                           negative_inputs_17_19_port, shift_in(18) => 
                           negative_inputs_17_18_port, shift_in(17) => 
                           negative_inputs_17_17_port, shift_in(16) => 
                           negative_inputs_17_16_port, shift_in(15) => 
                           negative_inputs_17_15_port, shift_in(14) => 
                           negative_inputs_17_14_port, shift_in(13) => 
                           negative_inputs_17_13_port, shift_in(12) => 
                           negative_inputs_17_12_port, shift_in(11) => 
                           negative_inputs_17_11_port, shift_in(10) => 
                           negative_inputs_17_10_port, shift_in(9) => 
                           negative_inputs_17_9_port, shift_in(8) => 
                           negative_inputs_17_8_port, shift_in(7) => 
                           negative_inputs_17_7_port, shift_in(6) => 
                           negative_inputs_17_6_port, shift_in(5) => 
                           negative_inputs_17_5_port, shift_in(4) => 
                           negative_inputs_17_4_port, shift_in(3) => 
                           negative_inputs_17_3_port, shift_in(2) => 
                           negative_inputs_17_2_port, shift_in(1) => 
                           negative_inputs_17_1_port, shift_in(0) => n8, 
                           shift_out(63) => negative_inputs_18_63_port, 
                           shift_out(62) => negative_inputs_18_62_port, 
                           shift_out(61) => negative_inputs_18_61_port, 
                           shift_out(60) => negative_inputs_18_60_port, 
                           shift_out(59) => negative_inputs_18_59_port, 
                           shift_out(58) => negative_inputs_18_58_port, 
                           shift_out(57) => negative_inputs_18_57_port, 
                           shift_out(56) => negative_inputs_18_56_port, 
                           shift_out(55) => negative_inputs_18_55_port, 
                           shift_out(54) => negative_inputs_18_54_port, 
                           shift_out(53) => negative_inputs_18_53_port, 
                           shift_out(52) => negative_inputs_18_52_port, 
                           shift_out(51) => negative_inputs_18_51_port, 
                           shift_out(50) => negative_inputs_18_50_port, 
                           shift_out(49) => negative_inputs_18_49_port, 
                           shift_out(48) => negative_inputs_18_48_port, 
                           shift_out(47) => negative_inputs_18_47_port, 
                           shift_out(46) => negative_inputs_18_46_port, 
                           shift_out(45) => negative_inputs_18_45_port, 
                           shift_out(44) => negative_inputs_18_44_port, 
                           shift_out(43) => negative_inputs_18_43_port, 
                           shift_out(42) => negative_inputs_18_42_port, 
                           shift_out(41) => negative_inputs_18_41_port, 
                           shift_out(40) => negative_inputs_18_40_port, 
                           shift_out(39) => negative_inputs_18_39_port, 
                           shift_out(38) => negative_inputs_18_38_port, 
                           shift_out(37) => negative_inputs_18_37_port, 
                           shift_out(36) => negative_inputs_18_36_port, 
                           shift_out(35) => negative_inputs_18_35_port, 
                           shift_out(34) => negative_inputs_18_34_port, 
                           shift_out(33) => negative_inputs_18_33_port, 
                           shift_out(32) => negative_inputs_18_32_port, 
                           shift_out(31) => negative_inputs_18_31_port, 
                           shift_out(30) => negative_inputs_18_30_port, 
                           shift_out(29) => negative_inputs_18_29_port, 
                           shift_out(28) => negative_inputs_18_28_port, 
                           shift_out(27) => negative_inputs_18_27_port, 
                           shift_out(26) => negative_inputs_18_26_port, 
                           shift_out(25) => negative_inputs_18_25_port, 
                           shift_out(24) => negative_inputs_18_24_port, 
                           shift_out(23) => negative_inputs_18_23_port, 
                           shift_out(22) => negative_inputs_18_22_port, 
                           shift_out(21) => negative_inputs_18_21_port, 
                           shift_out(20) => negative_inputs_18_20_port, 
                           shift_out(19) => negative_inputs_18_19_port, 
                           shift_out(18) => negative_inputs_18_18_port, 
                           shift_out(17) => negative_inputs_18_17_port, 
                           shift_out(16) => negative_inputs_18_16_port, 
                           shift_out(15) => negative_inputs_18_15_port, 
                           shift_out(14) => negative_inputs_18_14_port, 
                           shift_out(13) => negative_inputs_18_13_port, 
                           shift_out(12) => negative_inputs_18_12_port, 
                           shift_out(11) => negative_inputs_18_11_port, 
                           shift_out(10) => negative_inputs_18_10_port, 
                           shift_out(9) => negative_inputs_18_9_port, 
                           shift_out(8) => negative_inputs_18_8_port, 
                           shift_out(7) => negative_inputs_18_7_port, 
                           shift_out(6) => negative_inputs_18_6_port, 
                           shift_out(5) => negative_inputs_18_5_port, 
                           shift_out(4) => negative_inputs_18_4_port, 
                           shift_out(3) => negative_inputs_18_3_port, 
                           shift_out(2) => negative_inputs_18_2_port, 
                           shift_out(1) => negative_inputs_18_1_port, 
                           shift_out(0) => n_1113);
   shifted_neg_19 : leftshifter_NbitShifter64_76 port map( shift_in(63) => 
                           negative_inputs_18_63_port, shift_in(62) => 
                           negative_inputs_18_62_port, shift_in(61) => 
                           negative_inputs_18_61_port, shift_in(60) => 
                           negative_inputs_18_60_port, shift_in(59) => 
                           negative_inputs_18_59_port, shift_in(58) => 
                           negative_inputs_18_58_port, shift_in(57) => 
                           negative_inputs_18_57_port, shift_in(56) => 
                           negative_inputs_18_56_port, shift_in(55) => 
                           negative_inputs_18_55_port, shift_in(54) => 
                           negative_inputs_18_54_port, shift_in(53) => 
                           negative_inputs_18_53_port, shift_in(52) => 
                           negative_inputs_18_52_port, shift_in(51) => 
                           negative_inputs_18_51_port, shift_in(50) => 
                           negative_inputs_18_50_port, shift_in(49) => 
                           negative_inputs_18_49_port, shift_in(48) => 
                           negative_inputs_18_48_port, shift_in(47) => 
                           negative_inputs_18_47_port, shift_in(46) => 
                           negative_inputs_18_46_port, shift_in(45) => 
                           negative_inputs_18_45_port, shift_in(44) => 
                           negative_inputs_18_44_port, shift_in(43) => 
                           negative_inputs_18_43_port, shift_in(42) => 
                           negative_inputs_18_42_port, shift_in(41) => 
                           negative_inputs_18_41_port, shift_in(40) => 
                           negative_inputs_18_40_port, shift_in(39) => 
                           negative_inputs_18_39_port, shift_in(38) => 
                           negative_inputs_18_38_port, shift_in(37) => 
                           negative_inputs_18_37_port, shift_in(36) => 
                           negative_inputs_18_36_port, shift_in(35) => 
                           negative_inputs_18_35_port, shift_in(34) => 
                           negative_inputs_18_34_port, shift_in(33) => 
                           negative_inputs_18_33_port, shift_in(32) => 
                           negative_inputs_18_32_port, shift_in(31) => 
                           negative_inputs_18_31_port, shift_in(30) => 
                           negative_inputs_18_30_port, shift_in(29) => 
                           negative_inputs_18_29_port, shift_in(28) => 
                           negative_inputs_18_28_port, shift_in(27) => 
                           negative_inputs_18_27_port, shift_in(26) => 
                           negative_inputs_18_26_port, shift_in(25) => 
                           negative_inputs_18_25_port, shift_in(24) => 
                           negative_inputs_18_24_port, shift_in(23) => 
                           negative_inputs_18_23_port, shift_in(22) => 
                           negative_inputs_18_22_port, shift_in(21) => 
                           negative_inputs_18_21_port, shift_in(20) => 
                           negative_inputs_18_20_port, shift_in(19) => 
                           negative_inputs_18_19_port, shift_in(18) => 
                           negative_inputs_18_18_port, shift_in(17) => 
                           negative_inputs_18_17_port, shift_in(16) => 
                           negative_inputs_18_16_port, shift_in(15) => 
                           negative_inputs_18_15_port, shift_in(14) => 
                           negative_inputs_18_14_port, shift_in(13) => 
                           negative_inputs_18_13_port, shift_in(12) => 
                           negative_inputs_18_12_port, shift_in(11) => 
                           negative_inputs_18_11_port, shift_in(10) => 
                           negative_inputs_18_10_port, shift_in(9) => 
                           negative_inputs_18_9_port, shift_in(8) => 
                           negative_inputs_18_8_port, shift_in(7) => 
                           negative_inputs_18_7_port, shift_in(6) => 
                           negative_inputs_18_6_port, shift_in(5) => 
                           negative_inputs_18_5_port, shift_in(4) => 
                           negative_inputs_18_4_port, shift_in(3) => 
                           negative_inputs_18_3_port, shift_in(2) => 
                           negative_inputs_18_2_port, shift_in(1) => 
                           negative_inputs_18_1_port, shift_in(0) => n8, 
                           shift_out(63) => negative_inputs_19_63_port, 
                           shift_out(62) => negative_inputs_19_62_port, 
                           shift_out(61) => negative_inputs_19_61_port, 
                           shift_out(60) => negative_inputs_19_60_port, 
                           shift_out(59) => negative_inputs_19_59_port, 
                           shift_out(58) => negative_inputs_19_58_port, 
                           shift_out(57) => negative_inputs_19_57_port, 
                           shift_out(56) => negative_inputs_19_56_port, 
                           shift_out(55) => negative_inputs_19_55_port, 
                           shift_out(54) => negative_inputs_19_54_port, 
                           shift_out(53) => negative_inputs_19_53_port, 
                           shift_out(52) => negative_inputs_19_52_port, 
                           shift_out(51) => negative_inputs_19_51_port, 
                           shift_out(50) => negative_inputs_19_50_port, 
                           shift_out(49) => negative_inputs_19_49_port, 
                           shift_out(48) => negative_inputs_19_48_port, 
                           shift_out(47) => negative_inputs_19_47_port, 
                           shift_out(46) => negative_inputs_19_46_port, 
                           shift_out(45) => negative_inputs_19_45_port, 
                           shift_out(44) => negative_inputs_19_44_port, 
                           shift_out(43) => negative_inputs_19_43_port, 
                           shift_out(42) => negative_inputs_19_42_port, 
                           shift_out(41) => negative_inputs_19_41_port, 
                           shift_out(40) => negative_inputs_19_40_port, 
                           shift_out(39) => negative_inputs_19_39_port, 
                           shift_out(38) => negative_inputs_19_38_port, 
                           shift_out(37) => negative_inputs_19_37_port, 
                           shift_out(36) => negative_inputs_19_36_port, 
                           shift_out(35) => negative_inputs_19_35_port, 
                           shift_out(34) => negative_inputs_19_34_port, 
                           shift_out(33) => negative_inputs_19_33_port, 
                           shift_out(32) => negative_inputs_19_32_port, 
                           shift_out(31) => negative_inputs_19_31_port, 
                           shift_out(30) => negative_inputs_19_30_port, 
                           shift_out(29) => negative_inputs_19_29_port, 
                           shift_out(28) => negative_inputs_19_28_port, 
                           shift_out(27) => negative_inputs_19_27_port, 
                           shift_out(26) => negative_inputs_19_26_port, 
                           shift_out(25) => negative_inputs_19_25_port, 
                           shift_out(24) => negative_inputs_19_24_port, 
                           shift_out(23) => negative_inputs_19_23_port, 
                           shift_out(22) => negative_inputs_19_22_port, 
                           shift_out(21) => negative_inputs_19_21_port, 
                           shift_out(20) => negative_inputs_19_20_port, 
                           shift_out(19) => negative_inputs_19_19_port, 
                           shift_out(18) => negative_inputs_19_18_port, 
                           shift_out(17) => negative_inputs_19_17_port, 
                           shift_out(16) => negative_inputs_19_16_port, 
                           shift_out(15) => negative_inputs_19_15_port, 
                           shift_out(14) => negative_inputs_19_14_port, 
                           shift_out(13) => negative_inputs_19_13_port, 
                           shift_out(12) => negative_inputs_19_12_port, 
                           shift_out(11) => negative_inputs_19_11_port, 
                           shift_out(10) => negative_inputs_19_10_port, 
                           shift_out(9) => negative_inputs_19_9_port, 
                           shift_out(8) => negative_inputs_19_8_port, 
                           shift_out(7) => negative_inputs_19_7_port, 
                           shift_out(6) => negative_inputs_19_6_port, 
                           shift_out(5) => negative_inputs_19_5_port, 
                           shift_out(4) => negative_inputs_19_4_port, 
                           shift_out(3) => negative_inputs_19_3_port, 
                           shift_out(2) => negative_inputs_19_2_port, 
                           shift_out(1) => negative_inputs_19_1_port, 
                           shift_out(0) => n_1114);
   shifted_neg_20 : leftshifter_NbitShifter64_75 port map( shift_in(63) => 
                           negative_inputs_19_63_port, shift_in(62) => 
                           negative_inputs_19_62_port, shift_in(61) => 
                           negative_inputs_19_61_port, shift_in(60) => 
                           negative_inputs_19_60_port, shift_in(59) => 
                           negative_inputs_19_59_port, shift_in(58) => 
                           negative_inputs_19_58_port, shift_in(57) => 
                           negative_inputs_19_57_port, shift_in(56) => 
                           negative_inputs_19_56_port, shift_in(55) => 
                           negative_inputs_19_55_port, shift_in(54) => 
                           negative_inputs_19_54_port, shift_in(53) => 
                           negative_inputs_19_53_port, shift_in(52) => 
                           negative_inputs_19_52_port, shift_in(51) => 
                           negative_inputs_19_51_port, shift_in(50) => 
                           negative_inputs_19_50_port, shift_in(49) => 
                           negative_inputs_19_49_port, shift_in(48) => 
                           negative_inputs_19_48_port, shift_in(47) => 
                           negative_inputs_19_47_port, shift_in(46) => 
                           negative_inputs_19_46_port, shift_in(45) => 
                           negative_inputs_19_45_port, shift_in(44) => 
                           negative_inputs_19_44_port, shift_in(43) => 
                           negative_inputs_19_43_port, shift_in(42) => 
                           negative_inputs_19_42_port, shift_in(41) => 
                           negative_inputs_19_41_port, shift_in(40) => 
                           negative_inputs_19_40_port, shift_in(39) => 
                           negative_inputs_19_39_port, shift_in(38) => 
                           negative_inputs_19_38_port, shift_in(37) => 
                           negative_inputs_19_37_port, shift_in(36) => 
                           negative_inputs_19_36_port, shift_in(35) => 
                           negative_inputs_19_35_port, shift_in(34) => 
                           negative_inputs_19_34_port, shift_in(33) => 
                           negative_inputs_19_33_port, shift_in(32) => 
                           negative_inputs_19_32_port, shift_in(31) => 
                           negative_inputs_19_31_port, shift_in(30) => 
                           negative_inputs_19_30_port, shift_in(29) => 
                           negative_inputs_19_29_port, shift_in(28) => 
                           negative_inputs_19_28_port, shift_in(27) => 
                           negative_inputs_19_27_port, shift_in(26) => 
                           negative_inputs_19_26_port, shift_in(25) => 
                           negative_inputs_19_25_port, shift_in(24) => 
                           negative_inputs_19_24_port, shift_in(23) => 
                           negative_inputs_19_23_port, shift_in(22) => 
                           negative_inputs_19_22_port, shift_in(21) => 
                           negative_inputs_19_21_port, shift_in(20) => 
                           negative_inputs_19_20_port, shift_in(19) => 
                           negative_inputs_19_19_port, shift_in(18) => 
                           negative_inputs_19_18_port, shift_in(17) => 
                           negative_inputs_19_17_port, shift_in(16) => 
                           negative_inputs_19_16_port, shift_in(15) => 
                           negative_inputs_19_15_port, shift_in(14) => 
                           negative_inputs_19_14_port, shift_in(13) => 
                           negative_inputs_19_13_port, shift_in(12) => 
                           negative_inputs_19_12_port, shift_in(11) => 
                           negative_inputs_19_11_port, shift_in(10) => 
                           negative_inputs_19_10_port, shift_in(9) => 
                           negative_inputs_19_9_port, shift_in(8) => 
                           negative_inputs_19_8_port, shift_in(7) => 
                           negative_inputs_19_7_port, shift_in(6) => 
                           negative_inputs_19_6_port, shift_in(5) => 
                           negative_inputs_19_5_port, shift_in(4) => 
                           negative_inputs_19_4_port, shift_in(3) => 
                           negative_inputs_19_3_port, shift_in(2) => 
                           negative_inputs_19_2_port, shift_in(1) => 
                           negative_inputs_19_1_port, shift_in(0) => n8, 
                           shift_out(63) => negative_inputs_20_63_port, 
                           shift_out(62) => negative_inputs_20_62_port, 
                           shift_out(61) => negative_inputs_20_61_port, 
                           shift_out(60) => negative_inputs_20_60_port, 
                           shift_out(59) => negative_inputs_20_59_port, 
                           shift_out(58) => negative_inputs_20_58_port, 
                           shift_out(57) => negative_inputs_20_57_port, 
                           shift_out(56) => negative_inputs_20_56_port, 
                           shift_out(55) => negative_inputs_20_55_port, 
                           shift_out(54) => negative_inputs_20_54_port, 
                           shift_out(53) => negative_inputs_20_53_port, 
                           shift_out(52) => negative_inputs_20_52_port, 
                           shift_out(51) => negative_inputs_20_51_port, 
                           shift_out(50) => negative_inputs_20_50_port, 
                           shift_out(49) => negative_inputs_20_49_port, 
                           shift_out(48) => negative_inputs_20_48_port, 
                           shift_out(47) => negative_inputs_20_47_port, 
                           shift_out(46) => negative_inputs_20_46_port, 
                           shift_out(45) => negative_inputs_20_45_port, 
                           shift_out(44) => negative_inputs_20_44_port, 
                           shift_out(43) => negative_inputs_20_43_port, 
                           shift_out(42) => negative_inputs_20_42_port, 
                           shift_out(41) => negative_inputs_20_41_port, 
                           shift_out(40) => negative_inputs_20_40_port, 
                           shift_out(39) => negative_inputs_20_39_port, 
                           shift_out(38) => negative_inputs_20_38_port, 
                           shift_out(37) => negative_inputs_20_37_port, 
                           shift_out(36) => negative_inputs_20_36_port, 
                           shift_out(35) => negative_inputs_20_35_port, 
                           shift_out(34) => negative_inputs_20_34_port, 
                           shift_out(33) => negative_inputs_20_33_port, 
                           shift_out(32) => negative_inputs_20_32_port, 
                           shift_out(31) => negative_inputs_20_31_port, 
                           shift_out(30) => negative_inputs_20_30_port, 
                           shift_out(29) => negative_inputs_20_29_port, 
                           shift_out(28) => negative_inputs_20_28_port, 
                           shift_out(27) => negative_inputs_20_27_port, 
                           shift_out(26) => negative_inputs_20_26_port, 
                           shift_out(25) => negative_inputs_20_25_port, 
                           shift_out(24) => negative_inputs_20_24_port, 
                           shift_out(23) => negative_inputs_20_23_port, 
                           shift_out(22) => negative_inputs_20_22_port, 
                           shift_out(21) => negative_inputs_20_21_port, 
                           shift_out(20) => negative_inputs_20_20_port, 
                           shift_out(19) => negative_inputs_20_19_port, 
                           shift_out(18) => negative_inputs_20_18_port, 
                           shift_out(17) => negative_inputs_20_17_port, 
                           shift_out(16) => negative_inputs_20_16_port, 
                           shift_out(15) => negative_inputs_20_15_port, 
                           shift_out(14) => negative_inputs_20_14_port, 
                           shift_out(13) => negative_inputs_20_13_port, 
                           shift_out(12) => negative_inputs_20_12_port, 
                           shift_out(11) => negative_inputs_20_11_port, 
                           shift_out(10) => negative_inputs_20_10_port, 
                           shift_out(9) => negative_inputs_20_9_port, 
                           shift_out(8) => negative_inputs_20_8_port, 
                           shift_out(7) => negative_inputs_20_7_port, 
                           shift_out(6) => negative_inputs_20_6_port, 
                           shift_out(5) => negative_inputs_20_5_port, 
                           shift_out(4) => negative_inputs_20_4_port, 
                           shift_out(3) => negative_inputs_20_3_port, 
                           shift_out(2) => negative_inputs_20_2_port, 
                           shift_out(1) => negative_inputs_20_1_port, 
                           shift_out(0) => n_1115);
   shifted_neg_21 : leftshifter_NbitShifter64_74 port map( shift_in(63) => 
                           negative_inputs_20_63_port, shift_in(62) => 
                           negative_inputs_20_62_port, shift_in(61) => 
                           negative_inputs_20_61_port, shift_in(60) => 
                           negative_inputs_20_60_port, shift_in(59) => 
                           negative_inputs_20_59_port, shift_in(58) => 
                           negative_inputs_20_58_port, shift_in(57) => 
                           negative_inputs_20_57_port, shift_in(56) => 
                           negative_inputs_20_56_port, shift_in(55) => 
                           negative_inputs_20_55_port, shift_in(54) => 
                           negative_inputs_20_54_port, shift_in(53) => 
                           negative_inputs_20_53_port, shift_in(52) => 
                           negative_inputs_20_52_port, shift_in(51) => 
                           negative_inputs_20_51_port, shift_in(50) => 
                           negative_inputs_20_50_port, shift_in(49) => 
                           negative_inputs_20_49_port, shift_in(48) => 
                           negative_inputs_20_48_port, shift_in(47) => 
                           negative_inputs_20_47_port, shift_in(46) => 
                           negative_inputs_20_46_port, shift_in(45) => 
                           negative_inputs_20_45_port, shift_in(44) => 
                           negative_inputs_20_44_port, shift_in(43) => 
                           negative_inputs_20_43_port, shift_in(42) => 
                           negative_inputs_20_42_port, shift_in(41) => 
                           negative_inputs_20_41_port, shift_in(40) => 
                           negative_inputs_20_40_port, shift_in(39) => 
                           negative_inputs_20_39_port, shift_in(38) => 
                           negative_inputs_20_38_port, shift_in(37) => 
                           negative_inputs_20_37_port, shift_in(36) => 
                           negative_inputs_20_36_port, shift_in(35) => 
                           negative_inputs_20_35_port, shift_in(34) => 
                           negative_inputs_20_34_port, shift_in(33) => 
                           negative_inputs_20_33_port, shift_in(32) => 
                           negative_inputs_20_32_port, shift_in(31) => 
                           negative_inputs_20_31_port, shift_in(30) => 
                           negative_inputs_20_30_port, shift_in(29) => 
                           negative_inputs_20_29_port, shift_in(28) => 
                           negative_inputs_20_28_port, shift_in(27) => 
                           negative_inputs_20_27_port, shift_in(26) => 
                           negative_inputs_20_26_port, shift_in(25) => 
                           negative_inputs_20_25_port, shift_in(24) => 
                           negative_inputs_20_24_port, shift_in(23) => 
                           negative_inputs_20_23_port, shift_in(22) => 
                           negative_inputs_20_22_port, shift_in(21) => 
                           negative_inputs_20_21_port, shift_in(20) => 
                           negative_inputs_20_20_port, shift_in(19) => 
                           negative_inputs_20_19_port, shift_in(18) => 
                           negative_inputs_20_18_port, shift_in(17) => 
                           negative_inputs_20_17_port, shift_in(16) => 
                           negative_inputs_20_16_port, shift_in(15) => 
                           negative_inputs_20_15_port, shift_in(14) => 
                           negative_inputs_20_14_port, shift_in(13) => 
                           negative_inputs_20_13_port, shift_in(12) => 
                           negative_inputs_20_12_port, shift_in(11) => 
                           negative_inputs_20_11_port, shift_in(10) => 
                           negative_inputs_20_10_port, shift_in(9) => 
                           negative_inputs_20_9_port, shift_in(8) => 
                           negative_inputs_20_8_port, shift_in(7) => 
                           negative_inputs_20_7_port, shift_in(6) => 
                           negative_inputs_20_6_port, shift_in(5) => 
                           negative_inputs_20_5_port, shift_in(4) => 
                           negative_inputs_20_4_port, shift_in(3) => 
                           negative_inputs_20_3_port, shift_in(2) => 
                           negative_inputs_20_2_port, shift_in(1) => 
                           negative_inputs_20_1_port, shift_in(0) => n8, 
                           shift_out(63) => negative_inputs_21_63_port, 
                           shift_out(62) => negative_inputs_21_62_port, 
                           shift_out(61) => negative_inputs_21_61_port, 
                           shift_out(60) => negative_inputs_21_60_port, 
                           shift_out(59) => negative_inputs_21_59_port, 
                           shift_out(58) => negative_inputs_21_58_port, 
                           shift_out(57) => negative_inputs_21_57_port, 
                           shift_out(56) => negative_inputs_21_56_port, 
                           shift_out(55) => negative_inputs_21_55_port, 
                           shift_out(54) => negative_inputs_21_54_port, 
                           shift_out(53) => negative_inputs_21_53_port, 
                           shift_out(52) => negative_inputs_21_52_port, 
                           shift_out(51) => negative_inputs_21_51_port, 
                           shift_out(50) => negative_inputs_21_50_port, 
                           shift_out(49) => negative_inputs_21_49_port, 
                           shift_out(48) => negative_inputs_21_48_port, 
                           shift_out(47) => negative_inputs_21_47_port, 
                           shift_out(46) => negative_inputs_21_46_port, 
                           shift_out(45) => negative_inputs_21_45_port, 
                           shift_out(44) => negative_inputs_21_44_port, 
                           shift_out(43) => negative_inputs_21_43_port, 
                           shift_out(42) => negative_inputs_21_42_port, 
                           shift_out(41) => negative_inputs_21_41_port, 
                           shift_out(40) => negative_inputs_21_40_port, 
                           shift_out(39) => negative_inputs_21_39_port, 
                           shift_out(38) => negative_inputs_21_38_port, 
                           shift_out(37) => negative_inputs_21_37_port, 
                           shift_out(36) => negative_inputs_21_36_port, 
                           shift_out(35) => negative_inputs_21_35_port, 
                           shift_out(34) => negative_inputs_21_34_port, 
                           shift_out(33) => negative_inputs_21_33_port, 
                           shift_out(32) => negative_inputs_21_32_port, 
                           shift_out(31) => negative_inputs_21_31_port, 
                           shift_out(30) => negative_inputs_21_30_port, 
                           shift_out(29) => negative_inputs_21_29_port, 
                           shift_out(28) => negative_inputs_21_28_port, 
                           shift_out(27) => negative_inputs_21_27_port, 
                           shift_out(26) => negative_inputs_21_26_port, 
                           shift_out(25) => negative_inputs_21_25_port, 
                           shift_out(24) => negative_inputs_21_24_port, 
                           shift_out(23) => negative_inputs_21_23_port, 
                           shift_out(22) => negative_inputs_21_22_port, 
                           shift_out(21) => negative_inputs_21_21_port, 
                           shift_out(20) => negative_inputs_21_20_port, 
                           shift_out(19) => negative_inputs_21_19_port, 
                           shift_out(18) => negative_inputs_21_18_port, 
                           shift_out(17) => negative_inputs_21_17_port, 
                           shift_out(16) => negative_inputs_21_16_port, 
                           shift_out(15) => negative_inputs_21_15_port, 
                           shift_out(14) => negative_inputs_21_14_port, 
                           shift_out(13) => negative_inputs_21_13_port, 
                           shift_out(12) => negative_inputs_21_12_port, 
                           shift_out(11) => negative_inputs_21_11_port, 
                           shift_out(10) => negative_inputs_21_10_port, 
                           shift_out(9) => negative_inputs_21_9_port, 
                           shift_out(8) => negative_inputs_21_8_port, 
                           shift_out(7) => negative_inputs_21_7_port, 
                           shift_out(6) => negative_inputs_21_6_port, 
                           shift_out(5) => negative_inputs_21_5_port, 
                           shift_out(4) => negative_inputs_21_4_port, 
                           shift_out(3) => negative_inputs_21_3_port, 
                           shift_out(2) => negative_inputs_21_2_port, 
                           shift_out(1) => negative_inputs_21_1_port, 
                           shift_out(0) => n_1116);
   shifted_neg_22 : leftshifter_NbitShifter64_73 port map( shift_in(63) => 
                           negative_inputs_21_63_port, shift_in(62) => 
                           negative_inputs_21_62_port, shift_in(61) => 
                           negative_inputs_21_61_port, shift_in(60) => 
                           negative_inputs_21_60_port, shift_in(59) => 
                           negative_inputs_21_59_port, shift_in(58) => 
                           negative_inputs_21_58_port, shift_in(57) => 
                           negative_inputs_21_57_port, shift_in(56) => 
                           negative_inputs_21_56_port, shift_in(55) => 
                           negative_inputs_21_55_port, shift_in(54) => 
                           negative_inputs_21_54_port, shift_in(53) => 
                           negative_inputs_21_53_port, shift_in(52) => 
                           negative_inputs_21_52_port, shift_in(51) => 
                           negative_inputs_21_51_port, shift_in(50) => 
                           negative_inputs_21_50_port, shift_in(49) => 
                           negative_inputs_21_49_port, shift_in(48) => 
                           negative_inputs_21_48_port, shift_in(47) => 
                           negative_inputs_21_47_port, shift_in(46) => 
                           negative_inputs_21_46_port, shift_in(45) => 
                           negative_inputs_21_45_port, shift_in(44) => 
                           negative_inputs_21_44_port, shift_in(43) => 
                           negative_inputs_21_43_port, shift_in(42) => 
                           negative_inputs_21_42_port, shift_in(41) => 
                           negative_inputs_21_41_port, shift_in(40) => 
                           negative_inputs_21_40_port, shift_in(39) => 
                           negative_inputs_21_39_port, shift_in(38) => 
                           negative_inputs_21_38_port, shift_in(37) => 
                           negative_inputs_21_37_port, shift_in(36) => 
                           negative_inputs_21_36_port, shift_in(35) => 
                           negative_inputs_21_35_port, shift_in(34) => 
                           negative_inputs_21_34_port, shift_in(33) => 
                           negative_inputs_21_33_port, shift_in(32) => 
                           negative_inputs_21_32_port, shift_in(31) => 
                           negative_inputs_21_31_port, shift_in(30) => 
                           negative_inputs_21_30_port, shift_in(29) => 
                           negative_inputs_21_29_port, shift_in(28) => 
                           negative_inputs_21_28_port, shift_in(27) => 
                           negative_inputs_21_27_port, shift_in(26) => 
                           negative_inputs_21_26_port, shift_in(25) => 
                           negative_inputs_21_25_port, shift_in(24) => 
                           negative_inputs_21_24_port, shift_in(23) => 
                           negative_inputs_21_23_port, shift_in(22) => 
                           negative_inputs_21_22_port, shift_in(21) => 
                           negative_inputs_21_21_port, shift_in(20) => 
                           negative_inputs_21_20_port, shift_in(19) => 
                           negative_inputs_21_19_port, shift_in(18) => 
                           negative_inputs_21_18_port, shift_in(17) => 
                           negative_inputs_21_17_port, shift_in(16) => 
                           negative_inputs_21_16_port, shift_in(15) => 
                           negative_inputs_21_15_port, shift_in(14) => 
                           negative_inputs_21_14_port, shift_in(13) => 
                           negative_inputs_21_13_port, shift_in(12) => 
                           negative_inputs_21_12_port, shift_in(11) => 
                           negative_inputs_21_11_port, shift_in(10) => 
                           negative_inputs_21_10_port, shift_in(9) => 
                           negative_inputs_21_9_port, shift_in(8) => 
                           negative_inputs_21_8_port, shift_in(7) => 
                           negative_inputs_21_7_port, shift_in(6) => 
                           negative_inputs_21_6_port, shift_in(5) => 
                           negative_inputs_21_5_port, shift_in(4) => 
                           negative_inputs_21_4_port, shift_in(3) => 
                           negative_inputs_21_3_port, shift_in(2) => 
                           negative_inputs_21_2_port, shift_in(1) => 
                           negative_inputs_21_1_port, shift_in(0) => n8, 
                           shift_out(63) => negative_inputs_22_63_port, 
                           shift_out(62) => negative_inputs_22_62_port, 
                           shift_out(61) => negative_inputs_22_61_port, 
                           shift_out(60) => negative_inputs_22_60_port, 
                           shift_out(59) => negative_inputs_22_59_port, 
                           shift_out(58) => negative_inputs_22_58_port, 
                           shift_out(57) => negative_inputs_22_57_port, 
                           shift_out(56) => negative_inputs_22_56_port, 
                           shift_out(55) => negative_inputs_22_55_port, 
                           shift_out(54) => negative_inputs_22_54_port, 
                           shift_out(53) => negative_inputs_22_53_port, 
                           shift_out(52) => negative_inputs_22_52_port, 
                           shift_out(51) => negative_inputs_22_51_port, 
                           shift_out(50) => negative_inputs_22_50_port, 
                           shift_out(49) => negative_inputs_22_49_port, 
                           shift_out(48) => negative_inputs_22_48_port, 
                           shift_out(47) => negative_inputs_22_47_port, 
                           shift_out(46) => negative_inputs_22_46_port, 
                           shift_out(45) => negative_inputs_22_45_port, 
                           shift_out(44) => negative_inputs_22_44_port, 
                           shift_out(43) => negative_inputs_22_43_port, 
                           shift_out(42) => negative_inputs_22_42_port, 
                           shift_out(41) => negative_inputs_22_41_port, 
                           shift_out(40) => negative_inputs_22_40_port, 
                           shift_out(39) => negative_inputs_22_39_port, 
                           shift_out(38) => negative_inputs_22_38_port, 
                           shift_out(37) => negative_inputs_22_37_port, 
                           shift_out(36) => negative_inputs_22_36_port, 
                           shift_out(35) => negative_inputs_22_35_port, 
                           shift_out(34) => negative_inputs_22_34_port, 
                           shift_out(33) => negative_inputs_22_33_port, 
                           shift_out(32) => negative_inputs_22_32_port, 
                           shift_out(31) => negative_inputs_22_31_port, 
                           shift_out(30) => negative_inputs_22_30_port, 
                           shift_out(29) => negative_inputs_22_29_port, 
                           shift_out(28) => negative_inputs_22_28_port, 
                           shift_out(27) => negative_inputs_22_27_port, 
                           shift_out(26) => negative_inputs_22_26_port, 
                           shift_out(25) => negative_inputs_22_25_port, 
                           shift_out(24) => negative_inputs_22_24_port, 
                           shift_out(23) => negative_inputs_22_23_port, 
                           shift_out(22) => negative_inputs_22_22_port, 
                           shift_out(21) => negative_inputs_22_21_port, 
                           shift_out(20) => negative_inputs_22_20_port, 
                           shift_out(19) => negative_inputs_22_19_port, 
                           shift_out(18) => negative_inputs_22_18_port, 
                           shift_out(17) => negative_inputs_22_17_port, 
                           shift_out(16) => negative_inputs_22_16_port, 
                           shift_out(15) => negative_inputs_22_15_port, 
                           shift_out(14) => negative_inputs_22_14_port, 
                           shift_out(13) => negative_inputs_22_13_port, 
                           shift_out(12) => negative_inputs_22_12_port, 
                           shift_out(11) => negative_inputs_22_11_port, 
                           shift_out(10) => negative_inputs_22_10_port, 
                           shift_out(9) => negative_inputs_22_9_port, 
                           shift_out(8) => negative_inputs_22_8_port, 
                           shift_out(7) => negative_inputs_22_7_port, 
                           shift_out(6) => negative_inputs_22_6_port, 
                           shift_out(5) => negative_inputs_22_5_port, 
                           shift_out(4) => negative_inputs_22_4_port, 
                           shift_out(3) => negative_inputs_22_3_port, 
                           shift_out(2) => negative_inputs_22_2_port, 
                           shift_out(1) => negative_inputs_22_1_port, 
                           shift_out(0) => n_1117);
   shifted_neg_23 : leftshifter_NbitShifter64_72 port map( shift_in(63) => 
                           negative_inputs_22_63_port, shift_in(62) => 
                           negative_inputs_22_62_port, shift_in(61) => 
                           negative_inputs_22_61_port, shift_in(60) => 
                           negative_inputs_22_60_port, shift_in(59) => 
                           negative_inputs_22_59_port, shift_in(58) => 
                           negative_inputs_22_58_port, shift_in(57) => 
                           negative_inputs_22_57_port, shift_in(56) => 
                           negative_inputs_22_56_port, shift_in(55) => 
                           negative_inputs_22_55_port, shift_in(54) => 
                           negative_inputs_22_54_port, shift_in(53) => 
                           negative_inputs_22_53_port, shift_in(52) => 
                           negative_inputs_22_52_port, shift_in(51) => 
                           negative_inputs_22_51_port, shift_in(50) => 
                           negative_inputs_22_50_port, shift_in(49) => 
                           negative_inputs_22_49_port, shift_in(48) => 
                           negative_inputs_22_48_port, shift_in(47) => 
                           negative_inputs_22_47_port, shift_in(46) => 
                           negative_inputs_22_46_port, shift_in(45) => 
                           negative_inputs_22_45_port, shift_in(44) => 
                           negative_inputs_22_44_port, shift_in(43) => 
                           negative_inputs_22_43_port, shift_in(42) => 
                           negative_inputs_22_42_port, shift_in(41) => 
                           negative_inputs_22_41_port, shift_in(40) => 
                           negative_inputs_22_40_port, shift_in(39) => 
                           negative_inputs_22_39_port, shift_in(38) => 
                           negative_inputs_22_38_port, shift_in(37) => 
                           negative_inputs_22_37_port, shift_in(36) => 
                           negative_inputs_22_36_port, shift_in(35) => 
                           negative_inputs_22_35_port, shift_in(34) => 
                           negative_inputs_22_34_port, shift_in(33) => 
                           negative_inputs_22_33_port, shift_in(32) => 
                           negative_inputs_22_32_port, shift_in(31) => 
                           negative_inputs_22_31_port, shift_in(30) => 
                           negative_inputs_22_30_port, shift_in(29) => 
                           negative_inputs_22_29_port, shift_in(28) => 
                           negative_inputs_22_28_port, shift_in(27) => 
                           negative_inputs_22_27_port, shift_in(26) => 
                           negative_inputs_22_26_port, shift_in(25) => 
                           negative_inputs_22_25_port, shift_in(24) => 
                           negative_inputs_22_24_port, shift_in(23) => 
                           negative_inputs_22_23_port, shift_in(22) => 
                           negative_inputs_22_22_port, shift_in(21) => 
                           negative_inputs_22_21_port, shift_in(20) => 
                           negative_inputs_22_20_port, shift_in(19) => 
                           negative_inputs_22_19_port, shift_in(18) => 
                           negative_inputs_22_18_port, shift_in(17) => 
                           negative_inputs_22_17_port, shift_in(16) => 
                           negative_inputs_22_16_port, shift_in(15) => 
                           negative_inputs_22_15_port, shift_in(14) => 
                           negative_inputs_22_14_port, shift_in(13) => 
                           negative_inputs_22_13_port, shift_in(12) => 
                           negative_inputs_22_12_port, shift_in(11) => 
                           negative_inputs_22_11_port, shift_in(10) => 
                           negative_inputs_22_10_port, shift_in(9) => 
                           negative_inputs_22_9_port, shift_in(8) => 
                           negative_inputs_22_8_port, shift_in(7) => 
                           negative_inputs_22_7_port, shift_in(6) => 
                           negative_inputs_22_6_port, shift_in(5) => 
                           negative_inputs_22_5_port, shift_in(4) => 
                           negative_inputs_22_4_port, shift_in(3) => 
                           negative_inputs_22_3_port, shift_in(2) => 
                           negative_inputs_22_2_port, shift_in(1) => 
                           negative_inputs_22_1_port, shift_in(0) => n8, 
                           shift_out(63) => negative_inputs_23_63_port, 
                           shift_out(62) => negative_inputs_23_62_port, 
                           shift_out(61) => negative_inputs_23_61_port, 
                           shift_out(60) => negative_inputs_23_60_port, 
                           shift_out(59) => negative_inputs_23_59_port, 
                           shift_out(58) => negative_inputs_23_58_port, 
                           shift_out(57) => negative_inputs_23_57_port, 
                           shift_out(56) => negative_inputs_23_56_port, 
                           shift_out(55) => negative_inputs_23_55_port, 
                           shift_out(54) => negative_inputs_23_54_port, 
                           shift_out(53) => negative_inputs_23_53_port, 
                           shift_out(52) => negative_inputs_23_52_port, 
                           shift_out(51) => negative_inputs_23_51_port, 
                           shift_out(50) => negative_inputs_23_50_port, 
                           shift_out(49) => negative_inputs_23_49_port, 
                           shift_out(48) => negative_inputs_23_48_port, 
                           shift_out(47) => negative_inputs_23_47_port, 
                           shift_out(46) => negative_inputs_23_46_port, 
                           shift_out(45) => negative_inputs_23_45_port, 
                           shift_out(44) => negative_inputs_23_44_port, 
                           shift_out(43) => negative_inputs_23_43_port, 
                           shift_out(42) => negative_inputs_23_42_port, 
                           shift_out(41) => negative_inputs_23_41_port, 
                           shift_out(40) => negative_inputs_23_40_port, 
                           shift_out(39) => negative_inputs_23_39_port, 
                           shift_out(38) => negative_inputs_23_38_port, 
                           shift_out(37) => negative_inputs_23_37_port, 
                           shift_out(36) => negative_inputs_23_36_port, 
                           shift_out(35) => negative_inputs_23_35_port, 
                           shift_out(34) => negative_inputs_23_34_port, 
                           shift_out(33) => negative_inputs_23_33_port, 
                           shift_out(32) => negative_inputs_23_32_port, 
                           shift_out(31) => negative_inputs_23_31_port, 
                           shift_out(30) => negative_inputs_23_30_port, 
                           shift_out(29) => negative_inputs_23_29_port, 
                           shift_out(28) => negative_inputs_23_28_port, 
                           shift_out(27) => negative_inputs_23_27_port, 
                           shift_out(26) => negative_inputs_23_26_port, 
                           shift_out(25) => negative_inputs_23_25_port, 
                           shift_out(24) => negative_inputs_23_24_port, 
                           shift_out(23) => negative_inputs_23_23_port, 
                           shift_out(22) => negative_inputs_23_22_port, 
                           shift_out(21) => negative_inputs_23_21_port, 
                           shift_out(20) => negative_inputs_23_20_port, 
                           shift_out(19) => negative_inputs_23_19_port, 
                           shift_out(18) => negative_inputs_23_18_port, 
                           shift_out(17) => negative_inputs_23_17_port, 
                           shift_out(16) => negative_inputs_23_16_port, 
                           shift_out(15) => negative_inputs_23_15_port, 
                           shift_out(14) => negative_inputs_23_14_port, 
                           shift_out(13) => negative_inputs_23_13_port, 
                           shift_out(12) => negative_inputs_23_12_port, 
                           shift_out(11) => negative_inputs_23_11_port, 
                           shift_out(10) => negative_inputs_23_10_port, 
                           shift_out(9) => negative_inputs_23_9_port, 
                           shift_out(8) => negative_inputs_23_8_port, 
                           shift_out(7) => negative_inputs_23_7_port, 
                           shift_out(6) => negative_inputs_23_6_port, 
                           shift_out(5) => negative_inputs_23_5_port, 
                           shift_out(4) => negative_inputs_23_4_port, 
                           shift_out(3) => negative_inputs_23_3_port, 
                           shift_out(2) => negative_inputs_23_2_port, 
                           shift_out(1) => negative_inputs_23_1_port, 
                           shift_out(0) => n_1118);
   shifted_neg_24 : leftshifter_NbitShifter64_71 port map( shift_in(63) => 
                           negative_inputs_23_63_port, shift_in(62) => 
                           negative_inputs_23_62_port, shift_in(61) => 
                           negative_inputs_23_61_port, shift_in(60) => 
                           negative_inputs_23_60_port, shift_in(59) => 
                           negative_inputs_23_59_port, shift_in(58) => 
                           negative_inputs_23_58_port, shift_in(57) => 
                           negative_inputs_23_57_port, shift_in(56) => 
                           negative_inputs_23_56_port, shift_in(55) => 
                           negative_inputs_23_55_port, shift_in(54) => 
                           negative_inputs_23_54_port, shift_in(53) => 
                           negative_inputs_23_53_port, shift_in(52) => 
                           negative_inputs_23_52_port, shift_in(51) => 
                           negative_inputs_23_51_port, shift_in(50) => 
                           negative_inputs_23_50_port, shift_in(49) => 
                           negative_inputs_23_49_port, shift_in(48) => 
                           negative_inputs_23_48_port, shift_in(47) => 
                           negative_inputs_23_47_port, shift_in(46) => 
                           negative_inputs_23_46_port, shift_in(45) => 
                           negative_inputs_23_45_port, shift_in(44) => 
                           negative_inputs_23_44_port, shift_in(43) => 
                           negative_inputs_23_43_port, shift_in(42) => 
                           negative_inputs_23_42_port, shift_in(41) => 
                           negative_inputs_23_41_port, shift_in(40) => 
                           negative_inputs_23_40_port, shift_in(39) => 
                           negative_inputs_23_39_port, shift_in(38) => 
                           negative_inputs_23_38_port, shift_in(37) => 
                           negative_inputs_23_37_port, shift_in(36) => 
                           negative_inputs_23_36_port, shift_in(35) => 
                           negative_inputs_23_35_port, shift_in(34) => 
                           negative_inputs_23_34_port, shift_in(33) => 
                           negative_inputs_23_33_port, shift_in(32) => 
                           negative_inputs_23_32_port, shift_in(31) => 
                           negative_inputs_23_31_port, shift_in(30) => 
                           negative_inputs_23_30_port, shift_in(29) => 
                           negative_inputs_23_29_port, shift_in(28) => 
                           negative_inputs_23_28_port, shift_in(27) => 
                           negative_inputs_23_27_port, shift_in(26) => 
                           negative_inputs_23_26_port, shift_in(25) => 
                           negative_inputs_23_25_port, shift_in(24) => 
                           negative_inputs_23_24_port, shift_in(23) => 
                           negative_inputs_23_23_port, shift_in(22) => 
                           negative_inputs_23_22_port, shift_in(21) => 
                           negative_inputs_23_21_port, shift_in(20) => 
                           negative_inputs_23_20_port, shift_in(19) => 
                           negative_inputs_23_19_port, shift_in(18) => 
                           negative_inputs_23_18_port, shift_in(17) => 
                           negative_inputs_23_17_port, shift_in(16) => 
                           negative_inputs_23_16_port, shift_in(15) => 
                           negative_inputs_23_15_port, shift_in(14) => 
                           negative_inputs_23_14_port, shift_in(13) => 
                           negative_inputs_23_13_port, shift_in(12) => 
                           negative_inputs_23_12_port, shift_in(11) => 
                           negative_inputs_23_11_port, shift_in(10) => 
                           negative_inputs_23_10_port, shift_in(9) => 
                           negative_inputs_23_9_port, shift_in(8) => 
                           negative_inputs_23_8_port, shift_in(7) => 
                           negative_inputs_23_7_port, shift_in(6) => 
                           negative_inputs_23_6_port, shift_in(5) => 
                           negative_inputs_23_5_port, shift_in(4) => 
                           negative_inputs_23_4_port, shift_in(3) => 
                           negative_inputs_23_3_port, shift_in(2) => 
                           negative_inputs_23_2_port, shift_in(1) => 
                           negative_inputs_23_1_port, shift_in(0) => n8, 
                           shift_out(63) => negative_inputs_24_63_port, 
                           shift_out(62) => negative_inputs_24_62_port, 
                           shift_out(61) => negative_inputs_24_61_port, 
                           shift_out(60) => negative_inputs_24_60_port, 
                           shift_out(59) => negative_inputs_24_59_port, 
                           shift_out(58) => negative_inputs_24_58_port, 
                           shift_out(57) => negative_inputs_24_57_port, 
                           shift_out(56) => negative_inputs_24_56_port, 
                           shift_out(55) => negative_inputs_24_55_port, 
                           shift_out(54) => negative_inputs_24_54_port, 
                           shift_out(53) => negative_inputs_24_53_port, 
                           shift_out(52) => negative_inputs_24_52_port, 
                           shift_out(51) => negative_inputs_24_51_port, 
                           shift_out(50) => negative_inputs_24_50_port, 
                           shift_out(49) => negative_inputs_24_49_port, 
                           shift_out(48) => negative_inputs_24_48_port, 
                           shift_out(47) => negative_inputs_24_47_port, 
                           shift_out(46) => negative_inputs_24_46_port, 
                           shift_out(45) => negative_inputs_24_45_port, 
                           shift_out(44) => negative_inputs_24_44_port, 
                           shift_out(43) => negative_inputs_24_43_port, 
                           shift_out(42) => negative_inputs_24_42_port, 
                           shift_out(41) => negative_inputs_24_41_port, 
                           shift_out(40) => negative_inputs_24_40_port, 
                           shift_out(39) => negative_inputs_24_39_port, 
                           shift_out(38) => negative_inputs_24_38_port, 
                           shift_out(37) => negative_inputs_24_37_port, 
                           shift_out(36) => negative_inputs_24_36_port, 
                           shift_out(35) => negative_inputs_24_35_port, 
                           shift_out(34) => negative_inputs_24_34_port, 
                           shift_out(33) => negative_inputs_24_33_port, 
                           shift_out(32) => negative_inputs_24_32_port, 
                           shift_out(31) => negative_inputs_24_31_port, 
                           shift_out(30) => negative_inputs_24_30_port, 
                           shift_out(29) => negative_inputs_24_29_port, 
                           shift_out(28) => negative_inputs_24_28_port, 
                           shift_out(27) => negative_inputs_24_27_port, 
                           shift_out(26) => negative_inputs_24_26_port, 
                           shift_out(25) => negative_inputs_24_25_port, 
                           shift_out(24) => negative_inputs_24_24_port, 
                           shift_out(23) => negative_inputs_24_23_port, 
                           shift_out(22) => negative_inputs_24_22_port, 
                           shift_out(21) => negative_inputs_24_21_port, 
                           shift_out(20) => negative_inputs_24_20_port, 
                           shift_out(19) => negative_inputs_24_19_port, 
                           shift_out(18) => negative_inputs_24_18_port, 
                           shift_out(17) => negative_inputs_24_17_port, 
                           shift_out(16) => negative_inputs_24_16_port, 
                           shift_out(15) => negative_inputs_24_15_port, 
                           shift_out(14) => negative_inputs_24_14_port, 
                           shift_out(13) => negative_inputs_24_13_port, 
                           shift_out(12) => negative_inputs_24_12_port, 
                           shift_out(11) => negative_inputs_24_11_port, 
                           shift_out(10) => negative_inputs_24_10_port, 
                           shift_out(9) => negative_inputs_24_9_port, 
                           shift_out(8) => negative_inputs_24_8_port, 
                           shift_out(7) => negative_inputs_24_7_port, 
                           shift_out(6) => negative_inputs_24_6_port, 
                           shift_out(5) => negative_inputs_24_5_port, 
                           shift_out(4) => negative_inputs_24_4_port, 
                           shift_out(3) => negative_inputs_24_3_port, 
                           shift_out(2) => negative_inputs_24_2_port, 
                           shift_out(1) => negative_inputs_24_1_port, 
                           shift_out(0) => n_1119);
   shifted_neg_25 : leftshifter_NbitShifter64_70 port map( shift_in(63) => 
                           negative_inputs_24_63_port, shift_in(62) => 
                           negative_inputs_24_62_port, shift_in(61) => 
                           negative_inputs_24_61_port, shift_in(60) => 
                           negative_inputs_24_60_port, shift_in(59) => 
                           negative_inputs_24_59_port, shift_in(58) => 
                           negative_inputs_24_58_port, shift_in(57) => 
                           negative_inputs_24_57_port, shift_in(56) => 
                           negative_inputs_24_56_port, shift_in(55) => 
                           negative_inputs_24_55_port, shift_in(54) => 
                           negative_inputs_24_54_port, shift_in(53) => 
                           negative_inputs_24_53_port, shift_in(52) => 
                           negative_inputs_24_52_port, shift_in(51) => 
                           negative_inputs_24_51_port, shift_in(50) => 
                           negative_inputs_24_50_port, shift_in(49) => 
                           negative_inputs_24_49_port, shift_in(48) => 
                           negative_inputs_24_48_port, shift_in(47) => 
                           negative_inputs_24_47_port, shift_in(46) => 
                           negative_inputs_24_46_port, shift_in(45) => 
                           negative_inputs_24_45_port, shift_in(44) => 
                           negative_inputs_24_44_port, shift_in(43) => 
                           negative_inputs_24_43_port, shift_in(42) => 
                           negative_inputs_24_42_port, shift_in(41) => 
                           negative_inputs_24_41_port, shift_in(40) => 
                           negative_inputs_24_40_port, shift_in(39) => 
                           negative_inputs_24_39_port, shift_in(38) => 
                           negative_inputs_24_38_port, shift_in(37) => 
                           negative_inputs_24_37_port, shift_in(36) => 
                           negative_inputs_24_36_port, shift_in(35) => 
                           negative_inputs_24_35_port, shift_in(34) => 
                           negative_inputs_24_34_port, shift_in(33) => 
                           negative_inputs_24_33_port, shift_in(32) => 
                           negative_inputs_24_32_port, shift_in(31) => 
                           negative_inputs_24_31_port, shift_in(30) => 
                           negative_inputs_24_30_port, shift_in(29) => 
                           negative_inputs_24_29_port, shift_in(28) => 
                           negative_inputs_24_28_port, shift_in(27) => 
                           negative_inputs_24_27_port, shift_in(26) => 
                           negative_inputs_24_26_port, shift_in(25) => 
                           negative_inputs_24_25_port, shift_in(24) => 
                           negative_inputs_24_24_port, shift_in(23) => 
                           negative_inputs_24_23_port, shift_in(22) => 
                           negative_inputs_24_22_port, shift_in(21) => 
                           negative_inputs_24_21_port, shift_in(20) => 
                           negative_inputs_24_20_port, shift_in(19) => 
                           negative_inputs_24_19_port, shift_in(18) => 
                           negative_inputs_24_18_port, shift_in(17) => 
                           negative_inputs_24_17_port, shift_in(16) => 
                           negative_inputs_24_16_port, shift_in(15) => 
                           negative_inputs_24_15_port, shift_in(14) => 
                           negative_inputs_24_14_port, shift_in(13) => 
                           negative_inputs_24_13_port, shift_in(12) => 
                           negative_inputs_24_12_port, shift_in(11) => 
                           negative_inputs_24_11_port, shift_in(10) => 
                           negative_inputs_24_10_port, shift_in(9) => 
                           negative_inputs_24_9_port, shift_in(8) => 
                           negative_inputs_24_8_port, shift_in(7) => 
                           negative_inputs_24_7_port, shift_in(6) => 
                           negative_inputs_24_6_port, shift_in(5) => 
                           negative_inputs_24_5_port, shift_in(4) => 
                           negative_inputs_24_4_port, shift_in(3) => 
                           negative_inputs_24_3_port, shift_in(2) => 
                           negative_inputs_24_2_port, shift_in(1) => 
                           negative_inputs_24_1_port, shift_in(0) => n8, 
                           shift_out(63) => negative_inputs_25_63_port, 
                           shift_out(62) => negative_inputs_25_62_port, 
                           shift_out(61) => negative_inputs_25_61_port, 
                           shift_out(60) => negative_inputs_25_60_port, 
                           shift_out(59) => negative_inputs_25_59_port, 
                           shift_out(58) => negative_inputs_25_58_port, 
                           shift_out(57) => negative_inputs_25_57_port, 
                           shift_out(56) => negative_inputs_25_56_port, 
                           shift_out(55) => negative_inputs_25_55_port, 
                           shift_out(54) => negative_inputs_25_54_port, 
                           shift_out(53) => negative_inputs_25_53_port, 
                           shift_out(52) => negative_inputs_25_52_port, 
                           shift_out(51) => negative_inputs_25_51_port, 
                           shift_out(50) => negative_inputs_25_50_port, 
                           shift_out(49) => negative_inputs_25_49_port, 
                           shift_out(48) => negative_inputs_25_48_port, 
                           shift_out(47) => negative_inputs_25_47_port, 
                           shift_out(46) => negative_inputs_25_46_port, 
                           shift_out(45) => negative_inputs_25_45_port, 
                           shift_out(44) => negative_inputs_25_44_port, 
                           shift_out(43) => negative_inputs_25_43_port, 
                           shift_out(42) => negative_inputs_25_42_port, 
                           shift_out(41) => negative_inputs_25_41_port, 
                           shift_out(40) => negative_inputs_25_40_port, 
                           shift_out(39) => negative_inputs_25_39_port, 
                           shift_out(38) => negative_inputs_25_38_port, 
                           shift_out(37) => negative_inputs_25_37_port, 
                           shift_out(36) => negative_inputs_25_36_port, 
                           shift_out(35) => negative_inputs_25_35_port, 
                           shift_out(34) => negative_inputs_25_34_port, 
                           shift_out(33) => negative_inputs_25_33_port, 
                           shift_out(32) => negative_inputs_25_32_port, 
                           shift_out(31) => negative_inputs_25_31_port, 
                           shift_out(30) => negative_inputs_25_30_port, 
                           shift_out(29) => negative_inputs_25_29_port, 
                           shift_out(28) => negative_inputs_25_28_port, 
                           shift_out(27) => negative_inputs_25_27_port, 
                           shift_out(26) => negative_inputs_25_26_port, 
                           shift_out(25) => negative_inputs_25_25_port, 
                           shift_out(24) => negative_inputs_25_24_port, 
                           shift_out(23) => negative_inputs_25_23_port, 
                           shift_out(22) => negative_inputs_25_22_port, 
                           shift_out(21) => negative_inputs_25_21_port, 
                           shift_out(20) => negative_inputs_25_20_port, 
                           shift_out(19) => negative_inputs_25_19_port, 
                           shift_out(18) => negative_inputs_25_18_port, 
                           shift_out(17) => negative_inputs_25_17_port, 
                           shift_out(16) => negative_inputs_25_16_port, 
                           shift_out(15) => negative_inputs_25_15_port, 
                           shift_out(14) => negative_inputs_25_14_port, 
                           shift_out(13) => negative_inputs_25_13_port, 
                           shift_out(12) => negative_inputs_25_12_port, 
                           shift_out(11) => negative_inputs_25_11_port, 
                           shift_out(10) => negative_inputs_25_10_port, 
                           shift_out(9) => negative_inputs_25_9_port, 
                           shift_out(8) => negative_inputs_25_8_port, 
                           shift_out(7) => negative_inputs_25_7_port, 
                           shift_out(6) => negative_inputs_25_6_port, 
                           shift_out(5) => negative_inputs_25_5_port, 
                           shift_out(4) => negative_inputs_25_4_port, 
                           shift_out(3) => negative_inputs_25_3_port, 
                           shift_out(2) => negative_inputs_25_2_port, 
                           shift_out(1) => negative_inputs_25_1_port, 
                           shift_out(0) => n_1120);
   shifted_neg_26 : leftshifter_NbitShifter64_69 port map( shift_in(63) => 
                           negative_inputs_25_63_port, shift_in(62) => 
                           negative_inputs_25_62_port, shift_in(61) => 
                           negative_inputs_25_61_port, shift_in(60) => 
                           negative_inputs_25_60_port, shift_in(59) => 
                           negative_inputs_25_59_port, shift_in(58) => 
                           negative_inputs_25_58_port, shift_in(57) => 
                           negative_inputs_25_57_port, shift_in(56) => 
                           negative_inputs_25_56_port, shift_in(55) => 
                           negative_inputs_25_55_port, shift_in(54) => 
                           negative_inputs_25_54_port, shift_in(53) => 
                           negative_inputs_25_53_port, shift_in(52) => 
                           negative_inputs_25_52_port, shift_in(51) => 
                           negative_inputs_25_51_port, shift_in(50) => 
                           negative_inputs_25_50_port, shift_in(49) => 
                           negative_inputs_25_49_port, shift_in(48) => 
                           negative_inputs_25_48_port, shift_in(47) => 
                           negative_inputs_25_47_port, shift_in(46) => 
                           negative_inputs_25_46_port, shift_in(45) => 
                           negative_inputs_25_45_port, shift_in(44) => 
                           negative_inputs_25_44_port, shift_in(43) => 
                           negative_inputs_25_43_port, shift_in(42) => 
                           negative_inputs_25_42_port, shift_in(41) => 
                           negative_inputs_25_41_port, shift_in(40) => 
                           negative_inputs_25_40_port, shift_in(39) => 
                           negative_inputs_25_39_port, shift_in(38) => 
                           negative_inputs_25_38_port, shift_in(37) => 
                           negative_inputs_25_37_port, shift_in(36) => 
                           negative_inputs_25_36_port, shift_in(35) => 
                           negative_inputs_25_35_port, shift_in(34) => 
                           negative_inputs_25_34_port, shift_in(33) => 
                           negative_inputs_25_33_port, shift_in(32) => 
                           negative_inputs_25_32_port, shift_in(31) => 
                           negative_inputs_25_31_port, shift_in(30) => 
                           negative_inputs_25_30_port, shift_in(29) => 
                           negative_inputs_25_29_port, shift_in(28) => 
                           negative_inputs_25_28_port, shift_in(27) => 
                           negative_inputs_25_27_port, shift_in(26) => 
                           negative_inputs_25_26_port, shift_in(25) => 
                           negative_inputs_25_25_port, shift_in(24) => 
                           negative_inputs_25_24_port, shift_in(23) => 
                           negative_inputs_25_23_port, shift_in(22) => 
                           negative_inputs_25_22_port, shift_in(21) => 
                           negative_inputs_25_21_port, shift_in(20) => 
                           negative_inputs_25_20_port, shift_in(19) => 
                           negative_inputs_25_19_port, shift_in(18) => 
                           negative_inputs_25_18_port, shift_in(17) => 
                           negative_inputs_25_17_port, shift_in(16) => 
                           negative_inputs_25_16_port, shift_in(15) => 
                           negative_inputs_25_15_port, shift_in(14) => 
                           negative_inputs_25_14_port, shift_in(13) => 
                           negative_inputs_25_13_port, shift_in(12) => 
                           negative_inputs_25_12_port, shift_in(11) => 
                           negative_inputs_25_11_port, shift_in(10) => 
                           negative_inputs_25_10_port, shift_in(9) => 
                           negative_inputs_25_9_port, shift_in(8) => 
                           negative_inputs_25_8_port, shift_in(7) => 
                           negative_inputs_25_7_port, shift_in(6) => 
                           negative_inputs_25_6_port, shift_in(5) => 
                           negative_inputs_25_5_port, shift_in(4) => 
                           negative_inputs_25_4_port, shift_in(3) => 
                           negative_inputs_25_3_port, shift_in(2) => 
                           negative_inputs_25_2_port, shift_in(1) => 
                           negative_inputs_25_1_port, shift_in(0) => n8, 
                           shift_out(63) => negative_inputs_26_63_port, 
                           shift_out(62) => negative_inputs_26_62_port, 
                           shift_out(61) => negative_inputs_26_61_port, 
                           shift_out(60) => negative_inputs_26_60_port, 
                           shift_out(59) => negative_inputs_26_59_port, 
                           shift_out(58) => negative_inputs_26_58_port, 
                           shift_out(57) => negative_inputs_26_57_port, 
                           shift_out(56) => negative_inputs_26_56_port, 
                           shift_out(55) => negative_inputs_26_55_port, 
                           shift_out(54) => negative_inputs_26_54_port, 
                           shift_out(53) => negative_inputs_26_53_port, 
                           shift_out(52) => negative_inputs_26_52_port, 
                           shift_out(51) => negative_inputs_26_51_port, 
                           shift_out(50) => negative_inputs_26_50_port, 
                           shift_out(49) => negative_inputs_26_49_port, 
                           shift_out(48) => negative_inputs_26_48_port, 
                           shift_out(47) => negative_inputs_26_47_port, 
                           shift_out(46) => negative_inputs_26_46_port, 
                           shift_out(45) => negative_inputs_26_45_port, 
                           shift_out(44) => negative_inputs_26_44_port, 
                           shift_out(43) => negative_inputs_26_43_port, 
                           shift_out(42) => negative_inputs_26_42_port, 
                           shift_out(41) => negative_inputs_26_41_port, 
                           shift_out(40) => negative_inputs_26_40_port, 
                           shift_out(39) => negative_inputs_26_39_port, 
                           shift_out(38) => negative_inputs_26_38_port, 
                           shift_out(37) => negative_inputs_26_37_port, 
                           shift_out(36) => negative_inputs_26_36_port, 
                           shift_out(35) => negative_inputs_26_35_port, 
                           shift_out(34) => negative_inputs_26_34_port, 
                           shift_out(33) => negative_inputs_26_33_port, 
                           shift_out(32) => negative_inputs_26_32_port, 
                           shift_out(31) => negative_inputs_26_31_port, 
                           shift_out(30) => negative_inputs_26_30_port, 
                           shift_out(29) => negative_inputs_26_29_port, 
                           shift_out(28) => negative_inputs_26_28_port, 
                           shift_out(27) => negative_inputs_26_27_port, 
                           shift_out(26) => negative_inputs_26_26_port, 
                           shift_out(25) => negative_inputs_26_25_port, 
                           shift_out(24) => negative_inputs_26_24_port, 
                           shift_out(23) => negative_inputs_26_23_port, 
                           shift_out(22) => negative_inputs_26_22_port, 
                           shift_out(21) => negative_inputs_26_21_port, 
                           shift_out(20) => negative_inputs_26_20_port, 
                           shift_out(19) => negative_inputs_26_19_port, 
                           shift_out(18) => negative_inputs_26_18_port, 
                           shift_out(17) => negative_inputs_26_17_port, 
                           shift_out(16) => negative_inputs_26_16_port, 
                           shift_out(15) => negative_inputs_26_15_port, 
                           shift_out(14) => negative_inputs_26_14_port, 
                           shift_out(13) => negative_inputs_26_13_port, 
                           shift_out(12) => negative_inputs_26_12_port, 
                           shift_out(11) => negative_inputs_26_11_port, 
                           shift_out(10) => negative_inputs_26_10_port, 
                           shift_out(9) => negative_inputs_26_9_port, 
                           shift_out(8) => negative_inputs_26_8_port, 
                           shift_out(7) => negative_inputs_26_7_port, 
                           shift_out(6) => negative_inputs_26_6_port, 
                           shift_out(5) => negative_inputs_26_5_port, 
                           shift_out(4) => negative_inputs_26_4_port, 
                           shift_out(3) => negative_inputs_26_3_port, 
                           shift_out(2) => negative_inputs_26_2_port, 
                           shift_out(1) => negative_inputs_26_1_port, 
                           shift_out(0) => n_1121);
   shifted_neg_27 : leftshifter_NbitShifter64_68 port map( shift_in(63) => 
                           negative_inputs_26_63_port, shift_in(62) => 
                           negative_inputs_26_62_port, shift_in(61) => 
                           negative_inputs_26_61_port, shift_in(60) => 
                           negative_inputs_26_60_port, shift_in(59) => 
                           negative_inputs_26_59_port, shift_in(58) => 
                           negative_inputs_26_58_port, shift_in(57) => 
                           negative_inputs_26_57_port, shift_in(56) => 
                           negative_inputs_26_56_port, shift_in(55) => 
                           negative_inputs_26_55_port, shift_in(54) => 
                           negative_inputs_26_54_port, shift_in(53) => 
                           negative_inputs_26_53_port, shift_in(52) => 
                           negative_inputs_26_52_port, shift_in(51) => 
                           negative_inputs_26_51_port, shift_in(50) => 
                           negative_inputs_26_50_port, shift_in(49) => 
                           negative_inputs_26_49_port, shift_in(48) => 
                           negative_inputs_26_48_port, shift_in(47) => 
                           negative_inputs_26_47_port, shift_in(46) => 
                           negative_inputs_26_46_port, shift_in(45) => 
                           negative_inputs_26_45_port, shift_in(44) => 
                           negative_inputs_26_44_port, shift_in(43) => 
                           negative_inputs_26_43_port, shift_in(42) => 
                           negative_inputs_26_42_port, shift_in(41) => 
                           negative_inputs_26_41_port, shift_in(40) => 
                           negative_inputs_26_40_port, shift_in(39) => 
                           negative_inputs_26_39_port, shift_in(38) => 
                           negative_inputs_26_38_port, shift_in(37) => 
                           negative_inputs_26_37_port, shift_in(36) => 
                           negative_inputs_26_36_port, shift_in(35) => 
                           negative_inputs_26_35_port, shift_in(34) => 
                           negative_inputs_26_34_port, shift_in(33) => 
                           negative_inputs_26_33_port, shift_in(32) => 
                           negative_inputs_26_32_port, shift_in(31) => 
                           negative_inputs_26_31_port, shift_in(30) => 
                           negative_inputs_26_30_port, shift_in(29) => 
                           negative_inputs_26_29_port, shift_in(28) => 
                           negative_inputs_26_28_port, shift_in(27) => 
                           negative_inputs_26_27_port, shift_in(26) => 
                           negative_inputs_26_26_port, shift_in(25) => 
                           negative_inputs_26_25_port, shift_in(24) => 
                           negative_inputs_26_24_port, shift_in(23) => 
                           negative_inputs_26_23_port, shift_in(22) => 
                           negative_inputs_26_22_port, shift_in(21) => 
                           negative_inputs_26_21_port, shift_in(20) => 
                           negative_inputs_26_20_port, shift_in(19) => 
                           negative_inputs_26_19_port, shift_in(18) => 
                           negative_inputs_26_18_port, shift_in(17) => 
                           negative_inputs_26_17_port, shift_in(16) => 
                           negative_inputs_26_16_port, shift_in(15) => 
                           negative_inputs_26_15_port, shift_in(14) => 
                           negative_inputs_26_14_port, shift_in(13) => 
                           negative_inputs_26_13_port, shift_in(12) => 
                           negative_inputs_26_12_port, shift_in(11) => 
                           negative_inputs_26_11_port, shift_in(10) => 
                           negative_inputs_26_10_port, shift_in(9) => 
                           negative_inputs_26_9_port, shift_in(8) => 
                           negative_inputs_26_8_port, shift_in(7) => 
                           negative_inputs_26_7_port, shift_in(6) => 
                           negative_inputs_26_6_port, shift_in(5) => 
                           negative_inputs_26_5_port, shift_in(4) => 
                           negative_inputs_26_4_port, shift_in(3) => 
                           negative_inputs_26_3_port, shift_in(2) => 
                           negative_inputs_26_2_port, shift_in(1) => 
                           negative_inputs_26_1_port, shift_in(0) => n8, 
                           shift_out(63) => negative_inputs_27_63_port, 
                           shift_out(62) => negative_inputs_27_62_port, 
                           shift_out(61) => negative_inputs_27_61_port, 
                           shift_out(60) => negative_inputs_27_60_port, 
                           shift_out(59) => negative_inputs_27_59_port, 
                           shift_out(58) => negative_inputs_27_58_port, 
                           shift_out(57) => negative_inputs_27_57_port, 
                           shift_out(56) => negative_inputs_27_56_port, 
                           shift_out(55) => negative_inputs_27_55_port, 
                           shift_out(54) => negative_inputs_27_54_port, 
                           shift_out(53) => negative_inputs_27_53_port, 
                           shift_out(52) => negative_inputs_27_52_port, 
                           shift_out(51) => negative_inputs_27_51_port, 
                           shift_out(50) => negative_inputs_27_50_port, 
                           shift_out(49) => negative_inputs_27_49_port, 
                           shift_out(48) => negative_inputs_27_48_port, 
                           shift_out(47) => negative_inputs_27_47_port, 
                           shift_out(46) => negative_inputs_27_46_port, 
                           shift_out(45) => negative_inputs_27_45_port, 
                           shift_out(44) => negative_inputs_27_44_port, 
                           shift_out(43) => negative_inputs_27_43_port, 
                           shift_out(42) => negative_inputs_27_42_port, 
                           shift_out(41) => negative_inputs_27_41_port, 
                           shift_out(40) => negative_inputs_27_40_port, 
                           shift_out(39) => negative_inputs_27_39_port, 
                           shift_out(38) => negative_inputs_27_38_port, 
                           shift_out(37) => negative_inputs_27_37_port, 
                           shift_out(36) => negative_inputs_27_36_port, 
                           shift_out(35) => negative_inputs_27_35_port, 
                           shift_out(34) => negative_inputs_27_34_port, 
                           shift_out(33) => negative_inputs_27_33_port, 
                           shift_out(32) => negative_inputs_27_32_port, 
                           shift_out(31) => negative_inputs_27_31_port, 
                           shift_out(30) => negative_inputs_27_30_port, 
                           shift_out(29) => negative_inputs_27_29_port, 
                           shift_out(28) => negative_inputs_27_28_port, 
                           shift_out(27) => negative_inputs_27_27_port, 
                           shift_out(26) => negative_inputs_27_26_port, 
                           shift_out(25) => negative_inputs_27_25_port, 
                           shift_out(24) => negative_inputs_27_24_port, 
                           shift_out(23) => negative_inputs_27_23_port, 
                           shift_out(22) => negative_inputs_27_22_port, 
                           shift_out(21) => negative_inputs_27_21_port, 
                           shift_out(20) => negative_inputs_27_20_port, 
                           shift_out(19) => negative_inputs_27_19_port, 
                           shift_out(18) => negative_inputs_27_18_port, 
                           shift_out(17) => negative_inputs_27_17_port, 
                           shift_out(16) => negative_inputs_27_16_port, 
                           shift_out(15) => negative_inputs_27_15_port, 
                           shift_out(14) => negative_inputs_27_14_port, 
                           shift_out(13) => negative_inputs_27_13_port, 
                           shift_out(12) => negative_inputs_27_12_port, 
                           shift_out(11) => negative_inputs_27_11_port, 
                           shift_out(10) => negative_inputs_27_10_port, 
                           shift_out(9) => negative_inputs_27_9_port, 
                           shift_out(8) => negative_inputs_27_8_port, 
                           shift_out(7) => negative_inputs_27_7_port, 
                           shift_out(6) => negative_inputs_27_6_port, 
                           shift_out(5) => negative_inputs_27_5_port, 
                           shift_out(4) => negative_inputs_27_4_port, 
                           shift_out(3) => negative_inputs_27_3_port, 
                           shift_out(2) => negative_inputs_27_2_port, 
                           shift_out(1) => negative_inputs_27_1_port, 
                           shift_out(0) => n_1122);
   shifted_neg_28 : leftshifter_NbitShifter64_67 port map( shift_in(63) => 
                           negative_inputs_27_63_port, shift_in(62) => 
                           negative_inputs_27_62_port, shift_in(61) => 
                           negative_inputs_27_61_port, shift_in(60) => 
                           negative_inputs_27_60_port, shift_in(59) => 
                           negative_inputs_27_59_port, shift_in(58) => 
                           negative_inputs_27_58_port, shift_in(57) => 
                           negative_inputs_27_57_port, shift_in(56) => 
                           negative_inputs_27_56_port, shift_in(55) => 
                           negative_inputs_27_55_port, shift_in(54) => 
                           negative_inputs_27_54_port, shift_in(53) => 
                           negative_inputs_27_53_port, shift_in(52) => 
                           negative_inputs_27_52_port, shift_in(51) => 
                           negative_inputs_27_51_port, shift_in(50) => 
                           negative_inputs_27_50_port, shift_in(49) => 
                           negative_inputs_27_49_port, shift_in(48) => 
                           negative_inputs_27_48_port, shift_in(47) => 
                           negative_inputs_27_47_port, shift_in(46) => 
                           negative_inputs_27_46_port, shift_in(45) => 
                           negative_inputs_27_45_port, shift_in(44) => 
                           negative_inputs_27_44_port, shift_in(43) => 
                           negative_inputs_27_43_port, shift_in(42) => 
                           negative_inputs_27_42_port, shift_in(41) => 
                           negative_inputs_27_41_port, shift_in(40) => 
                           negative_inputs_27_40_port, shift_in(39) => 
                           negative_inputs_27_39_port, shift_in(38) => 
                           negative_inputs_27_38_port, shift_in(37) => 
                           negative_inputs_27_37_port, shift_in(36) => 
                           negative_inputs_27_36_port, shift_in(35) => 
                           negative_inputs_27_35_port, shift_in(34) => 
                           negative_inputs_27_34_port, shift_in(33) => 
                           negative_inputs_27_33_port, shift_in(32) => 
                           negative_inputs_27_32_port, shift_in(31) => 
                           negative_inputs_27_31_port, shift_in(30) => 
                           negative_inputs_27_30_port, shift_in(29) => 
                           negative_inputs_27_29_port, shift_in(28) => 
                           negative_inputs_27_28_port, shift_in(27) => 
                           negative_inputs_27_27_port, shift_in(26) => 
                           negative_inputs_27_26_port, shift_in(25) => 
                           negative_inputs_27_25_port, shift_in(24) => 
                           negative_inputs_27_24_port, shift_in(23) => 
                           negative_inputs_27_23_port, shift_in(22) => 
                           negative_inputs_27_22_port, shift_in(21) => 
                           negative_inputs_27_21_port, shift_in(20) => 
                           negative_inputs_27_20_port, shift_in(19) => 
                           negative_inputs_27_19_port, shift_in(18) => 
                           negative_inputs_27_18_port, shift_in(17) => 
                           negative_inputs_27_17_port, shift_in(16) => 
                           negative_inputs_27_16_port, shift_in(15) => 
                           negative_inputs_27_15_port, shift_in(14) => 
                           negative_inputs_27_14_port, shift_in(13) => 
                           negative_inputs_27_13_port, shift_in(12) => 
                           negative_inputs_27_12_port, shift_in(11) => 
                           negative_inputs_27_11_port, shift_in(10) => 
                           negative_inputs_27_10_port, shift_in(9) => 
                           negative_inputs_27_9_port, shift_in(8) => 
                           negative_inputs_27_8_port, shift_in(7) => 
                           negative_inputs_27_7_port, shift_in(6) => 
                           negative_inputs_27_6_port, shift_in(5) => 
                           negative_inputs_27_5_port, shift_in(4) => 
                           negative_inputs_27_4_port, shift_in(3) => 
                           negative_inputs_27_3_port, shift_in(2) => 
                           negative_inputs_27_2_port, shift_in(1) => 
                           negative_inputs_27_1_port, shift_in(0) => n8, 
                           shift_out(63) => negative_inputs_28_63_port, 
                           shift_out(62) => negative_inputs_28_62_port, 
                           shift_out(61) => negative_inputs_28_61_port, 
                           shift_out(60) => negative_inputs_28_60_port, 
                           shift_out(59) => negative_inputs_28_59_port, 
                           shift_out(58) => negative_inputs_28_58_port, 
                           shift_out(57) => negative_inputs_28_57_port, 
                           shift_out(56) => negative_inputs_28_56_port, 
                           shift_out(55) => negative_inputs_28_55_port, 
                           shift_out(54) => negative_inputs_28_54_port, 
                           shift_out(53) => negative_inputs_28_53_port, 
                           shift_out(52) => negative_inputs_28_52_port, 
                           shift_out(51) => negative_inputs_28_51_port, 
                           shift_out(50) => negative_inputs_28_50_port, 
                           shift_out(49) => negative_inputs_28_49_port, 
                           shift_out(48) => negative_inputs_28_48_port, 
                           shift_out(47) => negative_inputs_28_47_port, 
                           shift_out(46) => negative_inputs_28_46_port, 
                           shift_out(45) => negative_inputs_28_45_port, 
                           shift_out(44) => negative_inputs_28_44_port, 
                           shift_out(43) => negative_inputs_28_43_port, 
                           shift_out(42) => negative_inputs_28_42_port, 
                           shift_out(41) => negative_inputs_28_41_port, 
                           shift_out(40) => negative_inputs_28_40_port, 
                           shift_out(39) => negative_inputs_28_39_port, 
                           shift_out(38) => negative_inputs_28_38_port, 
                           shift_out(37) => negative_inputs_28_37_port, 
                           shift_out(36) => negative_inputs_28_36_port, 
                           shift_out(35) => negative_inputs_28_35_port, 
                           shift_out(34) => negative_inputs_28_34_port, 
                           shift_out(33) => negative_inputs_28_33_port, 
                           shift_out(32) => negative_inputs_28_32_port, 
                           shift_out(31) => negative_inputs_28_31_port, 
                           shift_out(30) => negative_inputs_28_30_port, 
                           shift_out(29) => negative_inputs_28_29_port, 
                           shift_out(28) => negative_inputs_28_28_port, 
                           shift_out(27) => negative_inputs_28_27_port, 
                           shift_out(26) => negative_inputs_28_26_port, 
                           shift_out(25) => negative_inputs_28_25_port, 
                           shift_out(24) => negative_inputs_28_24_port, 
                           shift_out(23) => negative_inputs_28_23_port, 
                           shift_out(22) => negative_inputs_28_22_port, 
                           shift_out(21) => negative_inputs_28_21_port, 
                           shift_out(20) => negative_inputs_28_20_port, 
                           shift_out(19) => negative_inputs_28_19_port, 
                           shift_out(18) => negative_inputs_28_18_port, 
                           shift_out(17) => negative_inputs_28_17_port, 
                           shift_out(16) => negative_inputs_28_16_port, 
                           shift_out(15) => negative_inputs_28_15_port, 
                           shift_out(14) => negative_inputs_28_14_port, 
                           shift_out(13) => negative_inputs_28_13_port, 
                           shift_out(12) => negative_inputs_28_12_port, 
                           shift_out(11) => negative_inputs_28_11_port, 
                           shift_out(10) => negative_inputs_28_10_port, 
                           shift_out(9) => negative_inputs_28_9_port, 
                           shift_out(8) => negative_inputs_28_8_port, 
                           shift_out(7) => negative_inputs_28_7_port, 
                           shift_out(6) => negative_inputs_28_6_port, 
                           shift_out(5) => negative_inputs_28_5_port, 
                           shift_out(4) => negative_inputs_28_4_port, 
                           shift_out(3) => negative_inputs_28_3_port, 
                           shift_out(2) => negative_inputs_28_2_port, 
                           shift_out(1) => negative_inputs_28_1_port, 
                           shift_out(0) => n_1123);
   shifted_neg_29 : leftshifter_NbitShifter64_66 port map( shift_in(63) => 
                           negative_inputs_28_63_port, shift_in(62) => 
                           negative_inputs_28_62_port, shift_in(61) => 
                           negative_inputs_28_61_port, shift_in(60) => 
                           negative_inputs_28_60_port, shift_in(59) => 
                           negative_inputs_28_59_port, shift_in(58) => 
                           negative_inputs_28_58_port, shift_in(57) => 
                           negative_inputs_28_57_port, shift_in(56) => 
                           negative_inputs_28_56_port, shift_in(55) => 
                           negative_inputs_28_55_port, shift_in(54) => 
                           negative_inputs_28_54_port, shift_in(53) => 
                           negative_inputs_28_53_port, shift_in(52) => 
                           negative_inputs_28_52_port, shift_in(51) => 
                           negative_inputs_28_51_port, shift_in(50) => 
                           negative_inputs_28_50_port, shift_in(49) => 
                           negative_inputs_28_49_port, shift_in(48) => 
                           negative_inputs_28_48_port, shift_in(47) => 
                           negative_inputs_28_47_port, shift_in(46) => 
                           negative_inputs_28_46_port, shift_in(45) => 
                           negative_inputs_28_45_port, shift_in(44) => 
                           negative_inputs_28_44_port, shift_in(43) => 
                           negative_inputs_28_43_port, shift_in(42) => 
                           negative_inputs_28_42_port, shift_in(41) => 
                           negative_inputs_28_41_port, shift_in(40) => 
                           negative_inputs_28_40_port, shift_in(39) => 
                           negative_inputs_28_39_port, shift_in(38) => 
                           negative_inputs_28_38_port, shift_in(37) => 
                           negative_inputs_28_37_port, shift_in(36) => 
                           negative_inputs_28_36_port, shift_in(35) => 
                           negative_inputs_28_35_port, shift_in(34) => 
                           negative_inputs_28_34_port, shift_in(33) => 
                           negative_inputs_28_33_port, shift_in(32) => 
                           negative_inputs_28_32_port, shift_in(31) => 
                           negative_inputs_28_31_port, shift_in(30) => 
                           negative_inputs_28_30_port, shift_in(29) => 
                           negative_inputs_28_29_port, shift_in(28) => 
                           negative_inputs_28_28_port, shift_in(27) => 
                           negative_inputs_28_27_port, shift_in(26) => 
                           negative_inputs_28_26_port, shift_in(25) => 
                           negative_inputs_28_25_port, shift_in(24) => 
                           negative_inputs_28_24_port, shift_in(23) => 
                           negative_inputs_28_23_port, shift_in(22) => 
                           negative_inputs_28_22_port, shift_in(21) => 
                           negative_inputs_28_21_port, shift_in(20) => 
                           negative_inputs_28_20_port, shift_in(19) => 
                           negative_inputs_28_19_port, shift_in(18) => 
                           negative_inputs_28_18_port, shift_in(17) => 
                           negative_inputs_28_17_port, shift_in(16) => 
                           negative_inputs_28_16_port, shift_in(15) => 
                           negative_inputs_28_15_port, shift_in(14) => 
                           negative_inputs_28_14_port, shift_in(13) => 
                           negative_inputs_28_13_port, shift_in(12) => 
                           negative_inputs_28_12_port, shift_in(11) => 
                           negative_inputs_28_11_port, shift_in(10) => 
                           negative_inputs_28_10_port, shift_in(9) => 
                           negative_inputs_28_9_port, shift_in(8) => 
                           negative_inputs_28_8_port, shift_in(7) => 
                           negative_inputs_28_7_port, shift_in(6) => 
                           negative_inputs_28_6_port, shift_in(5) => 
                           negative_inputs_28_5_port, shift_in(4) => 
                           negative_inputs_28_4_port, shift_in(3) => 
                           negative_inputs_28_3_port, shift_in(2) => 
                           negative_inputs_28_2_port, shift_in(1) => 
                           negative_inputs_28_1_port, shift_in(0) => n8, 
                           shift_out(63) => negative_inputs_29_63_port, 
                           shift_out(62) => negative_inputs_29_62_port, 
                           shift_out(61) => negative_inputs_29_61_port, 
                           shift_out(60) => negative_inputs_29_60_port, 
                           shift_out(59) => negative_inputs_29_59_port, 
                           shift_out(58) => negative_inputs_29_58_port, 
                           shift_out(57) => negative_inputs_29_57_port, 
                           shift_out(56) => negative_inputs_29_56_port, 
                           shift_out(55) => negative_inputs_29_55_port, 
                           shift_out(54) => negative_inputs_29_54_port, 
                           shift_out(53) => negative_inputs_29_53_port, 
                           shift_out(52) => negative_inputs_29_52_port, 
                           shift_out(51) => negative_inputs_29_51_port, 
                           shift_out(50) => negative_inputs_29_50_port, 
                           shift_out(49) => negative_inputs_29_49_port, 
                           shift_out(48) => negative_inputs_29_48_port, 
                           shift_out(47) => negative_inputs_29_47_port, 
                           shift_out(46) => negative_inputs_29_46_port, 
                           shift_out(45) => negative_inputs_29_45_port, 
                           shift_out(44) => negative_inputs_29_44_port, 
                           shift_out(43) => negative_inputs_29_43_port, 
                           shift_out(42) => negative_inputs_29_42_port, 
                           shift_out(41) => negative_inputs_29_41_port, 
                           shift_out(40) => negative_inputs_29_40_port, 
                           shift_out(39) => negative_inputs_29_39_port, 
                           shift_out(38) => negative_inputs_29_38_port, 
                           shift_out(37) => negative_inputs_29_37_port, 
                           shift_out(36) => negative_inputs_29_36_port, 
                           shift_out(35) => negative_inputs_29_35_port, 
                           shift_out(34) => negative_inputs_29_34_port, 
                           shift_out(33) => negative_inputs_29_33_port, 
                           shift_out(32) => negative_inputs_29_32_port, 
                           shift_out(31) => negative_inputs_29_31_port, 
                           shift_out(30) => negative_inputs_29_30_port, 
                           shift_out(29) => negative_inputs_29_29_port, 
                           shift_out(28) => negative_inputs_29_28_port, 
                           shift_out(27) => negative_inputs_29_27_port, 
                           shift_out(26) => negative_inputs_29_26_port, 
                           shift_out(25) => negative_inputs_29_25_port, 
                           shift_out(24) => negative_inputs_29_24_port, 
                           shift_out(23) => negative_inputs_29_23_port, 
                           shift_out(22) => negative_inputs_29_22_port, 
                           shift_out(21) => negative_inputs_29_21_port, 
                           shift_out(20) => negative_inputs_29_20_port, 
                           shift_out(19) => negative_inputs_29_19_port, 
                           shift_out(18) => negative_inputs_29_18_port, 
                           shift_out(17) => negative_inputs_29_17_port, 
                           shift_out(16) => negative_inputs_29_16_port, 
                           shift_out(15) => negative_inputs_29_15_port, 
                           shift_out(14) => negative_inputs_29_14_port, 
                           shift_out(13) => negative_inputs_29_13_port, 
                           shift_out(12) => negative_inputs_29_12_port, 
                           shift_out(11) => negative_inputs_29_11_port, 
                           shift_out(10) => negative_inputs_29_10_port, 
                           shift_out(9) => negative_inputs_29_9_port, 
                           shift_out(8) => negative_inputs_29_8_port, 
                           shift_out(7) => negative_inputs_29_7_port, 
                           shift_out(6) => negative_inputs_29_6_port, 
                           shift_out(5) => negative_inputs_29_5_port, 
                           shift_out(4) => negative_inputs_29_4_port, 
                           shift_out(3) => negative_inputs_29_3_port, 
                           shift_out(2) => negative_inputs_29_2_port, 
                           shift_out(1) => negative_inputs_29_1_port, 
                           shift_out(0) => n_1124);
   shifted_neg_30 : leftshifter_NbitShifter64_65 port map( shift_in(63) => 
                           negative_inputs_29_63_port, shift_in(62) => 
                           negative_inputs_29_62_port, shift_in(61) => 
                           negative_inputs_29_61_port, shift_in(60) => 
                           negative_inputs_29_60_port, shift_in(59) => 
                           negative_inputs_29_59_port, shift_in(58) => 
                           negative_inputs_29_58_port, shift_in(57) => 
                           negative_inputs_29_57_port, shift_in(56) => 
                           negative_inputs_29_56_port, shift_in(55) => 
                           negative_inputs_29_55_port, shift_in(54) => 
                           negative_inputs_29_54_port, shift_in(53) => 
                           negative_inputs_29_53_port, shift_in(52) => 
                           negative_inputs_29_52_port, shift_in(51) => 
                           negative_inputs_29_51_port, shift_in(50) => 
                           negative_inputs_29_50_port, shift_in(49) => 
                           negative_inputs_29_49_port, shift_in(48) => 
                           negative_inputs_29_48_port, shift_in(47) => 
                           negative_inputs_29_47_port, shift_in(46) => 
                           negative_inputs_29_46_port, shift_in(45) => 
                           negative_inputs_29_45_port, shift_in(44) => 
                           negative_inputs_29_44_port, shift_in(43) => 
                           negative_inputs_29_43_port, shift_in(42) => 
                           negative_inputs_29_42_port, shift_in(41) => 
                           negative_inputs_29_41_port, shift_in(40) => 
                           negative_inputs_29_40_port, shift_in(39) => 
                           negative_inputs_29_39_port, shift_in(38) => 
                           negative_inputs_29_38_port, shift_in(37) => 
                           negative_inputs_29_37_port, shift_in(36) => 
                           negative_inputs_29_36_port, shift_in(35) => 
                           negative_inputs_29_35_port, shift_in(34) => 
                           negative_inputs_29_34_port, shift_in(33) => 
                           negative_inputs_29_33_port, shift_in(32) => 
                           negative_inputs_29_32_port, shift_in(31) => 
                           negative_inputs_29_31_port, shift_in(30) => 
                           negative_inputs_29_30_port, shift_in(29) => 
                           negative_inputs_29_29_port, shift_in(28) => 
                           negative_inputs_29_28_port, shift_in(27) => 
                           negative_inputs_29_27_port, shift_in(26) => 
                           negative_inputs_29_26_port, shift_in(25) => 
                           negative_inputs_29_25_port, shift_in(24) => 
                           negative_inputs_29_24_port, shift_in(23) => 
                           negative_inputs_29_23_port, shift_in(22) => 
                           negative_inputs_29_22_port, shift_in(21) => 
                           negative_inputs_29_21_port, shift_in(20) => 
                           negative_inputs_29_20_port, shift_in(19) => 
                           negative_inputs_29_19_port, shift_in(18) => 
                           negative_inputs_29_18_port, shift_in(17) => 
                           negative_inputs_29_17_port, shift_in(16) => 
                           negative_inputs_29_16_port, shift_in(15) => 
                           negative_inputs_29_15_port, shift_in(14) => 
                           negative_inputs_29_14_port, shift_in(13) => 
                           negative_inputs_29_13_port, shift_in(12) => 
                           negative_inputs_29_12_port, shift_in(11) => 
                           negative_inputs_29_11_port, shift_in(10) => 
                           negative_inputs_29_10_port, shift_in(9) => 
                           negative_inputs_29_9_port, shift_in(8) => 
                           negative_inputs_29_8_port, shift_in(7) => 
                           negative_inputs_29_7_port, shift_in(6) => 
                           negative_inputs_29_6_port, shift_in(5) => 
                           negative_inputs_29_5_port, shift_in(4) => 
                           negative_inputs_29_4_port, shift_in(3) => 
                           negative_inputs_29_3_port, shift_in(2) => 
                           negative_inputs_29_2_port, shift_in(1) => 
                           negative_inputs_29_1_port, shift_in(0) => n8, 
                           shift_out(63) => negative_inputs_30_63_port, 
                           shift_out(62) => negative_inputs_30_62_port, 
                           shift_out(61) => negative_inputs_30_61_port, 
                           shift_out(60) => negative_inputs_30_60_port, 
                           shift_out(59) => negative_inputs_30_59_port, 
                           shift_out(58) => negative_inputs_30_58_port, 
                           shift_out(57) => negative_inputs_30_57_port, 
                           shift_out(56) => negative_inputs_30_56_port, 
                           shift_out(55) => negative_inputs_30_55_port, 
                           shift_out(54) => negative_inputs_30_54_port, 
                           shift_out(53) => negative_inputs_30_53_port, 
                           shift_out(52) => negative_inputs_30_52_port, 
                           shift_out(51) => negative_inputs_30_51_port, 
                           shift_out(50) => negative_inputs_30_50_port, 
                           shift_out(49) => negative_inputs_30_49_port, 
                           shift_out(48) => negative_inputs_30_48_port, 
                           shift_out(47) => negative_inputs_30_47_port, 
                           shift_out(46) => negative_inputs_30_46_port, 
                           shift_out(45) => negative_inputs_30_45_port, 
                           shift_out(44) => negative_inputs_30_44_port, 
                           shift_out(43) => negative_inputs_30_43_port, 
                           shift_out(42) => negative_inputs_30_42_port, 
                           shift_out(41) => negative_inputs_30_41_port, 
                           shift_out(40) => negative_inputs_30_40_port, 
                           shift_out(39) => negative_inputs_30_39_port, 
                           shift_out(38) => negative_inputs_30_38_port, 
                           shift_out(37) => negative_inputs_30_37_port, 
                           shift_out(36) => negative_inputs_30_36_port, 
                           shift_out(35) => negative_inputs_30_35_port, 
                           shift_out(34) => negative_inputs_30_34_port, 
                           shift_out(33) => negative_inputs_30_33_port, 
                           shift_out(32) => negative_inputs_30_32_port, 
                           shift_out(31) => negative_inputs_30_31_port, 
                           shift_out(30) => negative_inputs_30_30_port, 
                           shift_out(29) => negative_inputs_30_29_port, 
                           shift_out(28) => negative_inputs_30_28_port, 
                           shift_out(27) => negative_inputs_30_27_port, 
                           shift_out(26) => negative_inputs_30_26_port, 
                           shift_out(25) => negative_inputs_30_25_port, 
                           shift_out(24) => negative_inputs_30_24_port, 
                           shift_out(23) => negative_inputs_30_23_port, 
                           shift_out(22) => negative_inputs_30_22_port, 
                           shift_out(21) => negative_inputs_30_21_port, 
                           shift_out(20) => negative_inputs_30_20_port, 
                           shift_out(19) => negative_inputs_30_19_port, 
                           shift_out(18) => negative_inputs_30_18_port, 
                           shift_out(17) => negative_inputs_30_17_port, 
                           shift_out(16) => negative_inputs_30_16_port, 
                           shift_out(15) => negative_inputs_30_15_port, 
                           shift_out(14) => negative_inputs_30_14_port, 
                           shift_out(13) => negative_inputs_30_13_port, 
                           shift_out(12) => negative_inputs_30_12_port, 
                           shift_out(11) => negative_inputs_30_11_port, 
                           shift_out(10) => negative_inputs_30_10_port, 
                           shift_out(9) => negative_inputs_30_9_port, 
                           shift_out(8) => negative_inputs_30_8_port, 
                           shift_out(7) => negative_inputs_30_7_port, 
                           shift_out(6) => negative_inputs_30_6_port, 
                           shift_out(5) => negative_inputs_30_5_port, 
                           shift_out(4) => negative_inputs_30_4_port, 
                           shift_out(3) => negative_inputs_30_3_port, 
                           shift_out(2) => negative_inputs_30_2_port, 
                           shift_out(1) => negative_inputs_30_1_port, 
                           shift_out(0) => n_1125);
   shifted_neg_31 : leftshifter_NbitShifter64_64 port map( shift_in(63) => 
                           negative_inputs_30_63_port, shift_in(62) => 
                           negative_inputs_30_62_port, shift_in(61) => 
                           negative_inputs_30_61_port, shift_in(60) => 
                           negative_inputs_30_60_port, shift_in(59) => 
                           negative_inputs_30_59_port, shift_in(58) => 
                           negative_inputs_30_58_port, shift_in(57) => 
                           negative_inputs_30_57_port, shift_in(56) => 
                           negative_inputs_30_56_port, shift_in(55) => 
                           negative_inputs_30_55_port, shift_in(54) => 
                           negative_inputs_30_54_port, shift_in(53) => 
                           negative_inputs_30_53_port, shift_in(52) => 
                           negative_inputs_30_52_port, shift_in(51) => 
                           negative_inputs_30_51_port, shift_in(50) => 
                           negative_inputs_30_50_port, shift_in(49) => 
                           negative_inputs_30_49_port, shift_in(48) => 
                           negative_inputs_30_48_port, shift_in(47) => 
                           negative_inputs_30_47_port, shift_in(46) => 
                           negative_inputs_30_46_port, shift_in(45) => 
                           negative_inputs_30_45_port, shift_in(44) => 
                           negative_inputs_30_44_port, shift_in(43) => 
                           negative_inputs_30_43_port, shift_in(42) => 
                           negative_inputs_30_42_port, shift_in(41) => 
                           negative_inputs_30_41_port, shift_in(40) => 
                           negative_inputs_30_40_port, shift_in(39) => 
                           negative_inputs_30_39_port, shift_in(38) => 
                           negative_inputs_30_38_port, shift_in(37) => 
                           negative_inputs_30_37_port, shift_in(36) => 
                           negative_inputs_30_36_port, shift_in(35) => 
                           negative_inputs_30_35_port, shift_in(34) => 
                           negative_inputs_30_34_port, shift_in(33) => 
                           negative_inputs_30_33_port, shift_in(32) => 
                           negative_inputs_30_32_port, shift_in(31) => 
                           negative_inputs_30_31_port, shift_in(30) => 
                           negative_inputs_30_30_port, shift_in(29) => 
                           negative_inputs_30_29_port, shift_in(28) => 
                           negative_inputs_30_28_port, shift_in(27) => 
                           negative_inputs_30_27_port, shift_in(26) => 
                           negative_inputs_30_26_port, shift_in(25) => 
                           negative_inputs_30_25_port, shift_in(24) => 
                           negative_inputs_30_24_port, shift_in(23) => 
                           negative_inputs_30_23_port, shift_in(22) => 
                           negative_inputs_30_22_port, shift_in(21) => 
                           negative_inputs_30_21_port, shift_in(20) => 
                           negative_inputs_30_20_port, shift_in(19) => 
                           negative_inputs_30_19_port, shift_in(18) => 
                           negative_inputs_30_18_port, shift_in(17) => 
                           negative_inputs_30_17_port, shift_in(16) => 
                           negative_inputs_30_16_port, shift_in(15) => 
                           negative_inputs_30_15_port, shift_in(14) => 
                           negative_inputs_30_14_port, shift_in(13) => 
                           negative_inputs_30_13_port, shift_in(12) => 
                           negative_inputs_30_12_port, shift_in(11) => 
                           negative_inputs_30_11_port, shift_in(10) => 
                           negative_inputs_30_10_port, shift_in(9) => 
                           negative_inputs_30_9_port, shift_in(8) => 
                           negative_inputs_30_8_port, shift_in(7) => 
                           negative_inputs_30_7_port, shift_in(6) => 
                           negative_inputs_30_6_port, shift_in(5) => 
                           negative_inputs_30_5_port, shift_in(4) => 
                           negative_inputs_30_4_port, shift_in(3) => 
                           negative_inputs_30_3_port, shift_in(2) => 
                           negative_inputs_30_2_port, shift_in(1) => 
                           negative_inputs_30_1_port, shift_in(0) => n8, 
                           shift_out(63) => negative_inputs_31_63_port, 
                           shift_out(62) => negative_inputs_31_62_port, 
                           shift_out(61) => negative_inputs_31_61_port, 
                           shift_out(60) => negative_inputs_31_60_port, 
                           shift_out(59) => negative_inputs_31_59_port, 
                           shift_out(58) => negative_inputs_31_58_port, 
                           shift_out(57) => negative_inputs_31_57_port, 
                           shift_out(56) => negative_inputs_31_56_port, 
                           shift_out(55) => negative_inputs_31_55_port, 
                           shift_out(54) => negative_inputs_31_54_port, 
                           shift_out(53) => negative_inputs_31_53_port, 
                           shift_out(52) => negative_inputs_31_52_port, 
                           shift_out(51) => negative_inputs_31_51_port, 
                           shift_out(50) => negative_inputs_31_50_port, 
                           shift_out(49) => negative_inputs_31_49_port, 
                           shift_out(48) => negative_inputs_31_48_port, 
                           shift_out(47) => negative_inputs_31_47_port, 
                           shift_out(46) => negative_inputs_31_46_port, 
                           shift_out(45) => negative_inputs_31_45_port, 
                           shift_out(44) => negative_inputs_31_44_port, 
                           shift_out(43) => negative_inputs_31_43_port, 
                           shift_out(42) => negative_inputs_31_42_port, 
                           shift_out(41) => negative_inputs_31_41_port, 
                           shift_out(40) => negative_inputs_31_40_port, 
                           shift_out(39) => negative_inputs_31_39_port, 
                           shift_out(38) => negative_inputs_31_38_port, 
                           shift_out(37) => negative_inputs_31_37_port, 
                           shift_out(36) => negative_inputs_31_36_port, 
                           shift_out(35) => negative_inputs_31_35_port, 
                           shift_out(34) => negative_inputs_31_34_port, 
                           shift_out(33) => negative_inputs_31_33_port, 
                           shift_out(32) => negative_inputs_31_32_port, 
                           shift_out(31) => negative_inputs_31_31_port, 
                           shift_out(30) => negative_inputs_31_30_port, 
                           shift_out(29) => negative_inputs_31_29_port, 
                           shift_out(28) => negative_inputs_31_28_port, 
                           shift_out(27) => negative_inputs_31_27_port, 
                           shift_out(26) => negative_inputs_31_26_port, 
                           shift_out(25) => negative_inputs_31_25_port, 
                           shift_out(24) => negative_inputs_31_24_port, 
                           shift_out(23) => negative_inputs_31_23_port, 
                           shift_out(22) => negative_inputs_31_22_port, 
                           shift_out(21) => negative_inputs_31_21_port, 
                           shift_out(20) => negative_inputs_31_20_port, 
                           shift_out(19) => negative_inputs_31_19_port, 
                           shift_out(18) => negative_inputs_31_18_port, 
                           shift_out(17) => negative_inputs_31_17_port, 
                           shift_out(16) => negative_inputs_31_16_port, 
                           shift_out(15) => negative_inputs_31_15_port, 
                           shift_out(14) => negative_inputs_31_14_port, 
                           shift_out(13) => negative_inputs_31_13_port, 
                           shift_out(12) => negative_inputs_31_12_port, 
                           shift_out(11) => negative_inputs_31_11_port, 
                           shift_out(10) => negative_inputs_31_10_port, 
                           shift_out(9) => negative_inputs_31_9_port, 
                           shift_out(8) => negative_inputs_31_8_port, 
                           shift_out(7) => negative_inputs_31_7_port, 
                           shift_out(6) => negative_inputs_31_6_port, 
                           shift_out(5) => negative_inputs_31_5_port, 
                           shift_out(4) => negative_inputs_31_4_port, 
                           shift_out(3) => negative_inputs_31_3_port, 
                           shift_out(2) => negative_inputs_31_2_port, 
                           shift_out(1) => negative_inputs_31_1_port, 
                           shift_out(0) => n_1126);
   encoder0_0 : encoder_16 port map( pieceofB(2) => B(1), pieceofB(1) => B(0), 
                           pieceofB(0) => X_Logic0_port, sel(2) => sel_0_2_port
                           , sel(1) => sel_0_1_port, sel(0) => sel_0_0_port);
   MUX0_0 : MUX51_MuxNbit64_16 port map( zeroSignal(63) => X_Logic0_port, 
                           zeroSignal(62) => X_Logic0_port, zeroSignal(61) => 
                           X_Logic0_port, zeroSignal(60) => X_Logic0_port, 
                           zeroSignal(59) => X_Logic0_port, zeroSignal(58) => 
                           X_Logic0_port, zeroSignal(57) => X_Logic0_port, 
                           zeroSignal(56) => X_Logic0_port, zeroSignal(55) => 
                           X_Logic0_port, zeroSignal(54) => X_Logic0_port, 
                           zeroSignal(53) => X_Logic0_port, zeroSignal(52) => 
                           X_Logic0_port, zeroSignal(51) => X_Logic0_port, 
                           zeroSignal(50) => X_Logic0_port, zeroSignal(49) => 
                           X_Logic0_port, zeroSignal(48) => X_Logic0_port, 
                           zeroSignal(47) => X_Logic0_port, zeroSignal(46) => 
                           X_Logic0_port, zeroSignal(45) => X_Logic0_port, 
                           zeroSignal(44) => X_Logic0_port, zeroSignal(43) => 
                           X_Logic0_port, zeroSignal(42) => X_Logic0_port, 
                           zeroSignal(41) => X_Logic0_port, zeroSignal(40) => 
                           X_Logic0_port, zeroSignal(39) => X_Logic0_port, 
                           zeroSignal(38) => X_Logic0_port, zeroSignal(37) => 
                           X_Logic0_port, zeroSignal(36) => X_Logic0_port, 
                           zeroSignal(35) => X_Logic0_port, zeroSignal(34) => 
                           X_Logic0_port, zeroSignal(33) => X_Logic0_port, 
                           zeroSignal(32) => X_Logic0_port, zeroSignal(31) => 
                           X_Logic0_port, zeroSignal(30) => X_Logic0_port, 
                           zeroSignal(29) => X_Logic0_port, zeroSignal(28) => 
                           X_Logic0_port, zeroSignal(27) => X_Logic0_port, 
                           zeroSignal(26) => X_Logic0_port, zeroSignal(25) => 
                           X_Logic0_port, zeroSignal(24) => X_Logic0_port, 
                           zeroSignal(23) => X_Logic0_port, zeroSignal(22) => 
                           X_Logic0_port, zeroSignal(21) => X_Logic0_port, 
                           zeroSignal(20) => X_Logic0_port, zeroSignal(19) => 
                           X_Logic0_port, zeroSignal(18) => X_Logic0_port, 
                           zeroSignal(17) => X_Logic0_port, zeroSignal(16) => 
                           X_Logic0_port, zeroSignal(15) => X_Logic0_port, 
                           zeroSignal(14) => X_Logic0_port, zeroSignal(13) => 
                           X_Logic0_port, zeroSignal(12) => X_Logic0_port, 
                           zeroSignal(11) => X_Logic0_port, zeroSignal(10) => 
                           X_Logic0_port, zeroSignal(9) => X_Logic0_port, 
                           zeroSignal(8) => X_Logic0_port, zeroSignal(7) => 
                           X_Logic0_port, zeroSignal(6) => X_Logic0_port, 
                           zeroSignal(5) => X_Logic0_port, zeroSignal(4) => 
                           X_Logic0_port, zeroSignal(3) => X_Logic0_port, 
                           zeroSignal(2) => X_Logic0_port, zeroSignal(1) => 
                           X_Logic0_port, zeroSignal(0) => X_Logic0_port, 
                           A_signal(63) => A(31), A_signal(62) => A(31), 
                           A_signal(61) => A(31), A_signal(60) => A(31), 
                           A_signal(59) => A(31), A_signal(58) => A(31), 
                           A_signal(57) => A(31), A_signal(56) => A(31), 
                           A_signal(55) => A(31), A_signal(54) => A(31), 
                           A_signal(53) => A(31), A_signal(52) => A(31), 
                           A_signal(51) => A(31), A_signal(50) => A(31), 
                           A_signal(49) => A(31), A_signal(48) => A(31), 
                           A_signal(47) => A(31), A_signal(46) => A(31), 
                           A_signal(45) => A(31), A_signal(44) => A(31), 
                           A_signal(43) => A(31), A_signal(42) => A(31), 
                           A_signal(41) => A(31), A_signal(40) => A(31), 
                           A_signal(39) => A(31), A_signal(38) => A(31), 
                           A_signal(37) => A(31), A_signal(36) => A(31), 
                           A_signal(35) => A(31), A_signal(34) => A(31), 
                           A_signal(33) => A(31), A_signal(32) => A(31), 
                           A_signal(31) => A(31), A_signal(30) => A(30), 
                           A_signal(29) => A(29), A_signal(28) => A(28), 
                           A_signal(27) => A(27), A_signal(26) => A(26), 
                           A_signal(25) => A(25), A_signal(24) => A(24), 
                           A_signal(23) => A(23), A_signal(22) => A(22), 
                           A_signal(21) => A(21), A_signal(20) => A(20), 
                           A_signal(19) => A(19), A_signal(18) => A(18), 
                           A_signal(17) => A(17), A_signal(16) => A(16), 
                           A_signal(15) => A(15), A_signal(14) => A(14), 
                           A_signal(13) => A(13), A_signal(12) => A(12), 
                           A_signal(11) => A(11), A_signal(10) => A(10), 
                           A_signal(9) => A(9), A_signal(8) => A(8), 
                           A_signal(7) => A(7), A_signal(6) => A(6), 
                           A_signal(5) => A(5), A_signal(4) => A(4), 
                           A_signal(3) => A(3), A_signal(2) => A(2), 
                           A_signal(1) => n15, A_signal(0) => n18, A_neg(63) =>
                           negative_inputs_0_63_port, A_neg(62) => 
                           negative_inputs_0_62_port, A_neg(61) => 
                           negative_inputs_0_61_port, A_neg(60) => 
                           negative_inputs_0_60_port, A_neg(59) => 
                           negative_inputs_0_59_port, A_neg(58) => 
                           negative_inputs_0_58_port, A_neg(57) => 
                           negative_inputs_0_57_port, A_neg(56) => 
                           negative_inputs_0_56_port, A_neg(55) => 
                           negative_inputs_0_55_port, A_neg(54) => 
                           negative_inputs_0_54_port, A_neg(53) => 
                           negative_inputs_0_53_port, A_neg(52) => n40, 
                           A_neg(51) => n39, A_neg(50) => 
                           negative_inputs_0_50_port, A_neg(49) => n41, 
                           A_neg(48) => negative_inputs_0_48_port, A_neg(47) =>
                           negative_inputs_0_47_port, A_neg(46) => 
                           negative_inputs_0_46_port, A_neg(45) => 
                           negative_inputs_0_45_port, A_neg(44) => 
                           negative_inputs_0_44_port, A_neg(43) => 
                           negative_inputs_0_43_port, A_neg(42) => 
                           negative_inputs_0_42_port, A_neg(41) => 
                           negative_inputs_0_41_port, A_neg(40) => 
                           negative_inputs_0_40_port, A_neg(39) => 
                           negative_inputs_0_39_port, A_neg(38) => 
                           negative_inputs_0_38_port, A_neg(37) => 
                           negative_inputs_0_37_port, A_neg(36) => 
                           negative_inputs_0_36_port, A_neg(35) => 
                           negative_inputs_0_35_port, A_neg(34) => 
                           negative_inputs_0_34_port, A_neg(33) => 
                           negative_inputs_0_33_port, A_neg(32) => 
                           negative_inputs_0_32_port, A_neg(31) => 
                           negative_inputs_0_31_port, A_neg(30) => 
                           negative_inputs_0_30_port, A_neg(29) => 
                           negative_inputs_0_29_port, A_neg(28) => 
                           negative_inputs_0_28_port, A_neg(27) => 
                           negative_inputs_0_27_port, A_neg(26) => 
                           negative_inputs_0_26_port, A_neg(25) => 
                           negative_inputs_0_25_port, A_neg(24) => 
                           negative_inputs_0_24_port, A_neg(23) => 
                           negative_inputs_0_23_port, A_neg(22) => 
                           negative_inputs_0_22_port, A_neg(21) => 
                           negative_inputs_0_21_port, A_neg(20) => 
                           negative_inputs_0_20_port, A_neg(19) => 
                           negative_inputs_0_19_port, A_neg(18) => 
                           negative_inputs_0_18_port, A_neg(17) => 
                           negative_inputs_0_17_port, A_neg(16) => 
                           negative_inputs_0_16_port, A_neg(15) => 
                           negative_inputs_0_15_port, A_neg(14) => 
                           negative_inputs_0_14_port, A_neg(13) => 
                           negative_inputs_0_13_port, A_neg(12) => 
                           negative_inputs_0_12_port, A_neg(11) => 
                           negative_inputs_0_11_port, A_neg(10) => 
                           negative_inputs_0_10_port, A_neg(9) => 
                           negative_inputs_0_9_port, A_neg(8) => 
                           negative_inputs_0_8_port, A_neg(7) => 
                           negative_inputs_0_7_port, A_neg(6) => 
                           negative_inputs_0_6_port, A_neg(5) => 
                           negative_inputs_0_5_port, A_neg(4) => 
                           negative_inputs_0_4_port, A_neg(3) => 
                           negative_inputs_0_3_port, A_neg(2) => 
                           negative_inputs_0_2_port, A_neg(1) => 
                           negative_inputs_0_1_port, A_neg(0) => 
                           negative_inputs_0_0_port, A_shifted(63) => 
                           positive_inputs_1_63_port, A_shifted(62) => 
                           positive_inputs_1_62_port, A_shifted(61) => 
                           positive_inputs_1_61_port, A_shifted(60) => 
                           positive_inputs_1_60_port, A_shifted(59) => 
                           positive_inputs_1_59_port, A_shifted(58) => 
                           positive_inputs_1_58_port, A_shifted(57) => 
                           positive_inputs_1_57_port, A_shifted(56) => 
                           positive_inputs_1_56_port, A_shifted(55) => 
                           positive_inputs_1_55_port, A_shifted(54) => 
                           positive_inputs_1_54_port, A_shifted(53) => 
                           positive_inputs_1_53_port, A_shifted(52) => 
                           positive_inputs_1_52_port, A_shifted(51) => 
                           positive_inputs_1_51_port, A_shifted(50) => 
                           positive_inputs_1_50_port, A_shifted(49) => 
                           positive_inputs_1_49_port, A_shifted(48) => 
                           positive_inputs_1_48_port, A_shifted(47) => 
                           positive_inputs_1_47_port, A_shifted(46) => 
                           positive_inputs_1_46_port, A_shifted(45) => 
                           positive_inputs_1_45_port, A_shifted(44) => 
                           positive_inputs_1_44_port, A_shifted(43) => 
                           positive_inputs_1_43_port, A_shifted(42) => 
                           positive_inputs_1_42_port, A_shifted(41) => 
                           positive_inputs_1_41_port, A_shifted(40) => 
                           positive_inputs_1_40_port, A_shifted(39) => 
                           positive_inputs_1_39_port, A_shifted(38) => 
                           positive_inputs_1_38_port, A_shifted(37) => n24, 
                           A_shifted(36) => positive_inputs_1_36_port, 
                           A_shifted(35) => positive_inputs_1_35_port, 
                           A_shifted(34) => positive_inputs_1_34_port, 
                           A_shifted(33) => positive_inputs_1_33_port, 
                           A_shifted(32) => positive_inputs_1_32_port, 
                           A_shifted(31) => positive_inputs_1_31_port, 
                           A_shifted(30) => positive_inputs_1_30_port, 
                           A_shifted(29) => positive_inputs_1_29_port, 
                           A_shifted(28) => positive_inputs_1_28_port, 
                           A_shifted(27) => positive_inputs_1_27_port, 
                           A_shifted(26) => positive_inputs_1_26_port, 
                           A_shifted(25) => positive_inputs_1_25_port, 
                           A_shifted(24) => positive_inputs_1_24_port, 
                           A_shifted(23) => positive_inputs_1_23_port, 
                           A_shifted(22) => positive_inputs_1_22_port, 
                           A_shifted(21) => positive_inputs_1_21_port, 
                           A_shifted(20) => positive_inputs_1_20_port, 
                           A_shifted(19) => positive_inputs_1_19_port, 
                           A_shifted(18) => positive_inputs_1_18_port, 
                           A_shifted(17) => positive_inputs_1_17_port, 
                           A_shifted(16) => positive_inputs_1_16_port, 
                           A_shifted(15) => positive_inputs_1_15_port, 
                           A_shifted(14) => positive_inputs_1_14_port, 
                           A_shifted(13) => positive_inputs_1_13_port, 
                           A_shifted(12) => positive_inputs_1_12_port, 
                           A_shifted(11) => positive_inputs_1_11_port, 
                           A_shifted(10) => positive_inputs_1_10_port, 
                           A_shifted(9) => positive_inputs_1_9_port, 
                           A_shifted(8) => positive_inputs_1_8_port, 
                           A_shifted(7) => positive_inputs_1_7_port, 
                           A_shifted(6) => positive_inputs_1_6_port, 
                           A_shifted(5) => positive_inputs_1_5_port, 
                           A_shifted(4) => positive_inputs_1_4_port, 
                           A_shifted(3) => positive_inputs_1_3_port, 
                           A_shifted(2) => positive_inputs_1_2_port, 
                           A_shifted(1) => positive_inputs_1_1_port, 
                           A_shifted(0) => n8, A_neg_shifted(63) => 
                           negative_inputs_1_63_port, A_neg_shifted(62) => 
                           negative_inputs_1_62_port, A_neg_shifted(61) => 
                           negative_inputs_1_61_port, A_neg_shifted(60) => 
                           negative_inputs_1_60_port, A_neg_shifted(59) => 
                           negative_inputs_1_59_port, A_neg_shifted(58) => 
                           negative_inputs_1_58_port, A_neg_shifted(57) => 
                           negative_inputs_1_57_port, A_neg_shifted(56) => 
                           negative_inputs_1_56_port, A_neg_shifted(55) => 
                           negative_inputs_1_55_port, A_neg_shifted(54) => 
                           negative_inputs_1_54_port, A_neg_shifted(53) => 
                           negative_inputs_1_53_port, A_neg_shifted(52) => 
                           negative_inputs_1_52_port, A_neg_shifted(51) => 
                           negative_inputs_1_51_port, A_neg_shifted(50) => 
                           negative_inputs_1_50_port, A_neg_shifted(49) => 
                           negative_inputs_1_49_port, A_neg_shifted(48) => 
                           negative_inputs_1_48_port, A_neg_shifted(47) => 
                           negative_inputs_1_47_port, A_neg_shifted(46) => 
                           negative_inputs_1_46_port, A_neg_shifted(45) => 
                           negative_inputs_1_45_port, A_neg_shifted(44) => 
                           negative_inputs_1_44_port, A_neg_shifted(43) => 
                           negative_inputs_1_43_port, A_neg_shifted(42) => 
                           negative_inputs_1_42_port, A_neg_shifted(41) => 
                           negative_inputs_1_41_port, A_neg_shifted(40) => 
                           negative_inputs_1_40_port, A_neg_shifted(39) => 
                           negative_inputs_1_39_port, A_neg_shifted(38) => 
                           negative_inputs_1_38_port, A_neg_shifted(37) => n114
                           , A_neg_shifted(36) => negative_inputs_1_36_port, 
                           A_neg_shifted(35) => negative_inputs_1_35_port, 
                           A_neg_shifted(34) => negative_inputs_1_34_port, 
                           A_neg_shifted(33) => negative_inputs_1_33_port, 
                           A_neg_shifted(32) => negative_inputs_1_32_port, 
                           A_neg_shifted(31) => negative_inputs_1_31_port, 
                           A_neg_shifted(30) => negative_inputs_1_30_port, 
                           A_neg_shifted(29) => negative_inputs_1_29_port, 
                           A_neg_shifted(28) => negative_inputs_1_28_port, 
                           A_neg_shifted(27) => negative_inputs_1_27_port, 
                           A_neg_shifted(26) => negative_inputs_1_26_port, 
                           A_neg_shifted(25) => negative_inputs_1_25_port, 
                           A_neg_shifted(24) => negative_inputs_1_24_port, 
                           A_neg_shifted(23) => negative_inputs_1_23_port, 
                           A_neg_shifted(22) => negative_inputs_1_22_port, 
                           A_neg_shifted(21) => negative_inputs_1_21_port, 
                           A_neg_shifted(20) => negative_inputs_1_20_port, 
                           A_neg_shifted(19) => negative_inputs_1_19_port, 
                           A_neg_shifted(18) => negative_inputs_1_18_port, 
                           A_neg_shifted(17) => negative_inputs_1_17_port, 
                           A_neg_shifted(16) => negative_inputs_1_16_port, 
                           A_neg_shifted(15) => negative_inputs_1_15_port, 
                           A_neg_shifted(14) => negative_inputs_1_14_port, 
                           A_neg_shifted(13) => negative_inputs_1_13_port, 
                           A_neg_shifted(12) => negative_inputs_1_12_port, 
                           A_neg_shifted(11) => negative_inputs_1_11_port, 
                           A_neg_shifted(10) => negative_inputs_1_10_port, 
                           A_neg_shifted(9) => negative_inputs_1_9_port, 
                           A_neg_shifted(8) => negative_inputs_1_8_port, 
                           A_neg_shifted(7) => negative_inputs_1_7_port, 
                           A_neg_shifted(6) => negative_inputs_1_6_port, 
                           A_neg_shifted(5) => negative_inputs_1_5_port, 
                           A_neg_shifted(4) => negative_inputs_1_4_port, 
                           A_neg_shifted(3) => negative_inputs_1_3_port, 
                           A_neg_shifted(2) => negative_inputs_1_2_port, 
                           A_neg_shifted(1) => negative_inputs_1_1_port, 
                           A_neg_shifted(0) => n8, Sel(2) => sel_0_2_port, 
                           Sel(1) => sel_0_1_port, Sel(0) => sel_0_0_port, 
                           Y(63) => MuxOutputs_0_63_port, Y(62) => 
                           MuxOutputs_0_62_port, Y(61) => MuxOutputs_0_61_port,
                           Y(60) => MuxOutputs_0_60_port, Y(59) => 
                           MuxOutputs_0_59_port, Y(58) => MuxOutputs_0_58_port,
                           Y(57) => MuxOutputs_0_57_port, Y(56) => 
                           MuxOutputs_0_56_port, Y(55) => MuxOutputs_0_55_port,
                           Y(54) => MuxOutputs_0_54_port, Y(53) => 
                           MuxOutputs_0_53_port, Y(52) => MuxOutputs_0_52_port,
                           Y(51) => MuxOutputs_0_51_port, Y(50) => 
                           MuxOutputs_0_50_port, Y(49) => MuxOutputs_0_49_port,
                           Y(48) => MuxOutputs_0_48_port, Y(47) => 
                           MuxOutputs_0_47_port, Y(46) => MuxOutputs_0_46_port,
                           Y(45) => MuxOutputs_0_45_port, Y(44) => 
                           MuxOutputs_0_44_port, Y(43) => MuxOutputs_0_43_port,
                           Y(42) => MuxOutputs_0_42_port, Y(41) => 
                           MuxOutputs_0_41_port, Y(40) => MuxOutputs_0_40_port,
                           Y(39) => MuxOutputs_0_39_port, Y(38) => 
                           MuxOutputs_0_38_port, Y(37) => MuxOutputs_0_37_port,
                           Y(36) => MuxOutputs_0_36_port, Y(35) => 
                           MuxOutputs_0_35_port, Y(34) => MuxOutputs_0_34_port,
                           Y(33) => MuxOutputs_0_33_port, Y(32) => 
                           MuxOutputs_0_32_port, Y(31) => MuxOutputs_0_31_port,
                           Y(30) => MuxOutputs_0_30_port, Y(29) => 
                           MuxOutputs_0_29_port, Y(28) => MuxOutputs_0_28_port,
                           Y(27) => MuxOutputs_0_27_port, Y(26) => 
                           MuxOutputs_0_26_port, Y(25) => MuxOutputs_0_25_port,
                           Y(24) => MuxOutputs_0_24_port, Y(23) => 
                           MuxOutputs_0_23_port, Y(22) => MuxOutputs_0_22_port,
                           Y(21) => MuxOutputs_0_21_port, Y(20) => 
                           MuxOutputs_0_20_port, Y(19) => MuxOutputs_0_19_port,
                           Y(18) => MuxOutputs_0_18_port, Y(17) => 
                           MuxOutputs_0_17_port, Y(16) => MuxOutputs_0_16_port,
                           Y(15) => MuxOutputs_0_15_port, Y(14) => 
                           MuxOutputs_0_14_port, Y(13) => MuxOutputs_0_13_port,
                           Y(12) => MuxOutputs_0_12_port, Y(11) => 
                           MuxOutputs_0_11_port, Y(10) => MuxOutputs_0_10_port,
                           Y(9) => MuxOutputs_0_9_port, Y(8) => 
                           MuxOutputs_0_8_port, Y(7) => MuxOutputs_0_7_port, 
                           Y(6) => MuxOutputs_0_6_port, Y(5) => 
                           MuxOutputs_0_5_port, Y(4) => MuxOutputs_0_4_port, 
                           Y(3) => MuxOutputs_0_3_port, Y(2) => 
                           MuxOutputs_0_2_port, Y(1) => MuxOutputs_0_1_port, 
                           Y(0) => MuxOutputs_0_0_port);
   encoderI_1 : encoder_31 port map( pieceofB(2) => B(3), pieceofB(1) => B(2), 
                           pieceofB(0) => B(1), sel(2) => sel_1_2_port, sel(1) 
                           => sel_1_1_port, sel(0) => sel_1_0_port);
   MUXI_1 : MUX51_MuxNbit64_31 port map( zeroSignal(63) => X_Logic0_port, 
                           zeroSignal(62) => X_Logic0_port, zeroSignal(61) => 
                           X_Logic0_port, zeroSignal(60) => X_Logic0_port, 
                           zeroSignal(59) => X_Logic0_port, zeroSignal(58) => 
                           X_Logic0_port, zeroSignal(57) => X_Logic0_port, 
                           zeroSignal(56) => X_Logic0_port, zeroSignal(55) => 
                           X_Logic0_port, zeroSignal(54) => X_Logic0_port, 
                           zeroSignal(53) => X_Logic0_port, zeroSignal(52) => 
                           X_Logic0_port, zeroSignal(51) => X_Logic0_port, 
                           zeroSignal(50) => X_Logic0_port, zeroSignal(49) => 
                           X_Logic0_port, zeroSignal(48) => X_Logic0_port, 
                           zeroSignal(47) => X_Logic0_port, zeroSignal(46) => 
                           X_Logic0_port, zeroSignal(45) => X_Logic0_port, 
                           zeroSignal(44) => X_Logic0_port, zeroSignal(43) => 
                           X_Logic0_port, zeroSignal(42) => X_Logic0_port, 
                           zeroSignal(41) => X_Logic0_port, zeroSignal(40) => 
                           X_Logic0_port, zeroSignal(39) => X_Logic0_port, 
                           zeroSignal(38) => X_Logic0_port, zeroSignal(37) => 
                           X_Logic0_port, zeroSignal(36) => X_Logic0_port, 
                           zeroSignal(35) => X_Logic0_port, zeroSignal(34) => 
                           X_Logic0_port, zeroSignal(33) => X_Logic0_port, 
                           zeroSignal(32) => X_Logic0_port, zeroSignal(31) => 
                           X_Logic0_port, zeroSignal(30) => X_Logic0_port, 
                           zeroSignal(29) => X_Logic0_port, zeroSignal(28) => 
                           X_Logic0_port, zeroSignal(27) => X_Logic0_port, 
                           zeroSignal(26) => X_Logic0_port, zeroSignal(25) => 
                           X_Logic0_port, zeroSignal(24) => X_Logic0_port, 
                           zeroSignal(23) => X_Logic0_port, zeroSignal(22) => 
                           X_Logic0_port, zeroSignal(21) => X_Logic0_port, 
                           zeroSignal(20) => X_Logic0_port, zeroSignal(19) => 
                           X_Logic0_port, zeroSignal(18) => X_Logic0_port, 
                           zeroSignal(17) => X_Logic0_port, zeroSignal(16) => 
                           X_Logic0_port, zeroSignal(15) => X_Logic0_port, 
                           zeroSignal(14) => X_Logic0_port, zeroSignal(13) => 
                           X_Logic0_port, zeroSignal(12) => X_Logic0_port, 
                           zeroSignal(11) => X_Logic0_port, zeroSignal(10) => 
                           X_Logic0_port, zeroSignal(9) => X_Logic0_port, 
                           zeroSignal(8) => X_Logic0_port, zeroSignal(7) => 
                           X_Logic0_port, zeroSignal(6) => X_Logic0_port, 
                           zeroSignal(5) => X_Logic0_port, zeroSignal(4) => 
                           X_Logic0_port, zeroSignal(3) => X_Logic0_port, 
                           zeroSignal(2) => X_Logic0_port, zeroSignal(1) => 
                           X_Logic0_port, zeroSignal(0) => X_Logic0_port, 
                           A_signal(63) => positive_inputs_2_63_port, 
                           A_signal(62) => positive_inputs_2_62_port, 
                           A_signal(61) => positive_inputs_2_61_port, 
                           A_signal(60) => positive_inputs_2_60_port, 
                           A_signal(59) => positive_inputs_2_59_port, 
                           A_signal(58) => positive_inputs_2_58_port, 
                           A_signal(57) => positive_inputs_2_57_port, 
                           A_signal(56) => positive_inputs_2_56_port, 
                           A_signal(55) => positive_inputs_2_55_port, 
                           A_signal(54) => positive_inputs_2_54_port, 
                           A_signal(53) => positive_inputs_2_53_port, 
                           A_signal(52) => positive_inputs_2_52_port, 
                           A_signal(51) => positive_inputs_2_51_port, 
                           A_signal(50) => positive_inputs_2_50_port, 
                           A_signal(49) => positive_inputs_2_49_port, 
                           A_signal(48) => positive_inputs_2_48_port, 
                           A_signal(47) => n38, A_signal(46) => 
                           positive_inputs_2_46_port, A_signal(45) => 
                           positive_inputs_2_45_port, A_signal(44) => 
                           positive_inputs_2_44_port, A_signal(43) => 
                           positive_inputs_2_43_port, A_signal(42) => 
                           positive_inputs_2_42_port, A_signal(41) => 
                           positive_inputs_2_41_port, A_signal(40) => 
                           positive_inputs_2_40_port, A_signal(39) => 
                           positive_inputs_2_39_port, A_signal(38) => 
                           positive_inputs_2_38_port, A_signal(37) => n23, 
                           A_signal(36) => positive_inputs_2_36_port, 
                           A_signal(35) => positive_inputs_2_35_port, 
                           A_signal(34) => positive_inputs_2_34_port, 
                           A_signal(33) => positive_inputs_2_33_port, 
                           A_signal(32) => positive_inputs_2_32_port, 
                           A_signal(31) => positive_inputs_2_31_port, 
                           A_signal(30) => positive_inputs_2_30_port, 
                           A_signal(29) => positive_inputs_2_29_port, 
                           A_signal(28) => positive_inputs_2_28_port, 
                           A_signal(27) => positive_inputs_2_27_port, 
                           A_signal(26) => positive_inputs_2_26_port, 
                           A_signal(25) => positive_inputs_2_25_port, 
                           A_signal(24) => positive_inputs_2_24_port, 
                           A_signal(23) => positive_inputs_2_23_port, 
                           A_signal(22) => positive_inputs_2_22_port, 
                           A_signal(21) => positive_inputs_2_21_port, 
                           A_signal(20) => positive_inputs_2_20_port, 
                           A_signal(19) => positive_inputs_2_19_port, 
                           A_signal(18) => positive_inputs_2_18_port, 
                           A_signal(17) => positive_inputs_2_17_port, 
                           A_signal(16) => positive_inputs_2_16_port, 
                           A_signal(15) => positive_inputs_2_15_port, 
                           A_signal(14) => positive_inputs_2_14_port, 
                           A_signal(13) => positive_inputs_2_13_port, 
                           A_signal(12) => positive_inputs_2_12_port, 
                           A_signal(11) => positive_inputs_2_11_port, 
                           A_signal(10) => positive_inputs_2_10_port, 
                           A_signal(9) => positive_inputs_2_9_port, A_signal(8)
                           => positive_inputs_2_8_port, A_signal(7) => 
                           positive_inputs_2_7_port, A_signal(6) => 
                           positive_inputs_2_6_port, A_signal(5) => 
                           positive_inputs_2_5_port, A_signal(4) => 
                           positive_inputs_2_4_port, A_signal(3) => 
                           positive_inputs_2_3_port, A_signal(2) => 
                           positive_inputs_2_2_port, A_signal(1) => 
                           positive_inputs_2_1_port, A_signal(0) => n8, 
                           A_neg(63) => negative_inputs_2_63_port, A_neg(62) =>
                           negative_inputs_2_62_port, A_neg(61) => 
                           negative_inputs_2_61_port, A_neg(60) => 
                           negative_inputs_2_60_port, A_neg(59) => 
                           negative_inputs_2_59_port, A_neg(58) => 
                           negative_inputs_2_58_port, A_neg(57) => 
                           negative_inputs_2_57_port, A_neg(56) => 
                           negative_inputs_2_56_port, A_neg(55) => 
                           negative_inputs_2_55_port, A_neg(54) => 
                           negative_inputs_2_54_port, A_neg(53) => 
                           negative_inputs_2_53_port, A_neg(52) => 
                           negative_inputs_2_52_port, A_neg(51) => 
                           negative_inputs_2_51_port, A_neg(50) => 
                           negative_inputs_2_50_port, A_neg(49) => 
                           negative_inputs_2_49_port, A_neg(48) => 
                           negative_inputs_2_48_port, A_neg(47) => 
                           negative_inputs_2_47_port, A_neg(46) => 
                           negative_inputs_2_46_port, A_neg(45) => 
                           negative_inputs_2_45_port, A_neg(44) => 
                           negative_inputs_2_44_port, A_neg(43) => 
                           negative_inputs_2_43_port, A_neg(42) => 
                           negative_inputs_2_42_port, A_neg(41) => 
                           negative_inputs_2_41_port, A_neg(40) => 
                           negative_inputs_2_40_port, A_neg(39) => 
                           negative_inputs_2_39_port, A_neg(38) => 
                           negative_inputs_2_38_port, A_neg(37) => n112, 
                           A_neg(36) => negative_inputs_2_36_port, A_neg(35) =>
                           negative_inputs_2_35_port, A_neg(34) => 
                           negative_inputs_2_34_port, A_neg(33) => 
                           negative_inputs_2_33_port, A_neg(32) => 
                           negative_inputs_2_32_port, A_neg(31) => 
                           negative_inputs_2_31_port, A_neg(30) => 
                           negative_inputs_2_30_port, A_neg(29) => 
                           negative_inputs_2_29_port, A_neg(28) => 
                           negative_inputs_2_28_port, A_neg(27) => 
                           negative_inputs_2_27_port, A_neg(26) => 
                           negative_inputs_2_26_port, A_neg(25) => 
                           negative_inputs_2_25_port, A_neg(24) => 
                           negative_inputs_2_24_port, A_neg(23) => 
                           negative_inputs_2_23_port, A_neg(22) => 
                           negative_inputs_2_22_port, A_neg(21) => 
                           negative_inputs_2_21_port, A_neg(20) => 
                           negative_inputs_2_20_port, A_neg(19) => 
                           negative_inputs_2_19_port, A_neg(18) => 
                           negative_inputs_2_18_port, A_neg(17) => 
                           negative_inputs_2_17_port, A_neg(16) => 
                           negative_inputs_2_16_port, A_neg(15) => 
                           negative_inputs_2_15_port, A_neg(14) => 
                           negative_inputs_2_14_port, A_neg(13) => 
                           negative_inputs_2_13_port, A_neg(12) => 
                           negative_inputs_2_12_port, A_neg(11) => 
                           negative_inputs_2_11_port, A_neg(10) => 
                           negative_inputs_2_10_port, A_neg(9) => 
                           negative_inputs_2_9_port, A_neg(8) => 
                           negative_inputs_2_8_port, A_neg(7) => 
                           negative_inputs_2_7_port, A_neg(6) => 
                           negative_inputs_2_6_port, A_neg(5) => 
                           negative_inputs_2_5_port, A_neg(4) => 
                           negative_inputs_2_4_port, A_neg(3) => 
                           negative_inputs_2_3_port, A_neg(2) => 
                           negative_inputs_2_2_port, A_neg(1) => 
                           negative_inputs_2_1_port, A_neg(0) => n8, 
                           A_shifted(63) => positive_inputs_3_63_port, 
                           A_shifted(62) => positive_inputs_3_62_port, 
                           A_shifted(61) => positive_inputs_3_61_port, 
                           A_shifted(60) => positive_inputs_3_60_port, 
                           A_shifted(59) => positive_inputs_3_59_port, 
                           A_shifted(58) => positive_inputs_3_58_port, 
                           A_shifted(57) => positive_inputs_3_57_port, 
                           A_shifted(56) => positive_inputs_3_56_port, 
                           A_shifted(55) => positive_inputs_3_55_port, 
                           A_shifted(54) => positive_inputs_3_54_port, 
                           A_shifted(53) => positive_inputs_3_53_port, 
                           A_shifted(52) => positive_inputs_3_52_port, 
                           A_shifted(51) => positive_inputs_3_51_port, 
                           A_shifted(50) => positive_inputs_3_50_port, 
                           A_shifted(49) => positive_inputs_3_49_port, 
                           A_shifted(48) => positive_inputs_3_48_port, 
                           A_shifted(47) => positive_inputs_3_47_port, 
                           A_shifted(46) => positive_inputs_3_46_port, 
                           A_shifted(45) => positive_inputs_3_45_port, 
                           A_shifted(44) => positive_inputs_3_44_port, 
                           A_shifted(43) => positive_inputs_3_43_port, 
                           A_shifted(42) => positive_inputs_3_42_port, 
                           A_shifted(41) => positive_inputs_3_41_port, 
                           A_shifted(40) => positive_inputs_3_40_port, 
                           A_shifted(39) => positive_inputs_3_39_port, 
                           A_shifted(38) => positive_inputs_3_38_port, 
                           A_shifted(37) => n22, A_shifted(36) => 
                           positive_inputs_3_36_port, A_shifted(35) => 
                           positive_inputs_3_35_port, A_shifted(34) => 
                           positive_inputs_3_34_port, A_shifted(33) => 
                           positive_inputs_3_33_port, A_shifted(32) => 
                           positive_inputs_3_32_port, A_shifted(31) => 
                           positive_inputs_3_31_port, A_shifted(30) => 
                           positive_inputs_3_30_port, A_shifted(29) => 
                           positive_inputs_3_29_port, A_shifted(28) => 
                           positive_inputs_3_28_port, A_shifted(27) => 
                           positive_inputs_3_27_port, A_shifted(26) => 
                           positive_inputs_3_26_port, A_shifted(25) => 
                           positive_inputs_3_25_port, A_shifted(24) => 
                           positive_inputs_3_24_port, A_shifted(23) => 
                           positive_inputs_3_23_port, A_shifted(22) => 
                           positive_inputs_3_22_port, A_shifted(21) => 
                           positive_inputs_3_21_port, A_shifted(20) => 
                           positive_inputs_3_20_port, A_shifted(19) => 
                           positive_inputs_3_19_port, A_shifted(18) => 
                           positive_inputs_3_18_port, A_shifted(17) => 
                           positive_inputs_3_17_port, A_shifted(16) => 
                           positive_inputs_3_16_port, A_shifted(15) => 
                           positive_inputs_3_15_port, A_shifted(14) => 
                           positive_inputs_3_14_port, A_shifted(13) => 
                           positive_inputs_3_13_port, A_shifted(12) => 
                           positive_inputs_3_12_port, A_shifted(11) => 
                           positive_inputs_3_11_port, A_shifted(10) => 
                           positive_inputs_3_10_port, A_shifted(9) => 
                           positive_inputs_3_9_port, A_shifted(8) => 
                           positive_inputs_3_8_port, A_shifted(7) => 
                           positive_inputs_3_7_port, A_shifted(6) => 
                           positive_inputs_3_6_port, A_shifted(5) => 
                           positive_inputs_3_5_port, A_shifted(4) => 
                           positive_inputs_3_4_port, A_shifted(3) => 
                           positive_inputs_3_3_port, A_shifted(2) => 
                           positive_inputs_3_2_port, A_shifted(1) => 
                           positive_inputs_3_1_port, A_shifted(0) => n8, 
                           A_neg_shifted(63) => negative_inputs_3_63_port, 
                           A_neg_shifted(62) => negative_inputs_3_62_port, 
                           A_neg_shifted(61) => negative_inputs_3_61_port, 
                           A_neg_shifted(60) => negative_inputs_3_60_port, 
                           A_neg_shifted(59) => negative_inputs_3_59_port, 
                           A_neg_shifted(58) => negative_inputs_3_58_port, 
                           A_neg_shifted(57) => negative_inputs_3_57_port, 
                           A_neg_shifted(56) => negative_inputs_3_56_port, 
                           A_neg_shifted(55) => negative_inputs_3_55_port, 
                           A_neg_shifted(54) => negative_inputs_3_54_port, 
                           A_neg_shifted(53) => negative_inputs_3_53_port, 
                           A_neg_shifted(52) => negative_inputs_3_52_port, 
                           A_neg_shifted(51) => negative_inputs_3_51_port, 
                           A_neg_shifted(50) => negative_inputs_3_50_port, 
                           A_neg_shifted(49) => negative_inputs_3_49_port, 
                           A_neg_shifted(48) => negative_inputs_3_48_port, 
                           A_neg_shifted(47) => negative_inputs_3_47_port, 
                           A_neg_shifted(46) => negative_inputs_3_46_port, 
                           A_neg_shifted(45) => negative_inputs_3_45_port, 
                           A_neg_shifted(44) => negative_inputs_3_44_port, 
                           A_neg_shifted(43) => negative_inputs_3_43_port, 
                           A_neg_shifted(42) => negative_inputs_3_42_port, 
                           A_neg_shifted(41) => negative_inputs_3_41_port, 
                           A_neg_shifted(40) => negative_inputs_3_40_port, 
                           A_neg_shifted(39) => negative_inputs_3_39_port, 
                           A_neg_shifted(38) => negative_inputs_3_38_port, 
                           A_neg_shifted(37) => n110, A_neg_shifted(36) => 
                           negative_inputs_3_36_port, A_neg_shifted(35) => 
                           negative_inputs_3_35_port, A_neg_shifted(34) => 
                           negative_inputs_3_34_port, A_neg_shifted(33) => 
                           negative_inputs_3_33_port, A_neg_shifted(32) => 
                           negative_inputs_3_32_port, A_neg_shifted(31) => 
                           negative_inputs_3_31_port, A_neg_shifted(30) => 
                           negative_inputs_3_30_port, A_neg_shifted(29) => 
                           negative_inputs_3_29_port, A_neg_shifted(28) => 
                           negative_inputs_3_28_port, A_neg_shifted(27) => 
                           negative_inputs_3_27_port, A_neg_shifted(26) => 
                           negative_inputs_3_26_port, A_neg_shifted(25) => 
                           negative_inputs_3_25_port, A_neg_shifted(24) => 
                           negative_inputs_3_24_port, A_neg_shifted(23) => 
                           negative_inputs_3_23_port, A_neg_shifted(22) => 
                           negative_inputs_3_22_port, A_neg_shifted(21) => 
                           negative_inputs_3_21_port, A_neg_shifted(20) => 
                           negative_inputs_3_20_port, A_neg_shifted(19) => 
                           negative_inputs_3_19_port, A_neg_shifted(18) => 
                           negative_inputs_3_18_port, A_neg_shifted(17) => 
                           negative_inputs_3_17_port, A_neg_shifted(16) => 
                           negative_inputs_3_16_port, A_neg_shifted(15) => 
                           negative_inputs_3_15_port, A_neg_shifted(14) => 
                           negative_inputs_3_14_port, A_neg_shifted(13) => 
                           negative_inputs_3_13_port, A_neg_shifted(12) => 
                           negative_inputs_3_12_port, A_neg_shifted(11) => 
                           negative_inputs_3_11_port, A_neg_shifted(10) => 
                           negative_inputs_3_10_port, A_neg_shifted(9) => 
                           negative_inputs_3_9_port, A_neg_shifted(8) => 
                           negative_inputs_3_8_port, A_neg_shifted(7) => 
                           negative_inputs_3_7_port, A_neg_shifted(6) => 
                           negative_inputs_3_6_port, A_neg_shifted(5) => 
                           negative_inputs_3_5_port, A_neg_shifted(4) => 
                           negative_inputs_3_4_port, A_neg_shifted(3) => 
                           negative_inputs_3_3_port, A_neg_shifted(2) => 
                           negative_inputs_3_2_port, A_neg_shifted(1) => 
                           negative_inputs_3_1_port, A_neg_shifted(0) => n8, 
                           Sel(2) => sel_1_2_port, Sel(1) => sel_1_1_port, 
                           Sel(0) => sel_1_0_port, Y(63) => 
                           MuxOutputs_1_63_port, Y(62) => MuxOutputs_1_62_port,
                           Y(61) => MuxOutputs_1_61_port, Y(60) => 
                           MuxOutputs_1_60_port, Y(59) => MuxOutputs_1_59_port,
                           Y(58) => MuxOutputs_1_58_port, Y(57) => 
                           MuxOutputs_1_57_port, Y(56) => MuxOutputs_1_56_port,
                           Y(55) => MuxOutputs_1_55_port, Y(54) => 
                           MuxOutputs_1_54_port, Y(53) => MuxOutputs_1_53_port,
                           Y(52) => MuxOutputs_1_52_port, Y(51) => 
                           MuxOutputs_1_51_port, Y(50) => MuxOutputs_1_50_port,
                           Y(49) => MuxOutputs_1_49_port, Y(48) => 
                           MuxOutputs_1_48_port, Y(47) => MuxOutputs_1_47_port,
                           Y(46) => MuxOutputs_1_46_port, Y(45) => 
                           MuxOutputs_1_45_port, Y(44) => MuxOutputs_1_44_port,
                           Y(43) => MuxOutputs_1_43_port, Y(42) => 
                           MuxOutputs_1_42_port, Y(41) => MuxOutputs_1_41_port,
                           Y(40) => MuxOutputs_1_40_port, Y(39) => 
                           MuxOutputs_1_39_port, Y(38) => MuxOutputs_1_38_port,
                           Y(37) => MuxOutputs_1_37_port, Y(36) => 
                           MuxOutputs_1_36_port, Y(35) => MuxOutputs_1_35_port,
                           Y(34) => MuxOutputs_1_34_port, Y(33) => 
                           MuxOutputs_1_33_port, Y(32) => MuxOutputs_1_32_port,
                           Y(31) => MuxOutputs_1_31_port, Y(30) => 
                           MuxOutputs_1_30_port, Y(29) => MuxOutputs_1_29_port,
                           Y(28) => MuxOutputs_1_28_port, Y(27) => 
                           MuxOutputs_1_27_port, Y(26) => MuxOutputs_1_26_port,
                           Y(25) => MuxOutputs_1_25_port, Y(24) => 
                           MuxOutputs_1_24_port, Y(23) => MuxOutputs_1_23_port,
                           Y(22) => MuxOutputs_1_22_port, Y(21) => 
                           MuxOutputs_1_21_port, Y(20) => MuxOutputs_1_20_port,
                           Y(19) => MuxOutputs_1_19_port, Y(18) => 
                           MuxOutputs_1_18_port, Y(17) => MuxOutputs_1_17_port,
                           Y(16) => MuxOutputs_1_16_port, Y(15) => 
                           MuxOutputs_1_15_port, Y(14) => MuxOutputs_1_14_port,
                           Y(13) => MuxOutputs_1_13_port, Y(12) => 
                           MuxOutputs_1_12_port, Y(11) => MuxOutputs_1_11_port,
                           Y(10) => MuxOutputs_1_10_port, Y(9) => 
                           MuxOutputs_1_9_port, Y(8) => MuxOutputs_1_8_port, 
                           Y(7) => MuxOutputs_1_7_port, Y(6) => 
                           MuxOutputs_1_6_port, Y(5) => MuxOutputs_1_5_port, 
                           Y(4) => MuxOutputs_1_4_port, Y(3) => 
                           MuxOutputs_1_3_port, Y(2) => MuxOutputs_1_2_port, 
                           Y(1) => MuxOutputs_1_1_port, Y(0) => 
                           MuxOutputs_1_0_port);
   encoderI_2 : encoder_30 port map( pieceofB(2) => B(5), pieceofB(1) => B(4), 
                           pieceofB(0) => B(3), sel(2) => sel_2_2_port, sel(1) 
                           => sel_2_1_port, sel(0) => sel_2_0_port);
   MUXI_2 : MUX51_MuxNbit64_30 port map( zeroSignal(63) => X_Logic0_port, 
                           zeroSignal(62) => X_Logic0_port, zeroSignal(61) => 
                           X_Logic0_port, zeroSignal(60) => X_Logic0_port, 
                           zeroSignal(59) => X_Logic0_port, zeroSignal(58) => 
                           X_Logic0_port, zeroSignal(57) => X_Logic0_port, 
                           zeroSignal(56) => X_Logic0_port, zeroSignal(55) => 
                           X_Logic0_port, zeroSignal(54) => X_Logic0_port, 
                           zeroSignal(53) => X_Logic0_port, zeroSignal(52) => 
                           X_Logic0_port, zeroSignal(51) => X_Logic0_port, 
                           zeroSignal(50) => X_Logic0_port, zeroSignal(49) => 
                           X_Logic0_port, zeroSignal(48) => X_Logic0_port, 
                           zeroSignal(47) => X_Logic0_port, zeroSignal(46) => 
                           X_Logic0_port, zeroSignal(45) => X_Logic0_port, 
                           zeroSignal(44) => X_Logic0_port, zeroSignal(43) => 
                           X_Logic0_port, zeroSignal(42) => X_Logic0_port, 
                           zeroSignal(41) => X_Logic0_port, zeroSignal(40) => 
                           X_Logic0_port, zeroSignal(39) => X_Logic0_port, 
                           zeroSignal(38) => X_Logic0_port, zeroSignal(37) => 
                           X_Logic0_port, zeroSignal(36) => X_Logic0_port, 
                           zeroSignal(35) => X_Logic0_port, zeroSignal(34) => 
                           X_Logic0_port, zeroSignal(33) => X_Logic0_port, 
                           zeroSignal(32) => X_Logic0_port, zeroSignal(31) => 
                           X_Logic0_port, zeroSignal(30) => X_Logic0_port, 
                           zeroSignal(29) => X_Logic0_port, zeroSignal(28) => 
                           X_Logic0_port, zeroSignal(27) => X_Logic0_port, 
                           zeroSignal(26) => X_Logic0_port, zeroSignal(25) => 
                           X_Logic0_port, zeroSignal(24) => X_Logic0_port, 
                           zeroSignal(23) => X_Logic0_port, zeroSignal(22) => 
                           X_Logic0_port, zeroSignal(21) => X_Logic0_port, 
                           zeroSignal(20) => X_Logic0_port, zeroSignal(19) => 
                           X_Logic0_port, zeroSignal(18) => X_Logic0_port, 
                           zeroSignal(17) => X_Logic0_port, zeroSignal(16) => 
                           X_Logic0_port, zeroSignal(15) => X_Logic0_port, 
                           zeroSignal(14) => X_Logic0_port, zeroSignal(13) => 
                           X_Logic0_port, zeroSignal(12) => X_Logic0_port, 
                           zeroSignal(11) => X_Logic0_port, zeroSignal(10) => 
                           X_Logic0_port, zeroSignal(9) => X_Logic0_port, 
                           zeroSignal(8) => X_Logic0_port, zeroSignal(7) => 
                           X_Logic0_port, zeroSignal(6) => X_Logic0_port, 
                           zeroSignal(5) => X_Logic0_port, zeroSignal(4) => 
                           X_Logic0_port, zeroSignal(3) => X_Logic0_port, 
                           zeroSignal(2) => X_Logic0_port, zeroSignal(1) => 
                           X_Logic0_port, zeroSignal(0) => X_Logic0_port, 
                           A_signal(63) => positive_inputs_4_63_port, 
                           A_signal(62) => positive_inputs_4_62_port, 
                           A_signal(61) => positive_inputs_4_61_port, 
                           A_signal(60) => positive_inputs_4_60_port, 
                           A_signal(59) => positive_inputs_4_59_port, 
                           A_signal(58) => positive_inputs_4_58_port, 
                           A_signal(57) => positive_inputs_4_57_port, 
                           A_signal(56) => positive_inputs_4_56_port, 
                           A_signal(55) => positive_inputs_4_55_port, 
                           A_signal(54) => positive_inputs_4_54_port, 
                           A_signal(53) => positive_inputs_4_53_port, 
                           A_signal(52) => positive_inputs_4_52_port, 
                           A_signal(51) => positive_inputs_4_51_port, 
                           A_signal(50) => positive_inputs_4_50_port, 
                           A_signal(49) => positive_inputs_4_49_port, 
                           A_signal(48) => positive_inputs_4_48_port, 
                           A_signal(47) => n37, A_signal(46) => 
                           positive_inputs_4_46_port, A_signal(45) => 
                           positive_inputs_4_45_port, A_signal(44) => 
                           positive_inputs_4_44_port, A_signal(43) => 
                           positive_inputs_4_43_port, A_signal(42) => 
                           positive_inputs_4_42_port, A_signal(41) => 
                           positive_inputs_4_41_port, A_signal(40) => 
                           positive_inputs_4_40_port, A_signal(39) => 
                           positive_inputs_4_39_port, A_signal(38) => 
                           positive_inputs_4_38_port, A_signal(37) => n21, 
                           A_signal(36) => positive_inputs_4_36_port, 
                           A_signal(35) => positive_inputs_4_35_port, 
                           A_signal(34) => positive_inputs_4_34_port, 
                           A_signal(33) => positive_inputs_4_33_port, 
                           A_signal(32) => positive_inputs_4_32_port, 
                           A_signal(31) => positive_inputs_4_31_port, 
                           A_signal(30) => positive_inputs_4_30_port, 
                           A_signal(29) => positive_inputs_4_29_port, 
                           A_signal(28) => positive_inputs_4_28_port, 
                           A_signal(27) => positive_inputs_4_27_port, 
                           A_signal(26) => positive_inputs_4_26_port, 
                           A_signal(25) => positive_inputs_4_25_port, 
                           A_signal(24) => positive_inputs_4_24_port, 
                           A_signal(23) => positive_inputs_4_23_port, 
                           A_signal(22) => positive_inputs_4_22_port, 
                           A_signal(21) => positive_inputs_4_21_port, 
                           A_signal(20) => positive_inputs_4_20_port, 
                           A_signal(19) => positive_inputs_4_19_port, 
                           A_signal(18) => positive_inputs_4_18_port, 
                           A_signal(17) => positive_inputs_4_17_port, 
                           A_signal(16) => positive_inputs_4_16_port, 
                           A_signal(15) => positive_inputs_4_15_port, 
                           A_signal(14) => positive_inputs_4_14_port, 
                           A_signal(13) => positive_inputs_4_13_port, 
                           A_signal(12) => positive_inputs_4_12_port, 
                           A_signal(11) => positive_inputs_4_11_port, 
                           A_signal(10) => positive_inputs_4_10_port, 
                           A_signal(9) => positive_inputs_4_9_port, A_signal(8)
                           => positive_inputs_4_8_port, A_signal(7) => 
                           positive_inputs_4_7_port, A_signal(6) => 
                           positive_inputs_4_6_port, A_signal(5) => 
                           positive_inputs_4_5_port, A_signal(4) => 
                           positive_inputs_4_4_port, A_signal(3) => 
                           positive_inputs_4_3_port, A_signal(2) => 
                           positive_inputs_4_2_port, A_signal(1) => 
                           positive_inputs_4_1_port, A_signal(0) => n8, 
                           A_neg(63) => negative_inputs_4_63_port, A_neg(62) =>
                           negative_inputs_4_62_port, A_neg(61) => 
                           negative_inputs_4_61_port, A_neg(60) => 
                           negative_inputs_4_60_port, A_neg(59) => 
                           negative_inputs_4_59_port, A_neg(58) => 
                           negative_inputs_4_58_port, A_neg(57) => 
                           negative_inputs_4_57_port, A_neg(56) => 
                           negative_inputs_4_56_port, A_neg(55) => 
                           negative_inputs_4_55_port, A_neg(54) => 
                           negative_inputs_4_54_port, A_neg(53) => 
                           negative_inputs_4_53_port, A_neg(52) => 
                           negative_inputs_4_52_port, A_neg(51) => 
                           negative_inputs_4_51_port, A_neg(50) => 
                           negative_inputs_4_50_port, A_neg(49) => 
                           negative_inputs_4_49_port, A_neg(48) => 
                           negative_inputs_4_48_port, A_neg(47) => 
                           negative_inputs_4_47_port, A_neg(46) => 
                           negative_inputs_4_46_port, A_neg(45) => 
                           negative_inputs_4_45_port, A_neg(44) => 
                           negative_inputs_4_44_port, A_neg(43) => 
                           negative_inputs_4_43_port, A_neg(42) => 
                           negative_inputs_4_42_port, A_neg(41) => 
                           negative_inputs_4_41_port, A_neg(40) => 
                           negative_inputs_4_40_port, A_neg(39) => 
                           negative_inputs_4_39_port, A_neg(38) => 
                           negative_inputs_4_38_port, A_neg(37) => n108, 
                           A_neg(36) => negative_inputs_4_36_port, A_neg(35) =>
                           negative_inputs_4_35_port, A_neg(34) => 
                           negative_inputs_4_34_port, A_neg(33) => 
                           negative_inputs_4_33_port, A_neg(32) => 
                           negative_inputs_4_32_port, A_neg(31) => 
                           negative_inputs_4_31_port, A_neg(30) => 
                           negative_inputs_4_30_port, A_neg(29) => 
                           negative_inputs_4_29_port, A_neg(28) => 
                           negative_inputs_4_28_port, A_neg(27) => 
                           negative_inputs_4_27_port, A_neg(26) => 
                           negative_inputs_4_26_port, A_neg(25) => 
                           negative_inputs_4_25_port, A_neg(24) => 
                           negative_inputs_4_24_port, A_neg(23) => 
                           negative_inputs_4_23_port, A_neg(22) => 
                           negative_inputs_4_22_port, A_neg(21) => 
                           negative_inputs_4_21_port, A_neg(20) => 
                           negative_inputs_4_20_port, A_neg(19) => 
                           negative_inputs_4_19_port, A_neg(18) => 
                           negative_inputs_4_18_port, A_neg(17) => 
                           negative_inputs_4_17_port, A_neg(16) => 
                           negative_inputs_4_16_port, A_neg(15) => 
                           negative_inputs_4_15_port, A_neg(14) => 
                           negative_inputs_4_14_port, A_neg(13) => 
                           negative_inputs_4_13_port, A_neg(12) => 
                           negative_inputs_4_12_port, A_neg(11) => 
                           negative_inputs_4_11_port, A_neg(10) => 
                           negative_inputs_4_10_port, A_neg(9) => 
                           negative_inputs_4_9_port, A_neg(8) => 
                           negative_inputs_4_8_port, A_neg(7) => 
                           negative_inputs_4_7_port, A_neg(6) => 
                           negative_inputs_4_6_port, A_neg(5) => 
                           negative_inputs_4_5_port, A_neg(4) => 
                           negative_inputs_4_4_port, A_neg(3) => 
                           negative_inputs_4_3_port, A_neg(2) => 
                           negative_inputs_4_2_port, A_neg(1) => 
                           negative_inputs_4_1_port, A_neg(0) => n8, 
                           A_shifted(63) => positive_inputs_5_63_port, 
                           A_shifted(62) => positive_inputs_5_62_port, 
                           A_shifted(61) => positive_inputs_5_61_port, 
                           A_shifted(60) => positive_inputs_5_60_port, 
                           A_shifted(59) => positive_inputs_5_59_port, 
                           A_shifted(58) => positive_inputs_5_58_port, 
                           A_shifted(57) => positive_inputs_5_57_port, 
                           A_shifted(56) => positive_inputs_5_56_port, 
                           A_shifted(55) => positive_inputs_5_55_port, 
                           A_shifted(54) => positive_inputs_5_54_port, 
                           A_shifted(53) => positive_inputs_5_53_port, 
                           A_shifted(52) => positive_inputs_5_52_port, 
                           A_shifted(51) => positive_inputs_5_51_port, 
                           A_shifted(50) => positive_inputs_5_50_port, 
                           A_shifted(49) => positive_inputs_5_49_port, 
                           A_shifted(48) => positive_inputs_5_48_port, 
                           A_shifted(47) => n36, A_shifted(46) => 
                           positive_inputs_5_46_port, A_shifted(45) => 
                           positive_inputs_5_45_port, A_shifted(44) => 
                           positive_inputs_5_44_port, A_shifted(43) => 
                           positive_inputs_5_43_port, A_shifted(42) => 
                           positive_inputs_5_42_port, A_shifted(41) => 
                           positive_inputs_5_41_port, A_shifted(40) => 
                           positive_inputs_5_40_port, A_shifted(39) => 
                           positive_inputs_5_39_port, A_shifted(38) => 
                           positive_inputs_5_38_port, A_shifted(37) => n20, 
                           A_shifted(36) => n19, A_shifted(35) => n180, 
                           A_shifted(34) => n178, A_shifted(33) => n176, 
                           A_shifted(32) => n174, A_shifted(31) => n172, 
                           A_shifted(30) => n170, A_shifted(29) => n168, 
                           A_shifted(28) => n166, A_shifted(27) => n164, 
                           A_shifted(26) => n162, A_shifted(25) => n160, 
                           A_shifted(24) => n158, A_shifted(23) => n156, 
                           A_shifted(22) => n154, A_shifted(21) => n152, 
                           A_shifted(20) => n150, A_shifted(19) => n148, 
                           A_shifted(18) => n146, A_shifted(17) => n144, 
                           A_shifted(16) => n142, A_shifted(15) => n140, 
                           A_shifted(14) => n138, A_shifted(13) => n136, 
                           A_shifted(12) => n134, A_shifted(11) => n132, 
                           A_shifted(10) => n130, A_shifted(9) => n128, 
                           A_shifted(8) => n126, A_shifted(7) => n124, 
                           A_shifted(6) => n122, A_shifted(5) => n120, 
                           A_shifted(4) => positive_inputs_5_4_port, 
                           A_shifted(3) => positive_inputs_5_3_port, 
                           A_shifted(2) => positive_inputs_5_2_port, 
                           A_shifted(1) => positive_inputs_5_1_port, 
                           A_shifted(0) => n8, A_neg_shifted(63) => 
                           negative_inputs_5_63_port, A_neg_shifted(62) => 
                           negative_inputs_5_62_port, A_neg_shifted(61) => 
                           negative_inputs_5_61_port, A_neg_shifted(60) => 
                           negative_inputs_5_60_port, A_neg_shifted(59) => 
                           negative_inputs_5_59_port, A_neg_shifted(58) => 
                           negative_inputs_5_58_port, A_neg_shifted(57) => 
                           negative_inputs_5_57_port, A_neg_shifted(56) => 
                           negative_inputs_5_56_port, A_neg_shifted(55) => 
                           negative_inputs_5_55_port, A_neg_shifted(54) => 
                           negative_inputs_5_54_port, A_neg_shifted(53) => 
                           negative_inputs_5_53_port, A_neg_shifted(52) => 
                           negative_inputs_5_52_port, A_neg_shifted(51) => 
                           negative_inputs_5_51_port, A_neg_shifted(50) => 
                           negative_inputs_5_50_port, A_neg_shifted(49) => 
                           negative_inputs_5_49_port, A_neg_shifted(48) => 
                           negative_inputs_5_48_port, A_neg_shifted(47) => 
                           negative_inputs_5_47_port, A_neg_shifted(46) => 
                           negative_inputs_5_46_port, A_neg_shifted(45) => 
                           negative_inputs_5_45_port, A_neg_shifted(44) => 
                           negative_inputs_5_44_port, A_neg_shifted(43) => 
                           negative_inputs_5_43_port, A_neg_shifted(42) => 
                           negative_inputs_5_42_port, A_neg_shifted(41) => 
                           negative_inputs_5_41_port, A_neg_shifted(40) => 
                           negative_inputs_5_40_port, A_neg_shifted(39) => 
                           negative_inputs_5_39_port, A_neg_shifted(38) => 
                           negative_inputs_5_38_port, A_neg_shifted(37) => n106
                           , A_neg_shifted(36) => n104, A_neg_shifted(35) => 
                           n102, A_neg_shifted(34) => n100, A_neg_shifted(33) 
                           => n98, A_neg_shifted(32) => n96, A_neg_shifted(31) 
                           => n94, A_neg_shifted(30) => n92, A_neg_shifted(29) 
                           => n90, A_neg_shifted(28) => n88, A_neg_shifted(27) 
                           => n86, A_neg_shifted(26) => n84, A_neg_shifted(25) 
                           => n82, A_neg_shifted(24) => n80, A_neg_shifted(23) 
                           => n78, A_neg_shifted(22) => n76, A_neg_shifted(21) 
                           => n74, A_neg_shifted(20) => n72, A_neg_shifted(19) 
                           => n70, A_neg_shifted(18) => n68, A_neg_shifted(17) 
                           => n66, A_neg_shifted(16) => n64, A_neg_shifted(15) 
                           => n62, A_neg_shifted(14) => n60, A_neg_shifted(13) 
                           => n58, A_neg_shifted(12) => n56, A_neg_shifted(11) 
                           => n54, A_neg_shifted(10) => n52, A_neg_shifted(9) 
                           => n50, A_neg_shifted(8) => n48, A_neg_shifted(7) =>
                           n46, A_neg_shifted(6) => n44, A_neg_shifted(5) => 
                           n42, A_neg_shifted(4) => negative_inputs_5_4_port, 
                           A_neg_shifted(3) => negative_inputs_5_3_port, 
                           A_neg_shifted(2) => negative_inputs_5_2_port, 
                           A_neg_shifted(1) => negative_inputs_5_1_port, 
                           A_neg_shifted(0) => n8, Sel(2) => sel_2_2_port, 
                           Sel(1) => sel_2_1_port, Sel(0) => sel_2_0_port, 
                           Y(63) => MuxOutputs_2_63_port, Y(62) => 
                           MuxOutputs_2_62_port, Y(61) => MuxOutputs_2_61_port,
                           Y(60) => MuxOutputs_2_60_port, Y(59) => 
                           MuxOutputs_2_59_port, Y(58) => MuxOutputs_2_58_port,
                           Y(57) => MuxOutputs_2_57_port, Y(56) => 
                           MuxOutputs_2_56_port, Y(55) => MuxOutputs_2_55_port,
                           Y(54) => MuxOutputs_2_54_port, Y(53) => 
                           MuxOutputs_2_53_port, Y(52) => MuxOutputs_2_52_port,
                           Y(51) => MuxOutputs_2_51_port, Y(50) => 
                           MuxOutputs_2_50_port, Y(49) => MuxOutputs_2_49_port,
                           Y(48) => MuxOutputs_2_48_port, Y(47) => 
                           MuxOutputs_2_47_port, Y(46) => MuxOutputs_2_46_port,
                           Y(45) => MuxOutputs_2_45_port, Y(44) => 
                           MuxOutputs_2_44_port, Y(43) => MuxOutputs_2_43_port,
                           Y(42) => MuxOutputs_2_42_port, Y(41) => 
                           MuxOutputs_2_41_port, Y(40) => MuxOutputs_2_40_port,
                           Y(39) => MuxOutputs_2_39_port, Y(38) => 
                           MuxOutputs_2_38_port, Y(37) => MuxOutputs_2_37_port,
                           Y(36) => MuxOutputs_2_36_port, Y(35) => 
                           MuxOutputs_2_35_port, Y(34) => MuxOutputs_2_34_port,
                           Y(33) => MuxOutputs_2_33_port, Y(32) => 
                           MuxOutputs_2_32_port, Y(31) => MuxOutputs_2_31_port,
                           Y(30) => MuxOutputs_2_30_port, Y(29) => 
                           MuxOutputs_2_29_port, Y(28) => MuxOutputs_2_28_port,
                           Y(27) => MuxOutputs_2_27_port, Y(26) => 
                           MuxOutputs_2_26_port, Y(25) => MuxOutputs_2_25_port,
                           Y(24) => MuxOutputs_2_24_port, Y(23) => 
                           MuxOutputs_2_23_port, Y(22) => MuxOutputs_2_22_port,
                           Y(21) => MuxOutputs_2_21_port, Y(20) => 
                           MuxOutputs_2_20_port, Y(19) => MuxOutputs_2_19_port,
                           Y(18) => MuxOutputs_2_18_port, Y(17) => 
                           MuxOutputs_2_17_port, Y(16) => MuxOutputs_2_16_port,
                           Y(15) => MuxOutputs_2_15_port, Y(14) => 
                           MuxOutputs_2_14_port, Y(13) => MuxOutputs_2_13_port,
                           Y(12) => MuxOutputs_2_12_port, Y(11) => 
                           MuxOutputs_2_11_port, Y(10) => MuxOutputs_2_10_port,
                           Y(9) => MuxOutputs_2_9_port, Y(8) => 
                           MuxOutputs_2_8_port, Y(7) => MuxOutputs_2_7_port, 
                           Y(6) => MuxOutputs_2_6_port, Y(5) => 
                           MuxOutputs_2_5_port, Y(4) => MuxOutputs_2_4_port, 
                           Y(3) => MuxOutputs_2_3_port, Y(2) => 
                           MuxOutputs_2_2_port, Y(1) => MuxOutputs_2_1_port, 
                           Y(0) => MuxOutputs_2_0_port);
   encoderI_3 : encoder_29 port map( pieceofB(2) => B(7), pieceofB(1) => B(6), 
                           pieceofB(0) => B(5), sel(2) => sel_3_2_port, sel(1) 
                           => sel_3_1_port, sel(0) => sel_3_0_port);
   MUXI_3 : MUX51_MuxNbit64_29 port map( zeroSignal(63) => X_Logic0_port, 
                           zeroSignal(62) => X_Logic0_port, zeroSignal(61) => 
                           X_Logic0_port, zeroSignal(60) => X_Logic0_port, 
                           zeroSignal(59) => X_Logic0_port, zeroSignal(58) => 
                           X_Logic0_port, zeroSignal(57) => X_Logic0_port, 
                           zeroSignal(56) => X_Logic0_port, zeroSignal(55) => 
                           X_Logic0_port, zeroSignal(54) => X_Logic0_port, 
                           zeroSignal(53) => X_Logic0_port, zeroSignal(52) => 
                           X_Logic0_port, zeroSignal(51) => X_Logic0_port, 
                           zeroSignal(50) => X_Logic0_port, zeroSignal(49) => 
                           X_Logic0_port, zeroSignal(48) => X_Logic0_port, 
                           zeroSignal(47) => X_Logic0_port, zeroSignal(46) => 
                           X_Logic0_port, zeroSignal(45) => X_Logic0_port, 
                           zeroSignal(44) => X_Logic0_port, zeroSignal(43) => 
                           X_Logic0_port, zeroSignal(42) => X_Logic0_port, 
                           zeroSignal(41) => X_Logic0_port, zeroSignal(40) => 
                           X_Logic0_port, zeroSignal(39) => X_Logic0_port, 
                           zeroSignal(38) => X_Logic0_port, zeroSignal(37) => 
                           X_Logic0_port, zeroSignal(36) => X_Logic0_port, 
                           zeroSignal(35) => X_Logic0_port, zeroSignal(34) => 
                           X_Logic0_port, zeroSignal(33) => X_Logic0_port, 
                           zeroSignal(32) => X_Logic0_port, zeroSignal(31) => 
                           X_Logic0_port, zeroSignal(30) => X_Logic0_port, 
                           zeroSignal(29) => X_Logic0_port, zeroSignal(28) => 
                           X_Logic0_port, zeroSignal(27) => X_Logic0_port, 
                           zeroSignal(26) => X_Logic0_port, zeroSignal(25) => 
                           X_Logic0_port, zeroSignal(24) => X_Logic0_port, 
                           zeroSignal(23) => X_Logic0_port, zeroSignal(22) => 
                           X_Logic0_port, zeroSignal(21) => X_Logic0_port, 
                           zeroSignal(20) => X_Logic0_port, zeroSignal(19) => 
                           X_Logic0_port, zeroSignal(18) => X_Logic0_port, 
                           zeroSignal(17) => X_Logic0_port, zeroSignal(16) => 
                           X_Logic0_port, zeroSignal(15) => X_Logic0_port, 
                           zeroSignal(14) => X_Logic0_port, zeroSignal(13) => 
                           X_Logic0_port, zeroSignal(12) => X_Logic0_port, 
                           zeroSignal(11) => X_Logic0_port, zeroSignal(10) => 
                           X_Logic0_port, zeroSignal(9) => X_Logic0_port, 
                           zeroSignal(8) => X_Logic0_port, zeroSignal(7) => 
                           X_Logic0_port, zeroSignal(6) => X_Logic0_port, 
                           zeroSignal(5) => X_Logic0_port, zeroSignal(4) => 
                           X_Logic0_port, zeroSignal(3) => X_Logic0_port, 
                           zeroSignal(2) => X_Logic0_port, zeroSignal(1) => 
                           X_Logic0_port, zeroSignal(0) => X_Logic0_port, 
                           A_signal(63) => positive_inputs_6_63_port, 
                           A_signal(62) => positive_inputs_6_62_port, 
                           A_signal(61) => positive_inputs_6_61_port, 
                           A_signal(60) => positive_inputs_6_60_port, 
                           A_signal(59) => positive_inputs_6_59_port, 
                           A_signal(58) => positive_inputs_6_58_port, 
                           A_signal(57) => positive_inputs_6_57_port, 
                           A_signal(56) => positive_inputs_6_56_port, 
                           A_signal(55) => positive_inputs_6_55_port, 
                           A_signal(54) => positive_inputs_6_54_port, 
                           A_signal(53) => positive_inputs_6_53_port, 
                           A_signal(52) => positive_inputs_6_52_port, 
                           A_signal(51) => positive_inputs_6_51_port, 
                           A_signal(50) => positive_inputs_6_50_port, 
                           A_signal(49) => positive_inputs_6_49_port, 
                           A_signal(48) => positive_inputs_6_48_port, 
                           A_signal(47) => n35, A_signal(46) => 
                           positive_inputs_6_46_port, A_signal(45) => 
                           positive_inputs_6_45_port, A_signal(44) => 
                           positive_inputs_6_44_port, A_signal(43) => 
                           positive_inputs_6_43_port, A_signal(42) => 
                           positive_inputs_6_42_port, A_signal(41) => 
                           positive_inputs_6_41_port, A_signal(40) => 
                           positive_inputs_6_40_port, A_signal(39) => 
                           positive_inputs_6_39_port, A_signal(38) => 
                           positive_inputs_6_38_port, A_signal(37) => 
                           positive_inputs_6_37_port, A_signal(36) => 
                           positive_inputs_6_36_port, A_signal(35) => 
                           positive_inputs_6_35_port, A_signal(34) => 
                           positive_inputs_6_34_port, A_signal(33) => 
                           positive_inputs_6_33_port, A_signal(32) => 
                           positive_inputs_6_32_port, A_signal(31) => 
                           positive_inputs_6_31_port, A_signal(30) => 
                           positive_inputs_6_30_port, A_signal(29) => 
                           positive_inputs_6_29_port, A_signal(28) => 
                           positive_inputs_6_28_port, A_signal(27) => 
                           positive_inputs_6_27_port, A_signal(26) => 
                           positive_inputs_6_26_port, A_signal(25) => 
                           positive_inputs_6_25_port, A_signal(24) => 
                           positive_inputs_6_24_port, A_signal(23) => 
                           positive_inputs_6_23_port, A_signal(22) => 
                           positive_inputs_6_22_port, A_signal(21) => 
                           positive_inputs_6_21_port, A_signal(20) => 
                           positive_inputs_6_20_port, A_signal(19) => 
                           positive_inputs_6_19_port, A_signal(18) => 
                           positive_inputs_6_18_port, A_signal(17) => 
                           positive_inputs_6_17_port, A_signal(16) => 
                           positive_inputs_6_16_port, A_signal(15) => 
                           positive_inputs_6_15_port, A_signal(14) => 
                           positive_inputs_6_14_port, A_signal(13) => 
                           positive_inputs_6_13_port, A_signal(12) => 
                           positive_inputs_6_12_port, A_signal(11) => 
                           positive_inputs_6_11_port, A_signal(10) => 
                           positive_inputs_6_10_port, A_signal(9) => 
                           positive_inputs_6_9_port, A_signal(8) => 
                           positive_inputs_6_8_port, A_signal(7) => 
                           positive_inputs_6_7_port, A_signal(6) => 
                           positive_inputs_6_6_port, A_signal(5) => 
                           positive_inputs_6_5_port, A_signal(4) => 
                           positive_inputs_6_4_port, A_signal(3) => 
                           positive_inputs_6_3_port, A_signal(2) => 
                           positive_inputs_6_2_port, A_signal(1) => 
                           positive_inputs_6_1_port, A_signal(0) => n8, 
                           A_neg(63) => negative_inputs_6_63_port, A_neg(62) =>
                           negative_inputs_6_62_port, A_neg(61) => 
                           negative_inputs_6_61_port, A_neg(60) => 
                           negative_inputs_6_60_port, A_neg(59) => 
                           negative_inputs_6_59_port, A_neg(58) => 
                           negative_inputs_6_58_port, A_neg(57) => 
                           negative_inputs_6_57_port, A_neg(56) => 
                           negative_inputs_6_56_port, A_neg(55) => 
                           negative_inputs_6_55_port, A_neg(54) => 
                           negative_inputs_6_54_port, A_neg(53) => 
                           negative_inputs_6_53_port, A_neg(52) => 
                           negative_inputs_6_52_port, A_neg(51) => 
                           negative_inputs_6_51_port, A_neg(50) => 
                           negative_inputs_6_50_port, A_neg(49) => 
                           negative_inputs_6_49_port, A_neg(48) => 
                           negative_inputs_6_48_port, A_neg(47) => 
                           negative_inputs_6_47_port, A_neg(46) => 
                           negative_inputs_6_46_port, A_neg(45) => 
                           negative_inputs_6_45_port, A_neg(44) => 
                           negative_inputs_6_44_port, A_neg(43) => 
                           negative_inputs_6_43_port, A_neg(42) => 
                           negative_inputs_6_42_port, A_neg(41) => 
                           negative_inputs_6_41_port, A_neg(40) => 
                           negative_inputs_6_40_port, A_neg(39) => 
                           negative_inputs_6_39_port, A_neg(38) => 
                           negative_inputs_6_38_port, A_neg(37) => 
                           negative_inputs_6_37_port, A_neg(36) => 
                           negative_inputs_6_36_port, A_neg(35) => 
                           negative_inputs_6_35_port, A_neg(34) => 
                           negative_inputs_6_34_port, A_neg(33) => 
                           negative_inputs_6_33_port, A_neg(32) => 
                           negative_inputs_6_32_port, A_neg(31) => 
                           negative_inputs_6_31_port, A_neg(30) => 
                           negative_inputs_6_30_port, A_neg(29) => 
                           negative_inputs_6_29_port, A_neg(28) => 
                           negative_inputs_6_28_port, A_neg(27) => 
                           negative_inputs_6_27_port, A_neg(26) => 
                           negative_inputs_6_26_port, A_neg(25) => 
                           negative_inputs_6_25_port, A_neg(24) => 
                           negative_inputs_6_24_port, A_neg(23) => 
                           negative_inputs_6_23_port, A_neg(22) => 
                           negative_inputs_6_22_port, A_neg(21) => 
                           negative_inputs_6_21_port, A_neg(20) => 
                           negative_inputs_6_20_port, A_neg(19) => 
                           negative_inputs_6_19_port, A_neg(18) => 
                           negative_inputs_6_18_port, A_neg(17) => 
                           negative_inputs_6_17_port, A_neg(16) => 
                           negative_inputs_6_16_port, A_neg(15) => 
                           negative_inputs_6_15_port, A_neg(14) => 
                           negative_inputs_6_14_port, A_neg(13) => 
                           negative_inputs_6_13_port, A_neg(12) => 
                           negative_inputs_6_12_port, A_neg(11) => 
                           negative_inputs_6_11_port, A_neg(10) => 
                           negative_inputs_6_10_port, A_neg(9) => 
                           negative_inputs_6_9_port, A_neg(8) => 
                           negative_inputs_6_8_port, A_neg(7) => 
                           negative_inputs_6_7_port, A_neg(6) => 
                           negative_inputs_6_6_port, A_neg(5) => 
                           negative_inputs_6_5_port, A_neg(4) => 
                           negative_inputs_6_4_port, A_neg(3) => 
                           negative_inputs_6_3_port, A_neg(2) => 
                           negative_inputs_6_2_port, A_neg(1) => 
                           negative_inputs_6_1_port, A_neg(0) => n8, 
                           A_shifted(63) => positive_inputs_7_63_port, 
                           A_shifted(62) => positive_inputs_7_62_port, 
                           A_shifted(61) => positive_inputs_7_61_port, 
                           A_shifted(60) => positive_inputs_7_60_port, 
                           A_shifted(59) => positive_inputs_7_59_port, 
                           A_shifted(58) => positive_inputs_7_58_port, 
                           A_shifted(57) => positive_inputs_7_57_port, 
                           A_shifted(56) => positive_inputs_7_56_port, 
                           A_shifted(55) => positive_inputs_7_55_port, 
                           A_shifted(54) => positive_inputs_7_54_port, 
                           A_shifted(53) => positive_inputs_7_53_port, 
                           A_shifted(52) => positive_inputs_7_52_port, 
                           A_shifted(51) => positive_inputs_7_51_port, 
                           A_shifted(50) => positive_inputs_7_50_port, 
                           A_shifted(49) => positive_inputs_7_49_port, 
                           A_shifted(48) => positive_inputs_7_48_port, 
                           A_shifted(47) => n34, A_shifted(46) => 
                           positive_inputs_7_46_port, A_shifted(45) => 
                           positive_inputs_7_45_port, A_shifted(44) => 
                           positive_inputs_7_44_port, A_shifted(43) => 
                           positive_inputs_7_43_port, A_shifted(42) => 
                           positive_inputs_7_42_port, A_shifted(41) => 
                           positive_inputs_7_41_port, A_shifted(40) => 
                           positive_inputs_7_40_port, A_shifted(39) => 
                           positive_inputs_7_39_port, A_shifted(38) => 
                           positive_inputs_7_38_port, A_shifted(37) => 
                           positive_inputs_7_37_port, A_shifted(36) => 
                           positive_inputs_7_36_port, A_shifted(35) => 
                           positive_inputs_7_35_port, A_shifted(34) => 
                           positive_inputs_7_34_port, A_shifted(33) => 
                           positive_inputs_7_33_port, A_shifted(32) => 
                           positive_inputs_7_32_port, A_shifted(31) => 
                           positive_inputs_7_31_port, A_shifted(30) => 
                           positive_inputs_7_30_port, A_shifted(29) => 
                           positive_inputs_7_29_port, A_shifted(28) => 
                           positive_inputs_7_28_port, A_shifted(27) => 
                           positive_inputs_7_27_port, A_shifted(26) => 
                           positive_inputs_7_26_port, A_shifted(25) => 
                           positive_inputs_7_25_port, A_shifted(24) => 
                           positive_inputs_7_24_port, A_shifted(23) => 
                           positive_inputs_7_23_port, A_shifted(22) => 
                           positive_inputs_7_22_port, A_shifted(21) => 
                           positive_inputs_7_21_port, A_shifted(20) => 
                           positive_inputs_7_20_port, A_shifted(19) => 
                           positive_inputs_7_19_port, A_shifted(18) => 
                           positive_inputs_7_18_port, A_shifted(17) => 
                           positive_inputs_7_17_port, A_shifted(16) => 
                           positive_inputs_7_16_port, A_shifted(15) => 
                           positive_inputs_7_15_port, A_shifted(14) => 
                           positive_inputs_7_14_port, A_shifted(13) => 
                           positive_inputs_7_13_port, A_shifted(12) => 
                           positive_inputs_7_12_port, A_shifted(11) => 
                           positive_inputs_7_11_port, A_shifted(10) => 
                           positive_inputs_7_10_port, A_shifted(9) => 
                           positive_inputs_7_9_port, A_shifted(8) => 
                           positive_inputs_7_8_port, A_shifted(7) => 
                           positive_inputs_7_7_port, A_shifted(6) => 
                           positive_inputs_7_6_port, A_shifted(5) => 
                           positive_inputs_7_5_port, A_shifted(4) => 
                           positive_inputs_7_4_port, A_shifted(3) => 
                           positive_inputs_7_3_port, A_shifted(2) => 
                           positive_inputs_7_2_port, A_shifted(1) => 
                           positive_inputs_7_1_port, A_shifted(0) => n8, 
                           A_neg_shifted(63) => negative_inputs_7_63_port, 
                           A_neg_shifted(62) => negative_inputs_7_62_port, 
                           A_neg_shifted(61) => negative_inputs_7_61_port, 
                           A_neg_shifted(60) => negative_inputs_7_60_port, 
                           A_neg_shifted(59) => negative_inputs_7_59_port, 
                           A_neg_shifted(58) => negative_inputs_7_58_port, 
                           A_neg_shifted(57) => negative_inputs_7_57_port, 
                           A_neg_shifted(56) => negative_inputs_7_56_port, 
                           A_neg_shifted(55) => negative_inputs_7_55_port, 
                           A_neg_shifted(54) => negative_inputs_7_54_port, 
                           A_neg_shifted(53) => negative_inputs_7_53_port, 
                           A_neg_shifted(52) => negative_inputs_7_52_port, 
                           A_neg_shifted(51) => negative_inputs_7_51_port, 
                           A_neg_shifted(50) => negative_inputs_7_50_port, 
                           A_neg_shifted(49) => negative_inputs_7_49_port, 
                           A_neg_shifted(48) => negative_inputs_7_48_port, 
                           A_neg_shifted(47) => n119, A_neg_shifted(46) => 
                           negative_inputs_7_46_port, A_neg_shifted(45) => 
                           negative_inputs_7_45_port, A_neg_shifted(44) => 
                           negative_inputs_7_44_port, A_neg_shifted(43) => 
                           negative_inputs_7_43_port, A_neg_shifted(42) => 
                           negative_inputs_7_42_port, A_neg_shifted(41) => 
                           negative_inputs_7_41_port, A_neg_shifted(40) => 
                           negative_inputs_7_40_port, A_neg_shifted(39) => 
                           negative_inputs_7_39_port, A_neg_shifted(38) => 
                           negative_inputs_7_38_port, A_neg_shifted(37) => 
                           negative_inputs_7_37_port, A_neg_shifted(36) => 
                           negative_inputs_7_36_port, A_neg_shifted(35) => 
                           negative_inputs_7_35_port, A_neg_shifted(34) => 
                           negative_inputs_7_34_port, A_neg_shifted(33) => 
                           negative_inputs_7_33_port, A_neg_shifted(32) => 
                           negative_inputs_7_32_port, A_neg_shifted(31) => 
                           negative_inputs_7_31_port, A_neg_shifted(30) => 
                           negative_inputs_7_30_port, A_neg_shifted(29) => 
                           negative_inputs_7_29_port, A_neg_shifted(28) => 
                           negative_inputs_7_28_port, A_neg_shifted(27) => 
                           negative_inputs_7_27_port, A_neg_shifted(26) => 
                           negative_inputs_7_26_port, A_neg_shifted(25) => 
                           negative_inputs_7_25_port, A_neg_shifted(24) => 
                           negative_inputs_7_24_port, A_neg_shifted(23) => 
                           negative_inputs_7_23_port, A_neg_shifted(22) => 
                           negative_inputs_7_22_port, A_neg_shifted(21) => 
                           negative_inputs_7_21_port, A_neg_shifted(20) => 
                           negative_inputs_7_20_port, A_neg_shifted(19) => 
                           negative_inputs_7_19_port, A_neg_shifted(18) => 
                           negative_inputs_7_18_port, A_neg_shifted(17) => 
                           negative_inputs_7_17_port, A_neg_shifted(16) => 
                           negative_inputs_7_16_port, A_neg_shifted(15) => 
                           negative_inputs_7_15_port, A_neg_shifted(14) => 
                           negative_inputs_7_14_port, A_neg_shifted(13) => 
                           negative_inputs_7_13_port, A_neg_shifted(12) => 
                           negative_inputs_7_12_port, A_neg_shifted(11) => 
                           negative_inputs_7_11_port, A_neg_shifted(10) => 
                           negative_inputs_7_10_port, A_neg_shifted(9) => 
                           negative_inputs_7_9_port, A_neg_shifted(8) => 
                           negative_inputs_7_8_port, A_neg_shifted(7) => 
                           negative_inputs_7_7_port, A_neg_shifted(6) => 
                           negative_inputs_7_6_port, A_neg_shifted(5) => 
                           negative_inputs_7_5_port, A_neg_shifted(4) => 
                           negative_inputs_7_4_port, A_neg_shifted(3) => 
                           negative_inputs_7_3_port, A_neg_shifted(2) => 
                           negative_inputs_7_2_port, A_neg_shifted(1) => 
                           negative_inputs_7_1_port, A_neg_shifted(0) => n8, 
                           Sel(2) => sel_3_2_port, Sel(1) => sel_3_1_port, 
                           Sel(0) => sel_3_0_port, Y(63) => 
                           MuxOutputs_3_63_port, Y(62) => MuxOutputs_3_62_port,
                           Y(61) => MuxOutputs_3_61_port, Y(60) => 
                           MuxOutputs_3_60_port, Y(59) => MuxOutputs_3_59_port,
                           Y(58) => MuxOutputs_3_58_port, Y(57) => 
                           MuxOutputs_3_57_port, Y(56) => MuxOutputs_3_56_port,
                           Y(55) => MuxOutputs_3_55_port, Y(54) => 
                           MuxOutputs_3_54_port, Y(53) => MuxOutputs_3_53_port,
                           Y(52) => MuxOutputs_3_52_port, Y(51) => 
                           MuxOutputs_3_51_port, Y(50) => MuxOutputs_3_50_port,
                           Y(49) => MuxOutputs_3_49_port, Y(48) => 
                           MuxOutputs_3_48_port, Y(47) => MuxOutputs_3_47_port,
                           Y(46) => MuxOutputs_3_46_port, Y(45) => 
                           MuxOutputs_3_45_port, Y(44) => MuxOutputs_3_44_port,
                           Y(43) => MuxOutputs_3_43_port, Y(42) => 
                           MuxOutputs_3_42_port, Y(41) => MuxOutputs_3_41_port,
                           Y(40) => MuxOutputs_3_40_port, Y(39) => 
                           MuxOutputs_3_39_port, Y(38) => MuxOutputs_3_38_port,
                           Y(37) => MuxOutputs_3_37_port, Y(36) => 
                           MuxOutputs_3_36_port, Y(35) => MuxOutputs_3_35_port,
                           Y(34) => MuxOutputs_3_34_port, Y(33) => 
                           MuxOutputs_3_33_port, Y(32) => MuxOutputs_3_32_port,
                           Y(31) => MuxOutputs_3_31_port, Y(30) => 
                           MuxOutputs_3_30_port, Y(29) => MuxOutputs_3_29_port,
                           Y(28) => MuxOutputs_3_28_port, Y(27) => 
                           MuxOutputs_3_27_port, Y(26) => MuxOutputs_3_26_port,
                           Y(25) => MuxOutputs_3_25_port, Y(24) => 
                           MuxOutputs_3_24_port, Y(23) => MuxOutputs_3_23_port,
                           Y(22) => MuxOutputs_3_22_port, Y(21) => 
                           MuxOutputs_3_21_port, Y(20) => MuxOutputs_3_20_port,
                           Y(19) => MuxOutputs_3_19_port, Y(18) => 
                           MuxOutputs_3_18_port, Y(17) => MuxOutputs_3_17_port,
                           Y(16) => MuxOutputs_3_16_port, Y(15) => 
                           MuxOutputs_3_15_port, Y(14) => MuxOutputs_3_14_port,
                           Y(13) => MuxOutputs_3_13_port, Y(12) => 
                           MuxOutputs_3_12_port, Y(11) => MuxOutputs_3_11_port,
                           Y(10) => MuxOutputs_3_10_port, Y(9) => 
                           MuxOutputs_3_9_port, Y(8) => MuxOutputs_3_8_port, 
                           Y(7) => MuxOutputs_3_7_port, Y(6) => 
                           MuxOutputs_3_6_port, Y(5) => MuxOutputs_3_5_port, 
                           Y(4) => MuxOutputs_3_4_port, Y(3) => 
                           MuxOutputs_3_3_port, Y(2) => MuxOutputs_3_2_port, 
                           Y(1) => MuxOutputs_3_1_port, Y(0) => 
                           MuxOutputs_3_0_port);
   encoderI_4 : encoder_28 port map( pieceofB(2) => B(9), pieceofB(1) => B(8), 
                           pieceofB(0) => B(7), sel(2) => sel_4_2_port, sel(1) 
                           => sel_4_1_port, sel(0) => sel_4_0_port);
   MUXI_4 : MUX51_MuxNbit64_28 port map( zeroSignal(63) => X_Logic0_port, 
                           zeroSignal(62) => X_Logic0_port, zeroSignal(61) => 
                           X_Logic0_port, zeroSignal(60) => X_Logic0_port, 
                           zeroSignal(59) => X_Logic0_port, zeroSignal(58) => 
                           X_Logic0_port, zeroSignal(57) => X_Logic0_port, 
                           zeroSignal(56) => X_Logic0_port, zeroSignal(55) => 
                           X_Logic0_port, zeroSignal(54) => X_Logic0_port, 
                           zeroSignal(53) => X_Logic0_port, zeroSignal(52) => 
                           X_Logic0_port, zeroSignal(51) => X_Logic0_port, 
                           zeroSignal(50) => X_Logic0_port, zeroSignal(49) => 
                           X_Logic0_port, zeroSignal(48) => X_Logic0_port, 
                           zeroSignal(47) => X_Logic0_port, zeroSignal(46) => 
                           X_Logic0_port, zeroSignal(45) => X_Logic0_port, 
                           zeroSignal(44) => X_Logic0_port, zeroSignal(43) => 
                           X_Logic0_port, zeroSignal(42) => X_Logic0_port, 
                           zeroSignal(41) => X_Logic0_port, zeroSignal(40) => 
                           X_Logic0_port, zeroSignal(39) => X_Logic0_port, 
                           zeroSignal(38) => X_Logic0_port, zeroSignal(37) => 
                           X_Logic0_port, zeroSignal(36) => X_Logic0_port, 
                           zeroSignal(35) => X_Logic0_port, zeroSignal(34) => 
                           X_Logic0_port, zeroSignal(33) => X_Logic0_port, 
                           zeroSignal(32) => X_Logic0_port, zeroSignal(31) => 
                           X_Logic0_port, zeroSignal(30) => X_Logic0_port, 
                           zeroSignal(29) => X_Logic0_port, zeroSignal(28) => 
                           X_Logic0_port, zeroSignal(27) => X_Logic0_port, 
                           zeroSignal(26) => X_Logic0_port, zeroSignal(25) => 
                           X_Logic0_port, zeroSignal(24) => X_Logic0_port, 
                           zeroSignal(23) => X_Logic0_port, zeroSignal(22) => 
                           X_Logic0_port, zeroSignal(21) => X_Logic0_port, 
                           zeroSignal(20) => X_Logic0_port, zeroSignal(19) => 
                           X_Logic0_port, zeroSignal(18) => X_Logic0_port, 
                           zeroSignal(17) => X_Logic0_port, zeroSignal(16) => 
                           X_Logic0_port, zeroSignal(15) => X_Logic0_port, 
                           zeroSignal(14) => X_Logic0_port, zeroSignal(13) => 
                           X_Logic0_port, zeroSignal(12) => X_Logic0_port, 
                           zeroSignal(11) => X_Logic0_port, zeroSignal(10) => 
                           X_Logic0_port, zeroSignal(9) => X_Logic0_port, 
                           zeroSignal(8) => X_Logic0_port, zeroSignal(7) => 
                           X_Logic0_port, zeroSignal(6) => X_Logic0_port, 
                           zeroSignal(5) => X_Logic0_port, zeroSignal(4) => 
                           X_Logic0_port, zeroSignal(3) => X_Logic0_port, 
                           zeroSignal(2) => X_Logic0_port, zeroSignal(1) => 
                           X_Logic0_port, zeroSignal(0) => X_Logic0_port, 
                           A_signal(63) => positive_inputs_8_63_port, 
                           A_signal(62) => positive_inputs_8_62_port, 
                           A_signal(61) => positive_inputs_8_61_port, 
                           A_signal(60) => positive_inputs_8_60_port, 
                           A_signal(59) => positive_inputs_8_59_port, 
                           A_signal(58) => positive_inputs_8_58_port, 
                           A_signal(57) => positive_inputs_8_57_port, 
                           A_signal(56) => positive_inputs_8_56_port, 
                           A_signal(55) => positive_inputs_8_55_port, 
                           A_signal(54) => positive_inputs_8_54_port, 
                           A_signal(53) => positive_inputs_8_53_port, 
                           A_signal(52) => positive_inputs_8_52_port, 
                           A_signal(51) => positive_inputs_8_51_port, 
                           A_signal(50) => positive_inputs_8_50_port, 
                           A_signal(49) => positive_inputs_8_49_port, 
                           A_signal(48) => positive_inputs_8_48_port, 
                           A_signal(47) => n33, A_signal(46) => 
                           positive_inputs_8_46_port, A_signal(45) => 
                           positive_inputs_8_45_port, A_signal(44) => 
                           positive_inputs_8_44_port, A_signal(43) => 
                           positive_inputs_8_43_port, A_signal(42) => 
                           positive_inputs_8_42_port, A_signal(41) => 
                           positive_inputs_8_41_port, A_signal(40) => 
                           positive_inputs_8_40_port, A_signal(39) => 
                           positive_inputs_8_39_port, A_signal(38) => 
                           positive_inputs_8_38_port, A_signal(37) => 
                           positive_inputs_8_37_port, A_signal(36) => 
                           positive_inputs_8_36_port, A_signal(35) => 
                           positive_inputs_8_35_port, A_signal(34) => 
                           positive_inputs_8_34_port, A_signal(33) => 
                           positive_inputs_8_33_port, A_signal(32) => 
                           positive_inputs_8_32_port, A_signal(31) => 
                           positive_inputs_8_31_port, A_signal(30) => 
                           positive_inputs_8_30_port, A_signal(29) => 
                           positive_inputs_8_29_port, A_signal(28) => 
                           positive_inputs_8_28_port, A_signal(27) => 
                           positive_inputs_8_27_port, A_signal(26) => 
                           positive_inputs_8_26_port, A_signal(25) => 
                           positive_inputs_8_25_port, A_signal(24) => 
                           positive_inputs_8_24_port, A_signal(23) => 
                           positive_inputs_8_23_port, A_signal(22) => 
                           positive_inputs_8_22_port, A_signal(21) => 
                           positive_inputs_8_21_port, A_signal(20) => 
                           positive_inputs_8_20_port, A_signal(19) => 
                           positive_inputs_8_19_port, A_signal(18) => 
                           positive_inputs_8_18_port, A_signal(17) => 
                           positive_inputs_8_17_port, A_signal(16) => 
                           positive_inputs_8_16_port, A_signal(15) => 
                           positive_inputs_8_15_port, A_signal(14) => 
                           positive_inputs_8_14_port, A_signal(13) => 
                           positive_inputs_8_13_port, A_signal(12) => 
                           positive_inputs_8_12_port, A_signal(11) => 
                           positive_inputs_8_11_port, A_signal(10) => 
                           positive_inputs_8_10_port, A_signal(9) => 
                           positive_inputs_8_9_port, A_signal(8) => 
                           positive_inputs_8_8_port, A_signal(7) => 
                           positive_inputs_8_7_port, A_signal(6) => 
                           positive_inputs_8_6_port, A_signal(5) => 
                           positive_inputs_8_5_port, A_signal(4) => 
                           positive_inputs_8_4_port, A_signal(3) => 
                           positive_inputs_8_3_port, A_signal(2) => 
                           positive_inputs_8_2_port, A_signal(1) => 
                           positive_inputs_8_1_port, A_signal(0) => n8, 
                           A_neg(63) => negative_inputs_8_63_port, A_neg(62) =>
                           negative_inputs_8_62_port, A_neg(61) => 
                           negative_inputs_8_61_port, A_neg(60) => 
                           negative_inputs_8_60_port, A_neg(59) => 
                           negative_inputs_8_59_port, A_neg(58) => 
                           negative_inputs_8_58_port, A_neg(57) => 
                           negative_inputs_8_57_port, A_neg(56) => 
                           negative_inputs_8_56_port, A_neg(55) => 
                           negative_inputs_8_55_port, A_neg(54) => 
                           negative_inputs_8_54_port, A_neg(53) => 
                           negative_inputs_8_53_port, A_neg(52) => 
                           negative_inputs_8_52_port, A_neg(51) => 
                           negative_inputs_8_51_port, A_neg(50) => 
                           negative_inputs_8_50_port, A_neg(49) => 
                           negative_inputs_8_49_port, A_neg(48) => 
                           negative_inputs_8_48_port, A_neg(47) => n118, 
                           A_neg(46) => negative_inputs_8_46_port, A_neg(45) =>
                           negative_inputs_8_45_port, A_neg(44) => 
                           negative_inputs_8_44_port, A_neg(43) => 
                           negative_inputs_8_43_port, A_neg(42) => 
                           negative_inputs_8_42_port, A_neg(41) => 
                           negative_inputs_8_41_port, A_neg(40) => 
                           negative_inputs_8_40_port, A_neg(39) => 
                           negative_inputs_8_39_port, A_neg(38) => 
                           negative_inputs_8_38_port, A_neg(37) => 
                           negative_inputs_8_37_port, A_neg(36) => 
                           negative_inputs_8_36_port, A_neg(35) => 
                           negative_inputs_8_35_port, A_neg(34) => 
                           negative_inputs_8_34_port, A_neg(33) => 
                           negative_inputs_8_33_port, A_neg(32) => 
                           negative_inputs_8_32_port, A_neg(31) => 
                           negative_inputs_8_31_port, A_neg(30) => 
                           negative_inputs_8_30_port, A_neg(29) => 
                           negative_inputs_8_29_port, A_neg(28) => 
                           negative_inputs_8_28_port, A_neg(27) => 
                           negative_inputs_8_27_port, A_neg(26) => 
                           negative_inputs_8_26_port, A_neg(25) => 
                           negative_inputs_8_25_port, A_neg(24) => 
                           negative_inputs_8_24_port, A_neg(23) => 
                           negative_inputs_8_23_port, A_neg(22) => 
                           negative_inputs_8_22_port, A_neg(21) => 
                           negative_inputs_8_21_port, A_neg(20) => 
                           negative_inputs_8_20_port, A_neg(19) => 
                           negative_inputs_8_19_port, A_neg(18) => 
                           negative_inputs_8_18_port, A_neg(17) => 
                           negative_inputs_8_17_port, A_neg(16) => 
                           negative_inputs_8_16_port, A_neg(15) => 
                           negative_inputs_8_15_port, A_neg(14) => 
                           negative_inputs_8_14_port, A_neg(13) => 
                           negative_inputs_8_13_port, A_neg(12) => 
                           negative_inputs_8_12_port, A_neg(11) => 
                           negative_inputs_8_11_port, A_neg(10) => 
                           negative_inputs_8_10_port, A_neg(9) => 
                           negative_inputs_8_9_port, A_neg(8) => 
                           negative_inputs_8_8_port, A_neg(7) => 
                           negative_inputs_8_7_port, A_neg(6) => 
                           negative_inputs_8_6_port, A_neg(5) => 
                           negative_inputs_8_5_port, A_neg(4) => 
                           negative_inputs_8_4_port, A_neg(3) => 
                           negative_inputs_8_3_port, A_neg(2) => 
                           negative_inputs_8_2_port, A_neg(1) => 
                           negative_inputs_8_1_port, A_neg(0) => n8, 
                           A_shifted(63) => positive_inputs_9_63_port, 
                           A_shifted(62) => positive_inputs_9_62_port, 
                           A_shifted(61) => positive_inputs_9_61_port, 
                           A_shifted(60) => positive_inputs_9_60_port, 
                           A_shifted(59) => positive_inputs_9_59_port, 
                           A_shifted(58) => positive_inputs_9_58_port, 
                           A_shifted(57) => positive_inputs_9_57_port, 
                           A_shifted(56) => positive_inputs_9_56_port, 
                           A_shifted(55) => positive_inputs_9_55_port, 
                           A_shifted(54) => positive_inputs_9_54_port, 
                           A_shifted(53) => positive_inputs_9_53_port, 
                           A_shifted(52) => positive_inputs_9_52_port, 
                           A_shifted(51) => positive_inputs_9_51_port, 
                           A_shifted(50) => positive_inputs_9_50_port, 
                           A_shifted(49) => positive_inputs_9_49_port, 
                           A_shifted(48) => positive_inputs_9_48_port, 
                           A_shifted(47) => n32, A_shifted(46) => 
                           positive_inputs_9_46_port, A_shifted(45) => 
                           positive_inputs_9_45_port, A_shifted(44) => 
                           positive_inputs_9_44_port, A_shifted(43) => 
                           positive_inputs_9_43_port, A_shifted(42) => 
                           positive_inputs_9_42_port, A_shifted(41) => 
                           positive_inputs_9_41_port, A_shifted(40) => 
                           positive_inputs_9_40_port, A_shifted(39) => 
                           positive_inputs_9_39_port, A_shifted(38) => 
                           positive_inputs_9_38_port, A_shifted(37) => 
                           positive_inputs_9_37_port, A_shifted(36) => 
                           positive_inputs_9_36_port, A_shifted(35) => 
                           positive_inputs_9_35_port, A_shifted(34) => 
                           positive_inputs_9_34_port, A_shifted(33) => 
                           positive_inputs_9_33_port, A_shifted(32) => 
                           positive_inputs_9_32_port, A_shifted(31) => 
                           positive_inputs_9_31_port, A_shifted(30) => 
                           positive_inputs_9_30_port, A_shifted(29) => 
                           positive_inputs_9_29_port, A_shifted(28) => 
                           positive_inputs_9_28_port, A_shifted(27) => 
                           positive_inputs_9_27_port, A_shifted(26) => 
                           positive_inputs_9_26_port, A_shifted(25) => 
                           positive_inputs_9_25_port, A_shifted(24) => 
                           positive_inputs_9_24_port, A_shifted(23) => 
                           positive_inputs_9_23_port, A_shifted(22) => 
                           positive_inputs_9_22_port, A_shifted(21) => 
                           positive_inputs_9_21_port, A_shifted(20) => 
                           positive_inputs_9_20_port, A_shifted(19) => 
                           positive_inputs_9_19_port, A_shifted(18) => 
                           positive_inputs_9_18_port, A_shifted(17) => 
                           positive_inputs_9_17_port, A_shifted(16) => 
                           positive_inputs_9_16_port, A_shifted(15) => 
                           positive_inputs_9_15_port, A_shifted(14) => 
                           positive_inputs_9_14_port, A_shifted(13) => 
                           positive_inputs_9_13_port, A_shifted(12) => 
                           positive_inputs_9_12_port, A_shifted(11) => 
                           positive_inputs_9_11_port, A_shifted(10) => 
                           positive_inputs_9_10_port, A_shifted(9) => 
                           positive_inputs_9_9_port, A_shifted(8) => 
                           positive_inputs_9_8_port, A_shifted(7) => 
                           positive_inputs_9_7_port, A_shifted(6) => 
                           positive_inputs_9_6_port, A_shifted(5) => 
                           positive_inputs_9_5_port, A_shifted(4) => 
                           positive_inputs_9_4_port, A_shifted(3) => 
                           positive_inputs_9_3_port, A_shifted(2) => 
                           positive_inputs_9_2_port, A_shifted(1) => 
                           positive_inputs_9_1_port, A_shifted(0) => n8, 
                           A_neg_shifted(63) => negative_inputs_9_63_port, 
                           A_neg_shifted(62) => negative_inputs_9_62_port, 
                           A_neg_shifted(61) => negative_inputs_9_61_port, 
                           A_neg_shifted(60) => negative_inputs_9_60_port, 
                           A_neg_shifted(59) => negative_inputs_9_59_port, 
                           A_neg_shifted(58) => negative_inputs_9_58_port, 
                           A_neg_shifted(57) => negative_inputs_9_57_port, 
                           A_neg_shifted(56) => negative_inputs_9_56_port, 
                           A_neg_shifted(55) => negative_inputs_9_55_port, 
                           A_neg_shifted(54) => negative_inputs_9_54_port, 
                           A_neg_shifted(53) => negative_inputs_9_53_port, 
                           A_neg_shifted(52) => negative_inputs_9_52_port, 
                           A_neg_shifted(51) => negative_inputs_9_51_port, 
                           A_neg_shifted(50) => negative_inputs_9_50_port, 
                           A_neg_shifted(49) => negative_inputs_9_49_port, 
                           A_neg_shifted(48) => negative_inputs_9_48_port, 
                           A_neg_shifted(47) => n117, A_neg_shifted(46) => 
                           negative_inputs_9_46_port, A_neg_shifted(45) => 
                           negative_inputs_9_45_port, A_neg_shifted(44) => 
                           negative_inputs_9_44_port, A_neg_shifted(43) => 
                           negative_inputs_9_43_port, A_neg_shifted(42) => 
                           negative_inputs_9_42_port, A_neg_shifted(41) => 
                           negative_inputs_9_41_port, A_neg_shifted(40) => 
                           negative_inputs_9_40_port, A_neg_shifted(39) => 
                           negative_inputs_9_39_port, A_neg_shifted(38) => 
                           negative_inputs_9_38_port, A_neg_shifted(37) => 
                           negative_inputs_9_37_port, A_neg_shifted(36) => 
                           negative_inputs_9_36_port, A_neg_shifted(35) => 
                           negative_inputs_9_35_port, A_neg_shifted(34) => 
                           negative_inputs_9_34_port, A_neg_shifted(33) => 
                           negative_inputs_9_33_port, A_neg_shifted(32) => 
                           negative_inputs_9_32_port, A_neg_shifted(31) => 
                           negative_inputs_9_31_port, A_neg_shifted(30) => 
                           negative_inputs_9_30_port, A_neg_shifted(29) => 
                           negative_inputs_9_29_port, A_neg_shifted(28) => 
                           negative_inputs_9_28_port, A_neg_shifted(27) => 
                           negative_inputs_9_27_port, A_neg_shifted(26) => 
                           negative_inputs_9_26_port, A_neg_shifted(25) => 
                           negative_inputs_9_25_port, A_neg_shifted(24) => 
                           negative_inputs_9_24_port, A_neg_shifted(23) => 
                           negative_inputs_9_23_port, A_neg_shifted(22) => 
                           negative_inputs_9_22_port, A_neg_shifted(21) => 
                           negative_inputs_9_21_port, A_neg_shifted(20) => 
                           negative_inputs_9_20_port, A_neg_shifted(19) => 
                           negative_inputs_9_19_port, A_neg_shifted(18) => 
                           negative_inputs_9_18_port, A_neg_shifted(17) => 
                           negative_inputs_9_17_port, A_neg_shifted(16) => 
                           negative_inputs_9_16_port, A_neg_shifted(15) => 
                           negative_inputs_9_15_port, A_neg_shifted(14) => 
                           negative_inputs_9_14_port, A_neg_shifted(13) => 
                           negative_inputs_9_13_port, A_neg_shifted(12) => 
                           negative_inputs_9_12_port, A_neg_shifted(11) => 
                           negative_inputs_9_11_port, A_neg_shifted(10) => 
                           negative_inputs_9_10_port, A_neg_shifted(9) => 
                           negative_inputs_9_9_port, A_neg_shifted(8) => 
                           negative_inputs_9_8_port, A_neg_shifted(7) => 
                           negative_inputs_9_7_port, A_neg_shifted(6) => 
                           negative_inputs_9_6_port, A_neg_shifted(5) => 
                           negative_inputs_9_5_port, A_neg_shifted(4) => 
                           negative_inputs_9_4_port, A_neg_shifted(3) => 
                           negative_inputs_9_3_port, A_neg_shifted(2) => 
                           negative_inputs_9_2_port, A_neg_shifted(1) => 
                           negative_inputs_9_1_port, A_neg_shifted(0) => n8, 
                           Sel(2) => sel_4_2_port, Sel(1) => sel_4_1_port, 
                           Sel(0) => sel_4_0_port, Y(63) => 
                           MuxOutputs_4_63_port, Y(62) => MuxOutputs_4_62_port,
                           Y(61) => MuxOutputs_4_61_port, Y(60) => 
                           MuxOutputs_4_60_port, Y(59) => MuxOutputs_4_59_port,
                           Y(58) => MuxOutputs_4_58_port, Y(57) => 
                           MuxOutputs_4_57_port, Y(56) => MuxOutputs_4_56_port,
                           Y(55) => MuxOutputs_4_55_port, Y(54) => 
                           MuxOutputs_4_54_port, Y(53) => MuxOutputs_4_53_port,
                           Y(52) => MuxOutputs_4_52_port, Y(51) => 
                           MuxOutputs_4_51_port, Y(50) => MuxOutputs_4_50_port,
                           Y(49) => MuxOutputs_4_49_port, Y(48) => 
                           MuxOutputs_4_48_port, Y(47) => MuxOutputs_4_47_port,
                           Y(46) => MuxOutputs_4_46_port, Y(45) => 
                           MuxOutputs_4_45_port, Y(44) => MuxOutputs_4_44_port,
                           Y(43) => MuxOutputs_4_43_port, Y(42) => 
                           MuxOutputs_4_42_port, Y(41) => MuxOutputs_4_41_port,
                           Y(40) => MuxOutputs_4_40_port, Y(39) => 
                           MuxOutputs_4_39_port, Y(38) => MuxOutputs_4_38_port,
                           Y(37) => MuxOutputs_4_37_port, Y(36) => 
                           MuxOutputs_4_36_port, Y(35) => MuxOutputs_4_35_port,
                           Y(34) => MuxOutputs_4_34_port, Y(33) => 
                           MuxOutputs_4_33_port, Y(32) => MuxOutputs_4_32_port,
                           Y(31) => MuxOutputs_4_31_port, Y(30) => 
                           MuxOutputs_4_30_port, Y(29) => MuxOutputs_4_29_port,
                           Y(28) => MuxOutputs_4_28_port, Y(27) => 
                           MuxOutputs_4_27_port, Y(26) => MuxOutputs_4_26_port,
                           Y(25) => MuxOutputs_4_25_port, Y(24) => 
                           MuxOutputs_4_24_port, Y(23) => MuxOutputs_4_23_port,
                           Y(22) => MuxOutputs_4_22_port, Y(21) => 
                           MuxOutputs_4_21_port, Y(20) => MuxOutputs_4_20_port,
                           Y(19) => MuxOutputs_4_19_port, Y(18) => 
                           MuxOutputs_4_18_port, Y(17) => MuxOutputs_4_17_port,
                           Y(16) => MuxOutputs_4_16_port, Y(15) => 
                           MuxOutputs_4_15_port, Y(14) => MuxOutputs_4_14_port,
                           Y(13) => MuxOutputs_4_13_port, Y(12) => 
                           MuxOutputs_4_12_port, Y(11) => MuxOutputs_4_11_port,
                           Y(10) => MuxOutputs_4_10_port, Y(9) => 
                           MuxOutputs_4_9_port, Y(8) => MuxOutputs_4_8_port, 
                           Y(7) => MuxOutputs_4_7_port, Y(6) => 
                           MuxOutputs_4_6_port, Y(5) => MuxOutputs_4_5_port, 
                           Y(4) => MuxOutputs_4_4_port, Y(3) => 
                           MuxOutputs_4_3_port, Y(2) => MuxOutputs_4_2_port, 
                           Y(1) => MuxOutputs_4_1_port, Y(0) => 
                           MuxOutputs_4_0_port);
   encoderI_5 : encoder_27 port map( pieceofB(2) => B(11), pieceofB(1) => B(10)
                           , pieceofB(0) => B(9), sel(2) => sel_5_2_port, 
                           sel(1) => sel_5_1_port, sel(0) => sel_5_0_port);
   MUXI_5 : MUX51_MuxNbit64_27 port map( zeroSignal(63) => X_Logic0_port, 
                           zeroSignal(62) => X_Logic0_port, zeroSignal(61) => 
                           X_Logic0_port, zeroSignal(60) => X_Logic0_port, 
                           zeroSignal(59) => X_Logic0_port, zeroSignal(58) => 
                           X_Logic0_port, zeroSignal(57) => X_Logic0_port, 
                           zeroSignal(56) => X_Logic0_port, zeroSignal(55) => 
                           X_Logic0_port, zeroSignal(54) => X_Logic0_port, 
                           zeroSignal(53) => X_Logic0_port, zeroSignal(52) => 
                           X_Logic0_port, zeroSignal(51) => X_Logic0_port, 
                           zeroSignal(50) => X_Logic0_port, zeroSignal(49) => 
                           X_Logic0_port, zeroSignal(48) => X_Logic0_port, 
                           zeroSignal(47) => X_Logic0_port, zeroSignal(46) => 
                           X_Logic0_port, zeroSignal(45) => X_Logic0_port, 
                           zeroSignal(44) => X_Logic0_port, zeroSignal(43) => 
                           X_Logic0_port, zeroSignal(42) => X_Logic0_port, 
                           zeroSignal(41) => X_Logic0_port, zeroSignal(40) => 
                           X_Logic0_port, zeroSignal(39) => X_Logic0_port, 
                           zeroSignal(38) => X_Logic0_port, zeroSignal(37) => 
                           X_Logic0_port, zeroSignal(36) => X_Logic0_port, 
                           zeroSignal(35) => X_Logic0_port, zeroSignal(34) => 
                           X_Logic0_port, zeroSignal(33) => X_Logic0_port, 
                           zeroSignal(32) => X_Logic0_port, zeroSignal(31) => 
                           X_Logic0_port, zeroSignal(30) => X_Logic0_port, 
                           zeroSignal(29) => X_Logic0_port, zeroSignal(28) => 
                           X_Logic0_port, zeroSignal(27) => X_Logic0_port, 
                           zeroSignal(26) => X_Logic0_port, zeroSignal(25) => 
                           X_Logic0_port, zeroSignal(24) => X_Logic0_port, 
                           zeroSignal(23) => X_Logic0_port, zeroSignal(22) => 
                           X_Logic0_port, zeroSignal(21) => X_Logic0_port, 
                           zeroSignal(20) => X_Logic0_port, zeroSignal(19) => 
                           X_Logic0_port, zeroSignal(18) => X_Logic0_port, 
                           zeroSignal(17) => X_Logic0_port, zeroSignal(16) => 
                           X_Logic0_port, zeroSignal(15) => X_Logic0_port, 
                           zeroSignal(14) => X_Logic0_port, zeroSignal(13) => 
                           X_Logic0_port, zeroSignal(12) => X_Logic0_port, 
                           zeroSignal(11) => X_Logic0_port, zeroSignal(10) => 
                           X_Logic0_port, zeroSignal(9) => X_Logic0_port, 
                           zeroSignal(8) => X_Logic0_port, zeroSignal(7) => 
                           X_Logic0_port, zeroSignal(6) => X_Logic0_port, 
                           zeroSignal(5) => X_Logic0_port, zeroSignal(4) => 
                           X_Logic0_port, zeroSignal(3) => X_Logic0_port, 
                           zeroSignal(2) => X_Logic0_port, zeroSignal(1) => 
                           X_Logic0_port, zeroSignal(0) => X_Logic0_port, 
                           A_signal(63) => positive_inputs_10_63_port, 
                           A_signal(62) => positive_inputs_10_62_port, 
                           A_signal(61) => positive_inputs_10_61_port, 
                           A_signal(60) => positive_inputs_10_60_port, 
                           A_signal(59) => positive_inputs_10_59_port, 
                           A_signal(58) => positive_inputs_10_58_port, 
                           A_signal(57) => positive_inputs_10_57_port, 
                           A_signal(56) => positive_inputs_10_56_port, 
                           A_signal(55) => positive_inputs_10_55_port, 
                           A_signal(54) => positive_inputs_10_54_port, 
                           A_signal(53) => positive_inputs_10_53_port, 
                           A_signal(52) => positive_inputs_10_52_port, 
                           A_signal(51) => positive_inputs_10_51_port, 
                           A_signal(50) => positive_inputs_10_50_port, 
                           A_signal(49) => positive_inputs_10_49_port, 
                           A_signal(48) => positive_inputs_10_48_port, 
                           A_signal(47) => n31, A_signal(46) => 
                           positive_inputs_10_46_port, A_signal(45) => 
                           positive_inputs_10_45_port, A_signal(44) => 
                           positive_inputs_10_44_port, A_signal(43) => 
                           positive_inputs_10_43_port, A_signal(42) => 
                           positive_inputs_10_42_port, A_signal(41) => 
                           positive_inputs_10_41_port, A_signal(40) => 
                           positive_inputs_10_40_port, A_signal(39) => 
                           positive_inputs_10_39_port, A_signal(38) => 
                           positive_inputs_10_38_port, A_signal(37) => 
                           positive_inputs_10_37_port, A_signal(36) => 
                           positive_inputs_10_36_port, A_signal(35) => 
                           positive_inputs_10_35_port, A_signal(34) => 
                           positive_inputs_10_34_port, A_signal(33) => 
                           positive_inputs_10_33_port, A_signal(32) => 
                           positive_inputs_10_32_port, A_signal(31) => 
                           positive_inputs_10_31_port, A_signal(30) => 
                           positive_inputs_10_30_port, A_signal(29) => 
                           positive_inputs_10_29_port, A_signal(28) => 
                           positive_inputs_10_28_port, A_signal(27) => 
                           positive_inputs_10_27_port, A_signal(26) => 
                           positive_inputs_10_26_port, A_signal(25) => 
                           positive_inputs_10_25_port, A_signal(24) => 
                           positive_inputs_10_24_port, A_signal(23) => 
                           positive_inputs_10_23_port, A_signal(22) => 
                           positive_inputs_10_22_port, A_signal(21) => 
                           positive_inputs_10_21_port, A_signal(20) => 
                           positive_inputs_10_20_port, A_signal(19) => 
                           positive_inputs_10_19_port, A_signal(18) => 
                           positive_inputs_10_18_port, A_signal(17) => 
                           positive_inputs_10_17_port, A_signal(16) => 
                           positive_inputs_10_16_port, A_signal(15) => 
                           positive_inputs_10_15_port, A_signal(14) => 
                           positive_inputs_10_14_port, A_signal(13) => 
                           positive_inputs_10_13_port, A_signal(12) => 
                           positive_inputs_10_12_port, A_signal(11) => 
                           positive_inputs_10_11_port, A_signal(10) => 
                           positive_inputs_10_10_port, A_signal(9) => 
                           positive_inputs_10_9_port, A_signal(8) => 
                           positive_inputs_10_8_port, A_signal(7) => 
                           positive_inputs_10_7_port, A_signal(6) => 
                           positive_inputs_10_6_port, A_signal(5) => 
                           positive_inputs_10_5_port, A_signal(4) => 
                           positive_inputs_10_4_port, A_signal(3) => 
                           positive_inputs_10_3_port, A_signal(2) => 
                           positive_inputs_10_2_port, A_signal(1) => 
                           positive_inputs_10_1_port, A_signal(0) => n8, 
                           A_neg(63) => negative_inputs_10_63_port, A_neg(62) 
                           => negative_inputs_10_62_port, A_neg(61) => 
                           negative_inputs_10_61_port, A_neg(60) => 
                           negative_inputs_10_60_port, A_neg(59) => 
                           negative_inputs_10_59_port, A_neg(58) => 
                           negative_inputs_10_58_port, A_neg(57) => 
                           negative_inputs_10_57_port, A_neg(56) => 
                           negative_inputs_10_56_port, A_neg(55) => 
                           negative_inputs_10_55_port, A_neg(54) => 
                           negative_inputs_10_54_port, A_neg(53) => 
                           negative_inputs_10_53_port, A_neg(52) => 
                           negative_inputs_10_52_port, A_neg(51) => 
                           negative_inputs_10_51_port, A_neg(50) => 
                           negative_inputs_10_50_port, A_neg(49) => 
                           negative_inputs_10_49_port, A_neg(48) => 
                           negative_inputs_10_48_port, A_neg(47) => n116, 
                           A_neg(46) => negative_inputs_10_46_port, A_neg(45) 
                           => negative_inputs_10_45_port, A_neg(44) => 
                           negative_inputs_10_44_port, A_neg(43) => 
                           negative_inputs_10_43_port, A_neg(42) => 
                           negative_inputs_10_42_port, A_neg(41) => 
                           negative_inputs_10_41_port, A_neg(40) => 
                           negative_inputs_10_40_port, A_neg(39) => 
                           negative_inputs_10_39_port, A_neg(38) => 
                           negative_inputs_10_38_port, A_neg(37) => 
                           negative_inputs_10_37_port, A_neg(36) => 
                           negative_inputs_10_36_port, A_neg(35) => 
                           negative_inputs_10_35_port, A_neg(34) => 
                           negative_inputs_10_34_port, A_neg(33) => 
                           negative_inputs_10_33_port, A_neg(32) => 
                           negative_inputs_10_32_port, A_neg(31) => 
                           negative_inputs_10_31_port, A_neg(30) => 
                           negative_inputs_10_30_port, A_neg(29) => 
                           negative_inputs_10_29_port, A_neg(28) => 
                           negative_inputs_10_28_port, A_neg(27) => 
                           negative_inputs_10_27_port, A_neg(26) => 
                           negative_inputs_10_26_port, A_neg(25) => 
                           negative_inputs_10_25_port, A_neg(24) => 
                           negative_inputs_10_24_port, A_neg(23) => 
                           negative_inputs_10_23_port, A_neg(22) => 
                           negative_inputs_10_22_port, A_neg(21) => 
                           negative_inputs_10_21_port, A_neg(20) => 
                           negative_inputs_10_20_port, A_neg(19) => 
                           negative_inputs_10_19_port, A_neg(18) => 
                           negative_inputs_10_18_port, A_neg(17) => 
                           negative_inputs_10_17_port, A_neg(16) => 
                           negative_inputs_10_16_port, A_neg(15) => 
                           negative_inputs_10_15_port, A_neg(14) => 
                           negative_inputs_10_14_port, A_neg(13) => 
                           negative_inputs_10_13_port, A_neg(12) => 
                           negative_inputs_10_12_port, A_neg(11) => 
                           negative_inputs_10_11_port, A_neg(10) => 
                           negative_inputs_10_10_port, A_neg(9) => 
                           negative_inputs_10_9_port, A_neg(8) => 
                           negative_inputs_10_8_port, A_neg(7) => 
                           negative_inputs_10_7_port, A_neg(6) => 
                           negative_inputs_10_6_port, A_neg(5) => 
                           negative_inputs_10_5_port, A_neg(4) => 
                           negative_inputs_10_4_port, A_neg(3) => 
                           negative_inputs_10_3_port, A_neg(2) => 
                           negative_inputs_10_2_port, A_neg(1) => 
                           negative_inputs_10_1_port, A_neg(0) => n8, 
                           A_shifted(63) => positive_inputs_11_63_port, 
                           A_shifted(62) => positive_inputs_11_62_port, 
                           A_shifted(61) => positive_inputs_11_61_port, 
                           A_shifted(60) => positive_inputs_11_60_port, 
                           A_shifted(59) => positive_inputs_11_59_port, 
                           A_shifted(58) => positive_inputs_11_58_port, 
                           A_shifted(57) => positive_inputs_11_57_port, 
                           A_shifted(56) => positive_inputs_11_56_port, 
                           A_shifted(55) => positive_inputs_11_55_port, 
                           A_shifted(54) => positive_inputs_11_54_port, 
                           A_shifted(53) => positive_inputs_11_53_port, 
                           A_shifted(52) => positive_inputs_11_52_port, 
                           A_shifted(51) => positive_inputs_11_51_port, 
                           A_shifted(50) => positive_inputs_11_50_port, 
                           A_shifted(49) => positive_inputs_11_49_port, 
                           A_shifted(48) => positive_inputs_11_48_port, 
                           A_shifted(47) => n30, A_shifted(46) => 
                           positive_inputs_11_46_port, A_shifted(45) => 
                           positive_inputs_11_45_port, A_shifted(44) => 
                           positive_inputs_11_44_port, A_shifted(43) => 
                           positive_inputs_11_43_port, A_shifted(42) => 
                           positive_inputs_11_42_port, A_shifted(41) => 
                           positive_inputs_11_41_port, A_shifted(40) => 
                           positive_inputs_11_40_port, A_shifted(39) => 
                           positive_inputs_11_39_port, A_shifted(38) => 
                           positive_inputs_11_38_port, A_shifted(37) => 
                           positive_inputs_11_37_port, A_shifted(36) => 
                           positive_inputs_11_36_port, A_shifted(35) => 
                           positive_inputs_11_35_port, A_shifted(34) => 
                           positive_inputs_11_34_port, A_shifted(33) => 
                           positive_inputs_11_33_port, A_shifted(32) => 
                           positive_inputs_11_32_port, A_shifted(31) => 
                           positive_inputs_11_31_port, A_shifted(30) => 
                           positive_inputs_11_30_port, A_shifted(29) => 
                           positive_inputs_11_29_port, A_shifted(28) => 
                           positive_inputs_11_28_port, A_shifted(27) => 
                           positive_inputs_11_27_port, A_shifted(26) => 
                           positive_inputs_11_26_port, A_shifted(25) => 
                           positive_inputs_11_25_port, A_shifted(24) => 
                           positive_inputs_11_24_port, A_shifted(23) => 
                           positive_inputs_11_23_port, A_shifted(22) => 
                           positive_inputs_11_22_port, A_shifted(21) => 
                           positive_inputs_11_21_port, A_shifted(20) => 
                           positive_inputs_11_20_port, A_shifted(19) => 
                           positive_inputs_11_19_port, A_shifted(18) => 
                           positive_inputs_11_18_port, A_shifted(17) => 
                           positive_inputs_11_17_port, A_shifted(16) => 
                           positive_inputs_11_16_port, A_shifted(15) => 
                           positive_inputs_11_15_port, A_shifted(14) => 
                           positive_inputs_11_14_port, A_shifted(13) => 
                           positive_inputs_11_13_port, A_shifted(12) => 
                           positive_inputs_11_12_port, A_shifted(11) => 
                           positive_inputs_11_11_port, A_shifted(10) => 
                           positive_inputs_11_10_port, A_shifted(9) => 
                           positive_inputs_11_9_port, A_shifted(8) => 
                           positive_inputs_11_8_port, A_shifted(7) => 
                           positive_inputs_11_7_port, A_shifted(6) => 
                           positive_inputs_11_6_port, A_shifted(5) => 
                           positive_inputs_11_5_port, A_shifted(4) => 
                           positive_inputs_11_4_port, A_shifted(3) => 
                           positive_inputs_11_3_port, A_shifted(2) => 
                           positive_inputs_11_2_port, A_shifted(1) => 
                           positive_inputs_11_1_port, A_shifted(0) => n8, 
                           A_neg_shifted(63) => negative_inputs_11_63_port, 
                           A_neg_shifted(62) => negative_inputs_11_62_port, 
                           A_neg_shifted(61) => negative_inputs_11_61_port, 
                           A_neg_shifted(60) => negative_inputs_11_60_port, 
                           A_neg_shifted(59) => negative_inputs_11_59_port, 
                           A_neg_shifted(58) => negative_inputs_11_58_port, 
                           A_neg_shifted(57) => negative_inputs_11_57_port, 
                           A_neg_shifted(56) => negative_inputs_11_56_port, 
                           A_neg_shifted(55) => negative_inputs_11_55_port, 
                           A_neg_shifted(54) => negative_inputs_11_54_port, 
                           A_neg_shifted(53) => negative_inputs_11_53_port, 
                           A_neg_shifted(52) => negative_inputs_11_52_port, 
                           A_neg_shifted(51) => negative_inputs_11_51_port, 
                           A_neg_shifted(50) => negative_inputs_11_50_port, 
                           A_neg_shifted(49) => negative_inputs_11_49_port, 
                           A_neg_shifted(48) => negative_inputs_11_48_port, 
                           A_neg_shifted(47) => n115, A_neg_shifted(46) => 
                           negative_inputs_11_46_port, A_neg_shifted(45) => 
                           negative_inputs_11_45_port, A_neg_shifted(44) => 
                           negative_inputs_11_44_port, A_neg_shifted(43) => 
                           negative_inputs_11_43_port, A_neg_shifted(42) => 
                           negative_inputs_11_42_port, A_neg_shifted(41) => 
                           negative_inputs_11_41_port, A_neg_shifted(40) => 
                           negative_inputs_11_40_port, A_neg_shifted(39) => 
                           negative_inputs_11_39_port, A_neg_shifted(38) => 
                           negative_inputs_11_38_port, A_neg_shifted(37) => 
                           negative_inputs_11_37_port, A_neg_shifted(36) => 
                           negative_inputs_11_36_port, A_neg_shifted(35) => 
                           negative_inputs_11_35_port, A_neg_shifted(34) => 
                           negative_inputs_11_34_port, A_neg_shifted(33) => 
                           negative_inputs_11_33_port, A_neg_shifted(32) => 
                           negative_inputs_11_32_port, A_neg_shifted(31) => 
                           negative_inputs_11_31_port, A_neg_shifted(30) => 
                           negative_inputs_11_30_port, A_neg_shifted(29) => 
                           negative_inputs_11_29_port, A_neg_shifted(28) => 
                           negative_inputs_11_28_port, A_neg_shifted(27) => 
                           negative_inputs_11_27_port, A_neg_shifted(26) => 
                           negative_inputs_11_26_port, A_neg_shifted(25) => 
                           negative_inputs_11_25_port, A_neg_shifted(24) => 
                           negative_inputs_11_24_port, A_neg_shifted(23) => 
                           negative_inputs_11_23_port, A_neg_shifted(22) => 
                           negative_inputs_11_22_port, A_neg_shifted(21) => 
                           negative_inputs_11_21_port, A_neg_shifted(20) => 
                           negative_inputs_11_20_port, A_neg_shifted(19) => 
                           negative_inputs_11_19_port, A_neg_shifted(18) => 
                           negative_inputs_11_18_port, A_neg_shifted(17) => 
                           negative_inputs_11_17_port, A_neg_shifted(16) => 
                           negative_inputs_11_16_port, A_neg_shifted(15) => 
                           negative_inputs_11_15_port, A_neg_shifted(14) => 
                           negative_inputs_11_14_port, A_neg_shifted(13) => 
                           negative_inputs_11_13_port, A_neg_shifted(12) => 
                           negative_inputs_11_12_port, A_neg_shifted(11) => 
                           negative_inputs_11_11_port, A_neg_shifted(10) => 
                           negative_inputs_11_10_port, A_neg_shifted(9) => 
                           negative_inputs_11_9_port, A_neg_shifted(8) => 
                           negative_inputs_11_8_port, A_neg_shifted(7) => 
                           negative_inputs_11_7_port, A_neg_shifted(6) => 
                           negative_inputs_11_6_port, A_neg_shifted(5) => 
                           negative_inputs_11_5_port, A_neg_shifted(4) => 
                           negative_inputs_11_4_port, A_neg_shifted(3) => 
                           negative_inputs_11_3_port, A_neg_shifted(2) => 
                           negative_inputs_11_2_port, A_neg_shifted(1) => 
                           negative_inputs_11_1_port, A_neg_shifted(0) => n8, 
                           Sel(2) => sel_5_2_port, Sel(1) => sel_5_1_port, 
                           Sel(0) => sel_5_0_port, Y(63) => 
                           MuxOutputs_5_63_port, Y(62) => MuxOutputs_5_62_port,
                           Y(61) => MuxOutputs_5_61_port, Y(60) => 
                           MuxOutputs_5_60_port, Y(59) => MuxOutputs_5_59_port,
                           Y(58) => MuxOutputs_5_58_port, Y(57) => 
                           MuxOutputs_5_57_port, Y(56) => MuxOutputs_5_56_port,
                           Y(55) => MuxOutputs_5_55_port, Y(54) => 
                           MuxOutputs_5_54_port, Y(53) => MuxOutputs_5_53_port,
                           Y(52) => MuxOutputs_5_52_port, Y(51) => 
                           MuxOutputs_5_51_port, Y(50) => MuxOutputs_5_50_port,
                           Y(49) => MuxOutputs_5_49_port, Y(48) => 
                           MuxOutputs_5_48_port, Y(47) => MuxOutputs_5_47_port,
                           Y(46) => MuxOutputs_5_46_port, Y(45) => 
                           MuxOutputs_5_45_port, Y(44) => MuxOutputs_5_44_port,
                           Y(43) => MuxOutputs_5_43_port, Y(42) => 
                           MuxOutputs_5_42_port, Y(41) => MuxOutputs_5_41_port,
                           Y(40) => MuxOutputs_5_40_port, Y(39) => 
                           MuxOutputs_5_39_port, Y(38) => MuxOutputs_5_38_port,
                           Y(37) => MuxOutputs_5_37_port, Y(36) => 
                           MuxOutputs_5_36_port, Y(35) => MuxOutputs_5_35_port,
                           Y(34) => MuxOutputs_5_34_port, Y(33) => 
                           MuxOutputs_5_33_port, Y(32) => MuxOutputs_5_32_port,
                           Y(31) => MuxOutputs_5_31_port, Y(30) => 
                           MuxOutputs_5_30_port, Y(29) => MuxOutputs_5_29_port,
                           Y(28) => MuxOutputs_5_28_port, Y(27) => 
                           MuxOutputs_5_27_port, Y(26) => MuxOutputs_5_26_port,
                           Y(25) => MuxOutputs_5_25_port, Y(24) => 
                           MuxOutputs_5_24_port, Y(23) => MuxOutputs_5_23_port,
                           Y(22) => MuxOutputs_5_22_port, Y(21) => 
                           MuxOutputs_5_21_port, Y(20) => MuxOutputs_5_20_port,
                           Y(19) => MuxOutputs_5_19_port, Y(18) => 
                           MuxOutputs_5_18_port, Y(17) => MuxOutputs_5_17_port,
                           Y(16) => MuxOutputs_5_16_port, Y(15) => 
                           MuxOutputs_5_15_port, Y(14) => MuxOutputs_5_14_port,
                           Y(13) => MuxOutputs_5_13_port, Y(12) => 
                           MuxOutputs_5_12_port, Y(11) => MuxOutputs_5_11_port,
                           Y(10) => MuxOutputs_5_10_port, Y(9) => 
                           MuxOutputs_5_9_port, Y(8) => MuxOutputs_5_8_port, 
                           Y(7) => MuxOutputs_5_7_port, Y(6) => 
                           MuxOutputs_5_6_port, Y(5) => MuxOutputs_5_5_port, 
                           Y(4) => MuxOutputs_5_4_port, Y(3) => 
                           MuxOutputs_5_3_port, Y(2) => MuxOutputs_5_2_port, 
                           Y(1) => MuxOutputs_5_1_port, Y(0) => 
                           MuxOutputs_5_0_port);
   encoderI_6 : encoder_26 port map( pieceofB(2) => B(13), pieceofB(1) => B(12)
                           , pieceofB(0) => B(11), sel(2) => sel_6_2_port, 
                           sel(1) => sel_6_1_port, sel(0) => sel_6_0_port);
   MUXI_6 : MUX51_MuxNbit64_26 port map( zeroSignal(63) => X_Logic0_port, 
                           zeroSignal(62) => X_Logic0_port, zeroSignal(61) => 
                           X_Logic0_port, zeroSignal(60) => X_Logic0_port, 
                           zeroSignal(59) => X_Logic0_port, zeroSignal(58) => 
                           X_Logic0_port, zeroSignal(57) => X_Logic0_port, 
                           zeroSignal(56) => X_Logic0_port, zeroSignal(55) => 
                           X_Logic0_port, zeroSignal(54) => X_Logic0_port, 
                           zeroSignal(53) => X_Logic0_port, zeroSignal(52) => 
                           X_Logic0_port, zeroSignal(51) => X_Logic0_port, 
                           zeroSignal(50) => X_Logic0_port, zeroSignal(49) => 
                           X_Logic0_port, zeroSignal(48) => X_Logic0_port, 
                           zeroSignal(47) => X_Logic0_port, zeroSignal(46) => 
                           X_Logic0_port, zeroSignal(45) => X_Logic0_port, 
                           zeroSignal(44) => X_Logic0_port, zeroSignal(43) => 
                           X_Logic0_port, zeroSignal(42) => X_Logic0_port, 
                           zeroSignal(41) => X_Logic0_port, zeroSignal(40) => 
                           X_Logic0_port, zeroSignal(39) => X_Logic0_port, 
                           zeroSignal(38) => X_Logic0_port, zeroSignal(37) => 
                           X_Logic0_port, zeroSignal(36) => X_Logic0_port, 
                           zeroSignal(35) => X_Logic0_port, zeroSignal(34) => 
                           X_Logic0_port, zeroSignal(33) => X_Logic0_port, 
                           zeroSignal(32) => X_Logic0_port, zeroSignal(31) => 
                           X_Logic0_port, zeroSignal(30) => X_Logic0_port, 
                           zeroSignal(29) => X_Logic0_port, zeroSignal(28) => 
                           X_Logic0_port, zeroSignal(27) => X_Logic0_port, 
                           zeroSignal(26) => X_Logic0_port, zeroSignal(25) => 
                           X_Logic0_port, zeroSignal(24) => X_Logic0_port, 
                           zeroSignal(23) => X_Logic0_port, zeroSignal(22) => 
                           X_Logic0_port, zeroSignal(21) => X_Logic0_port, 
                           zeroSignal(20) => X_Logic0_port, zeroSignal(19) => 
                           X_Logic0_port, zeroSignal(18) => X_Logic0_port, 
                           zeroSignal(17) => X_Logic0_port, zeroSignal(16) => 
                           X_Logic0_port, zeroSignal(15) => X_Logic0_port, 
                           zeroSignal(14) => X_Logic0_port, zeroSignal(13) => 
                           X_Logic0_port, zeroSignal(12) => X_Logic0_port, 
                           zeroSignal(11) => X_Logic0_port, zeroSignal(10) => 
                           X_Logic0_port, zeroSignal(9) => X_Logic0_port, 
                           zeroSignal(8) => X_Logic0_port, zeroSignal(7) => 
                           X_Logic0_port, zeroSignal(6) => X_Logic0_port, 
                           zeroSignal(5) => X_Logic0_port, zeroSignal(4) => 
                           X_Logic0_port, zeroSignal(3) => X_Logic0_port, 
                           zeroSignal(2) => X_Logic0_port, zeroSignal(1) => 
                           X_Logic0_port, zeroSignal(0) => X_Logic0_port, 
                           A_signal(63) => positive_inputs_12_63_port, 
                           A_signal(62) => positive_inputs_12_62_port, 
                           A_signal(61) => positive_inputs_12_61_port, 
                           A_signal(60) => positive_inputs_12_60_port, 
                           A_signal(59) => positive_inputs_12_59_port, 
                           A_signal(58) => positive_inputs_12_58_port, 
                           A_signal(57) => positive_inputs_12_57_port, 
                           A_signal(56) => positive_inputs_12_56_port, 
                           A_signal(55) => positive_inputs_12_55_port, 
                           A_signal(54) => positive_inputs_12_54_port, 
                           A_signal(53) => positive_inputs_12_53_port, 
                           A_signal(52) => positive_inputs_12_52_port, 
                           A_signal(51) => positive_inputs_12_51_port, 
                           A_signal(50) => positive_inputs_12_50_port, 
                           A_signal(49) => positive_inputs_12_49_port, 
                           A_signal(48) => positive_inputs_12_48_port, 
                           A_signal(47) => n29, A_signal(46) => 
                           positive_inputs_12_46_port, A_signal(45) => 
                           positive_inputs_12_45_port, A_signal(44) => 
                           positive_inputs_12_44_port, A_signal(43) => 
                           positive_inputs_12_43_port, A_signal(42) => 
                           positive_inputs_12_42_port, A_signal(41) => 
                           positive_inputs_12_41_port, A_signal(40) => 
                           positive_inputs_12_40_port, A_signal(39) => 
                           positive_inputs_12_39_port, A_signal(38) => 
                           positive_inputs_12_38_port, A_signal(37) => 
                           positive_inputs_12_37_port, A_signal(36) => 
                           positive_inputs_12_36_port, A_signal(35) => 
                           positive_inputs_12_35_port, A_signal(34) => 
                           positive_inputs_12_34_port, A_signal(33) => 
                           positive_inputs_12_33_port, A_signal(32) => 
                           positive_inputs_12_32_port, A_signal(31) => 
                           positive_inputs_12_31_port, A_signal(30) => 
                           positive_inputs_12_30_port, A_signal(29) => 
                           positive_inputs_12_29_port, A_signal(28) => 
                           positive_inputs_12_28_port, A_signal(27) => 
                           positive_inputs_12_27_port, A_signal(26) => 
                           positive_inputs_12_26_port, A_signal(25) => 
                           positive_inputs_12_25_port, A_signal(24) => 
                           positive_inputs_12_24_port, A_signal(23) => 
                           positive_inputs_12_23_port, A_signal(22) => 
                           positive_inputs_12_22_port, A_signal(21) => 
                           positive_inputs_12_21_port, A_signal(20) => 
                           positive_inputs_12_20_port, A_signal(19) => 
                           positive_inputs_12_19_port, A_signal(18) => 
                           positive_inputs_12_18_port, A_signal(17) => 
                           positive_inputs_12_17_port, A_signal(16) => 
                           positive_inputs_12_16_port, A_signal(15) => 
                           positive_inputs_12_15_port, A_signal(14) => 
                           positive_inputs_12_14_port, A_signal(13) => 
                           positive_inputs_12_13_port, A_signal(12) => 
                           positive_inputs_12_12_port, A_signal(11) => 
                           positive_inputs_12_11_port, A_signal(10) => 
                           positive_inputs_12_10_port, A_signal(9) => 
                           positive_inputs_12_9_port, A_signal(8) => 
                           positive_inputs_12_8_port, A_signal(7) => 
                           positive_inputs_12_7_port, A_signal(6) => 
                           positive_inputs_12_6_port, A_signal(5) => 
                           positive_inputs_12_5_port, A_signal(4) => 
                           positive_inputs_12_4_port, A_signal(3) => 
                           positive_inputs_12_3_port, A_signal(2) => 
                           positive_inputs_12_2_port, A_signal(1) => 
                           positive_inputs_12_1_port, A_signal(0) => n8, 
                           A_neg(63) => negative_inputs_12_63_port, A_neg(62) 
                           => negative_inputs_12_62_port, A_neg(61) => 
                           negative_inputs_12_61_port, A_neg(60) => 
                           negative_inputs_12_60_port, A_neg(59) => 
                           negative_inputs_12_59_port, A_neg(58) => 
                           negative_inputs_12_58_port, A_neg(57) => 
                           negative_inputs_12_57_port, A_neg(56) => 
                           negative_inputs_12_56_port, A_neg(55) => 
                           negative_inputs_12_55_port, A_neg(54) => 
                           negative_inputs_12_54_port, A_neg(53) => 
                           negative_inputs_12_53_port, A_neg(52) => 
                           negative_inputs_12_52_port, A_neg(51) => 
                           negative_inputs_12_51_port, A_neg(50) => 
                           negative_inputs_12_50_port, A_neg(49) => 
                           negative_inputs_12_49_port, A_neg(48) => 
                           negative_inputs_12_48_port, A_neg(47) => n113, 
                           A_neg(46) => negative_inputs_12_46_port, A_neg(45) 
                           => negative_inputs_12_45_port, A_neg(44) => 
                           negative_inputs_12_44_port, A_neg(43) => 
                           negative_inputs_12_43_port, A_neg(42) => 
                           negative_inputs_12_42_port, A_neg(41) => 
                           negative_inputs_12_41_port, A_neg(40) => 
                           negative_inputs_12_40_port, A_neg(39) => 
                           negative_inputs_12_39_port, A_neg(38) => 
                           negative_inputs_12_38_port, A_neg(37) => 
                           negative_inputs_12_37_port, A_neg(36) => 
                           negative_inputs_12_36_port, A_neg(35) => 
                           negative_inputs_12_35_port, A_neg(34) => 
                           negative_inputs_12_34_port, A_neg(33) => 
                           negative_inputs_12_33_port, A_neg(32) => 
                           negative_inputs_12_32_port, A_neg(31) => 
                           negative_inputs_12_31_port, A_neg(30) => 
                           negative_inputs_12_30_port, A_neg(29) => 
                           negative_inputs_12_29_port, A_neg(28) => 
                           negative_inputs_12_28_port, A_neg(27) => 
                           negative_inputs_12_27_port, A_neg(26) => 
                           negative_inputs_12_26_port, A_neg(25) => 
                           negative_inputs_12_25_port, A_neg(24) => 
                           negative_inputs_12_24_port, A_neg(23) => 
                           negative_inputs_12_23_port, A_neg(22) => 
                           negative_inputs_12_22_port, A_neg(21) => 
                           negative_inputs_12_21_port, A_neg(20) => 
                           negative_inputs_12_20_port, A_neg(19) => 
                           negative_inputs_12_19_port, A_neg(18) => 
                           negative_inputs_12_18_port, A_neg(17) => 
                           negative_inputs_12_17_port, A_neg(16) => 
                           negative_inputs_12_16_port, A_neg(15) => 
                           negative_inputs_12_15_port, A_neg(14) => 
                           negative_inputs_12_14_port, A_neg(13) => 
                           negative_inputs_12_13_port, A_neg(12) => 
                           negative_inputs_12_12_port, A_neg(11) => 
                           negative_inputs_12_11_port, A_neg(10) => 
                           negative_inputs_12_10_port, A_neg(9) => 
                           negative_inputs_12_9_port, A_neg(8) => 
                           negative_inputs_12_8_port, A_neg(7) => 
                           negative_inputs_12_7_port, A_neg(6) => 
                           negative_inputs_12_6_port, A_neg(5) => 
                           negative_inputs_12_5_port, A_neg(4) => 
                           negative_inputs_12_4_port, A_neg(3) => 
                           negative_inputs_12_3_port, A_neg(2) => 
                           negative_inputs_12_2_port, A_neg(1) => 
                           negative_inputs_12_1_port, A_neg(0) => n8, 
                           A_shifted(63) => positive_inputs_13_63_port, 
                           A_shifted(62) => positive_inputs_13_62_port, 
                           A_shifted(61) => positive_inputs_13_61_port, 
                           A_shifted(60) => positive_inputs_13_60_port, 
                           A_shifted(59) => positive_inputs_13_59_port, 
                           A_shifted(58) => positive_inputs_13_58_port, 
                           A_shifted(57) => positive_inputs_13_57_port, 
                           A_shifted(56) => positive_inputs_13_56_port, 
                           A_shifted(55) => positive_inputs_13_55_port, 
                           A_shifted(54) => positive_inputs_13_54_port, 
                           A_shifted(53) => positive_inputs_13_53_port, 
                           A_shifted(52) => positive_inputs_13_52_port, 
                           A_shifted(51) => positive_inputs_13_51_port, 
                           A_shifted(50) => positive_inputs_13_50_port, 
                           A_shifted(49) => positive_inputs_13_49_port, 
                           A_shifted(48) => positive_inputs_13_48_port, 
                           A_shifted(47) => n28, A_shifted(46) => 
                           positive_inputs_13_46_port, A_shifted(45) => 
                           positive_inputs_13_45_port, A_shifted(44) => 
                           positive_inputs_13_44_port, A_shifted(43) => 
                           positive_inputs_13_43_port, A_shifted(42) => 
                           positive_inputs_13_42_port, A_shifted(41) => 
                           positive_inputs_13_41_port, A_shifted(40) => 
                           positive_inputs_13_40_port, A_shifted(39) => 
                           positive_inputs_13_39_port, A_shifted(38) => 
                           positive_inputs_13_38_port, A_shifted(37) => 
                           positive_inputs_13_37_port, A_shifted(36) => 
                           positive_inputs_13_36_port, A_shifted(35) => 
                           positive_inputs_13_35_port, A_shifted(34) => 
                           positive_inputs_13_34_port, A_shifted(33) => 
                           positive_inputs_13_33_port, A_shifted(32) => 
                           positive_inputs_13_32_port, A_shifted(31) => 
                           positive_inputs_13_31_port, A_shifted(30) => 
                           positive_inputs_13_30_port, A_shifted(29) => 
                           positive_inputs_13_29_port, A_shifted(28) => 
                           positive_inputs_13_28_port, A_shifted(27) => 
                           positive_inputs_13_27_port, A_shifted(26) => 
                           positive_inputs_13_26_port, A_shifted(25) => 
                           positive_inputs_13_25_port, A_shifted(24) => 
                           positive_inputs_13_24_port, A_shifted(23) => 
                           positive_inputs_13_23_port, A_shifted(22) => 
                           positive_inputs_13_22_port, A_shifted(21) => 
                           positive_inputs_13_21_port, A_shifted(20) => 
                           positive_inputs_13_20_port, A_shifted(19) => 
                           positive_inputs_13_19_port, A_shifted(18) => 
                           positive_inputs_13_18_port, A_shifted(17) => 
                           positive_inputs_13_17_port, A_shifted(16) => 
                           positive_inputs_13_16_port, A_shifted(15) => 
                           positive_inputs_13_15_port, A_shifted(14) => 
                           positive_inputs_13_14_port, A_shifted(13) => 
                           positive_inputs_13_13_port, A_shifted(12) => 
                           positive_inputs_13_12_port, A_shifted(11) => 
                           positive_inputs_13_11_port, A_shifted(10) => 
                           positive_inputs_13_10_port, A_shifted(9) => 
                           positive_inputs_13_9_port, A_shifted(8) => 
                           positive_inputs_13_8_port, A_shifted(7) => 
                           positive_inputs_13_7_port, A_shifted(6) => 
                           positive_inputs_13_6_port, A_shifted(5) => 
                           positive_inputs_13_5_port, A_shifted(4) => 
                           positive_inputs_13_4_port, A_shifted(3) => 
                           positive_inputs_13_3_port, A_shifted(2) => 
                           positive_inputs_13_2_port, A_shifted(1) => 
                           positive_inputs_13_1_port, A_shifted(0) => n8, 
                           A_neg_shifted(63) => negative_inputs_13_63_port, 
                           A_neg_shifted(62) => negative_inputs_13_62_port, 
                           A_neg_shifted(61) => negative_inputs_13_61_port, 
                           A_neg_shifted(60) => negative_inputs_13_60_port, 
                           A_neg_shifted(59) => negative_inputs_13_59_port, 
                           A_neg_shifted(58) => negative_inputs_13_58_port, 
                           A_neg_shifted(57) => negative_inputs_13_57_port, 
                           A_neg_shifted(56) => negative_inputs_13_56_port, 
                           A_neg_shifted(55) => negative_inputs_13_55_port, 
                           A_neg_shifted(54) => negative_inputs_13_54_port, 
                           A_neg_shifted(53) => negative_inputs_13_53_port, 
                           A_neg_shifted(52) => negative_inputs_13_52_port, 
                           A_neg_shifted(51) => negative_inputs_13_51_port, 
                           A_neg_shifted(50) => negative_inputs_13_50_port, 
                           A_neg_shifted(49) => negative_inputs_13_49_port, 
                           A_neg_shifted(48) => negative_inputs_13_48_port, 
                           A_neg_shifted(47) => n111, A_neg_shifted(46) => 
                           negative_inputs_13_46_port, A_neg_shifted(45) => 
                           negative_inputs_13_45_port, A_neg_shifted(44) => 
                           negative_inputs_13_44_port, A_neg_shifted(43) => 
                           negative_inputs_13_43_port, A_neg_shifted(42) => 
                           negative_inputs_13_42_port, A_neg_shifted(41) => 
                           negative_inputs_13_41_port, A_neg_shifted(40) => 
                           negative_inputs_13_40_port, A_neg_shifted(39) => 
                           negative_inputs_13_39_port, A_neg_shifted(38) => 
                           negative_inputs_13_38_port, A_neg_shifted(37) => 
                           negative_inputs_13_37_port, A_neg_shifted(36) => 
                           negative_inputs_13_36_port, A_neg_shifted(35) => 
                           negative_inputs_13_35_port, A_neg_shifted(34) => 
                           negative_inputs_13_34_port, A_neg_shifted(33) => 
                           negative_inputs_13_33_port, A_neg_shifted(32) => 
                           negative_inputs_13_32_port, A_neg_shifted(31) => 
                           negative_inputs_13_31_port, A_neg_shifted(30) => 
                           negative_inputs_13_30_port, A_neg_shifted(29) => 
                           negative_inputs_13_29_port, A_neg_shifted(28) => 
                           negative_inputs_13_28_port, A_neg_shifted(27) => 
                           negative_inputs_13_27_port, A_neg_shifted(26) => 
                           negative_inputs_13_26_port, A_neg_shifted(25) => 
                           negative_inputs_13_25_port, A_neg_shifted(24) => 
                           negative_inputs_13_24_port, A_neg_shifted(23) => 
                           negative_inputs_13_23_port, A_neg_shifted(22) => 
                           negative_inputs_13_22_port, A_neg_shifted(21) => 
                           negative_inputs_13_21_port, A_neg_shifted(20) => 
                           negative_inputs_13_20_port, A_neg_shifted(19) => 
                           negative_inputs_13_19_port, A_neg_shifted(18) => 
                           negative_inputs_13_18_port, A_neg_shifted(17) => 
                           negative_inputs_13_17_port, A_neg_shifted(16) => 
                           negative_inputs_13_16_port, A_neg_shifted(15) => 
                           negative_inputs_13_15_port, A_neg_shifted(14) => 
                           negative_inputs_13_14_port, A_neg_shifted(13) => 
                           negative_inputs_13_13_port, A_neg_shifted(12) => 
                           negative_inputs_13_12_port, A_neg_shifted(11) => 
                           negative_inputs_13_11_port, A_neg_shifted(10) => 
                           negative_inputs_13_10_port, A_neg_shifted(9) => 
                           negative_inputs_13_9_port, A_neg_shifted(8) => 
                           negative_inputs_13_8_port, A_neg_shifted(7) => 
                           negative_inputs_13_7_port, A_neg_shifted(6) => 
                           negative_inputs_13_6_port, A_neg_shifted(5) => 
                           negative_inputs_13_5_port, A_neg_shifted(4) => 
                           negative_inputs_13_4_port, A_neg_shifted(3) => 
                           negative_inputs_13_3_port, A_neg_shifted(2) => 
                           negative_inputs_13_2_port, A_neg_shifted(1) => 
                           negative_inputs_13_1_port, A_neg_shifted(0) => n8, 
                           Sel(2) => sel_6_2_port, Sel(1) => sel_6_1_port, 
                           Sel(0) => sel_6_0_port, Y(63) => 
                           MuxOutputs_6_63_port, Y(62) => MuxOutputs_6_62_port,
                           Y(61) => MuxOutputs_6_61_port, Y(60) => 
                           MuxOutputs_6_60_port, Y(59) => MuxOutputs_6_59_port,
                           Y(58) => MuxOutputs_6_58_port, Y(57) => 
                           MuxOutputs_6_57_port, Y(56) => MuxOutputs_6_56_port,
                           Y(55) => MuxOutputs_6_55_port, Y(54) => 
                           MuxOutputs_6_54_port, Y(53) => MuxOutputs_6_53_port,
                           Y(52) => MuxOutputs_6_52_port, Y(51) => 
                           MuxOutputs_6_51_port, Y(50) => MuxOutputs_6_50_port,
                           Y(49) => MuxOutputs_6_49_port, Y(48) => 
                           MuxOutputs_6_48_port, Y(47) => MuxOutputs_6_47_port,
                           Y(46) => MuxOutputs_6_46_port, Y(45) => 
                           MuxOutputs_6_45_port, Y(44) => MuxOutputs_6_44_port,
                           Y(43) => MuxOutputs_6_43_port, Y(42) => 
                           MuxOutputs_6_42_port, Y(41) => MuxOutputs_6_41_port,
                           Y(40) => MuxOutputs_6_40_port, Y(39) => 
                           MuxOutputs_6_39_port, Y(38) => MuxOutputs_6_38_port,
                           Y(37) => MuxOutputs_6_37_port, Y(36) => 
                           MuxOutputs_6_36_port, Y(35) => MuxOutputs_6_35_port,
                           Y(34) => MuxOutputs_6_34_port, Y(33) => 
                           MuxOutputs_6_33_port, Y(32) => MuxOutputs_6_32_port,
                           Y(31) => MuxOutputs_6_31_port, Y(30) => 
                           MuxOutputs_6_30_port, Y(29) => MuxOutputs_6_29_port,
                           Y(28) => MuxOutputs_6_28_port, Y(27) => 
                           MuxOutputs_6_27_port, Y(26) => MuxOutputs_6_26_port,
                           Y(25) => MuxOutputs_6_25_port, Y(24) => 
                           MuxOutputs_6_24_port, Y(23) => MuxOutputs_6_23_port,
                           Y(22) => MuxOutputs_6_22_port, Y(21) => 
                           MuxOutputs_6_21_port, Y(20) => MuxOutputs_6_20_port,
                           Y(19) => MuxOutputs_6_19_port, Y(18) => 
                           MuxOutputs_6_18_port, Y(17) => MuxOutputs_6_17_port,
                           Y(16) => MuxOutputs_6_16_port, Y(15) => 
                           MuxOutputs_6_15_port, Y(14) => MuxOutputs_6_14_port,
                           Y(13) => MuxOutputs_6_13_port, Y(12) => 
                           MuxOutputs_6_12_port, Y(11) => MuxOutputs_6_11_port,
                           Y(10) => MuxOutputs_6_10_port, Y(9) => 
                           MuxOutputs_6_9_port, Y(8) => MuxOutputs_6_8_port, 
                           Y(7) => MuxOutputs_6_7_port, Y(6) => 
                           MuxOutputs_6_6_port, Y(5) => MuxOutputs_6_5_port, 
                           Y(4) => MuxOutputs_6_4_port, Y(3) => 
                           MuxOutputs_6_3_port, Y(2) => MuxOutputs_6_2_port, 
                           Y(1) => MuxOutputs_6_1_port, Y(0) => 
                           MuxOutputs_6_0_port);
   encoderI_7 : encoder_25 port map( pieceofB(2) => B(15), pieceofB(1) => B(14)
                           , pieceofB(0) => B(13), sel(2) => sel_7_2_port, 
                           sel(1) => sel_7_1_port, sel(0) => sel_7_0_port);
   MUXI_7 : MUX51_MuxNbit64_25 port map( zeroSignal(63) => X_Logic0_port, 
                           zeroSignal(62) => X_Logic0_port, zeroSignal(61) => 
                           X_Logic0_port, zeroSignal(60) => X_Logic0_port, 
                           zeroSignal(59) => X_Logic0_port, zeroSignal(58) => 
                           X_Logic0_port, zeroSignal(57) => X_Logic0_port, 
                           zeroSignal(56) => X_Logic0_port, zeroSignal(55) => 
                           X_Logic0_port, zeroSignal(54) => X_Logic0_port, 
                           zeroSignal(53) => X_Logic0_port, zeroSignal(52) => 
                           X_Logic0_port, zeroSignal(51) => X_Logic0_port, 
                           zeroSignal(50) => X_Logic0_port, zeroSignal(49) => 
                           X_Logic0_port, zeroSignal(48) => X_Logic0_port, 
                           zeroSignal(47) => X_Logic0_port, zeroSignal(46) => 
                           X_Logic0_port, zeroSignal(45) => X_Logic0_port, 
                           zeroSignal(44) => X_Logic0_port, zeroSignal(43) => 
                           X_Logic0_port, zeroSignal(42) => X_Logic0_port, 
                           zeroSignal(41) => X_Logic0_port, zeroSignal(40) => 
                           X_Logic0_port, zeroSignal(39) => X_Logic0_port, 
                           zeroSignal(38) => X_Logic0_port, zeroSignal(37) => 
                           X_Logic0_port, zeroSignal(36) => X_Logic0_port, 
                           zeroSignal(35) => X_Logic0_port, zeroSignal(34) => 
                           X_Logic0_port, zeroSignal(33) => X_Logic0_port, 
                           zeroSignal(32) => X_Logic0_port, zeroSignal(31) => 
                           X_Logic0_port, zeroSignal(30) => X_Logic0_port, 
                           zeroSignal(29) => X_Logic0_port, zeroSignal(28) => 
                           X_Logic0_port, zeroSignal(27) => X_Logic0_port, 
                           zeroSignal(26) => X_Logic0_port, zeroSignal(25) => 
                           X_Logic0_port, zeroSignal(24) => X_Logic0_port, 
                           zeroSignal(23) => X_Logic0_port, zeroSignal(22) => 
                           X_Logic0_port, zeroSignal(21) => X_Logic0_port, 
                           zeroSignal(20) => X_Logic0_port, zeroSignal(19) => 
                           X_Logic0_port, zeroSignal(18) => X_Logic0_port, 
                           zeroSignal(17) => X_Logic0_port, zeroSignal(16) => 
                           X_Logic0_port, zeroSignal(15) => X_Logic0_port, 
                           zeroSignal(14) => X_Logic0_port, zeroSignal(13) => 
                           X_Logic0_port, zeroSignal(12) => X_Logic0_port, 
                           zeroSignal(11) => X_Logic0_port, zeroSignal(10) => 
                           X_Logic0_port, zeroSignal(9) => X_Logic0_port, 
                           zeroSignal(8) => X_Logic0_port, zeroSignal(7) => 
                           X_Logic0_port, zeroSignal(6) => X_Logic0_port, 
                           zeroSignal(5) => X_Logic0_port, zeroSignal(4) => 
                           X_Logic0_port, zeroSignal(3) => X_Logic0_port, 
                           zeroSignal(2) => X_Logic0_port, zeroSignal(1) => 
                           X_Logic0_port, zeroSignal(0) => X_Logic0_port, 
                           A_signal(63) => positive_inputs_14_63_port, 
                           A_signal(62) => positive_inputs_14_62_port, 
                           A_signal(61) => positive_inputs_14_61_port, 
                           A_signal(60) => positive_inputs_14_60_port, 
                           A_signal(59) => positive_inputs_14_59_port, 
                           A_signal(58) => positive_inputs_14_58_port, 
                           A_signal(57) => positive_inputs_14_57_port, 
                           A_signal(56) => positive_inputs_14_56_port, 
                           A_signal(55) => positive_inputs_14_55_port, 
                           A_signal(54) => positive_inputs_14_54_port, 
                           A_signal(53) => positive_inputs_14_53_port, 
                           A_signal(52) => positive_inputs_14_52_port, 
                           A_signal(51) => positive_inputs_14_51_port, 
                           A_signal(50) => positive_inputs_14_50_port, 
                           A_signal(49) => positive_inputs_14_49_port, 
                           A_signal(48) => positive_inputs_14_48_port, 
                           A_signal(47) => n27, A_signal(46) => 
                           positive_inputs_14_46_port, A_signal(45) => 
                           positive_inputs_14_45_port, A_signal(44) => 
                           positive_inputs_14_44_port, A_signal(43) => 
                           positive_inputs_14_43_port, A_signal(42) => 
                           positive_inputs_14_42_port, A_signal(41) => 
                           positive_inputs_14_41_port, A_signal(40) => 
                           positive_inputs_14_40_port, A_signal(39) => 
                           positive_inputs_14_39_port, A_signal(38) => 
                           positive_inputs_14_38_port, A_signal(37) => 
                           positive_inputs_14_37_port, A_signal(36) => 
                           positive_inputs_14_36_port, A_signal(35) => 
                           positive_inputs_14_35_port, A_signal(34) => 
                           positive_inputs_14_34_port, A_signal(33) => 
                           positive_inputs_14_33_port, A_signal(32) => 
                           positive_inputs_14_32_port, A_signal(31) => 
                           positive_inputs_14_31_port, A_signal(30) => 
                           positive_inputs_14_30_port, A_signal(29) => 
                           positive_inputs_14_29_port, A_signal(28) => 
                           positive_inputs_14_28_port, A_signal(27) => 
                           positive_inputs_14_27_port, A_signal(26) => 
                           positive_inputs_14_26_port, A_signal(25) => 
                           positive_inputs_14_25_port, A_signal(24) => 
                           positive_inputs_14_24_port, A_signal(23) => 
                           positive_inputs_14_23_port, A_signal(22) => 
                           positive_inputs_14_22_port, A_signal(21) => 
                           positive_inputs_14_21_port, A_signal(20) => 
                           positive_inputs_14_20_port, A_signal(19) => 
                           positive_inputs_14_19_port, A_signal(18) => 
                           positive_inputs_14_18_port, A_signal(17) => 
                           positive_inputs_14_17_port, A_signal(16) => 
                           positive_inputs_14_16_port, A_signal(15) => 
                           positive_inputs_14_15_port, A_signal(14) => 
                           positive_inputs_14_14_port, A_signal(13) => 
                           positive_inputs_14_13_port, A_signal(12) => 
                           positive_inputs_14_12_port, A_signal(11) => 
                           positive_inputs_14_11_port, A_signal(10) => 
                           positive_inputs_14_10_port, A_signal(9) => 
                           positive_inputs_14_9_port, A_signal(8) => 
                           positive_inputs_14_8_port, A_signal(7) => 
                           positive_inputs_14_7_port, A_signal(6) => 
                           positive_inputs_14_6_port, A_signal(5) => 
                           positive_inputs_14_5_port, A_signal(4) => 
                           positive_inputs_14_4_port, A_signal(3) => 
                           positive_inputs_14_3_port, A_signal(2) => 
                           positive_inputs_14_2_port, A_signal(1) => 
                           positive_inputs_14_1_port, A_signal(0) => n8, 
                           A_neg(63) => negative_inputs_14_63_port, A_neg(62) 
                           => negative_inputs_14_62_port, A_neg(61) => 
                           negative_inputs_14_61_port, A_neg(60) => 
                           negative_inputs_14_60_port, A_neg(59) => 
                           negative_inputs_14_59_port, A_neg(58) => 
                           negative_inputs_14_58_port, A_neg(57) => 
                           negative_inputs_14_57_port, A_neg(56) => 
                           negative_inputs_14_56_port, A_neg(55) => 
                           negative_inputs_14_55_port, A_neg(54) => 
                           negative_inputs_14_54_port, A_neg(53) => 
                           negative_inputs_14_53_port, A_neg(52) => 
                           negative_inputs_14_52_port, A_neg(51) => 
                           negative_inputs_14_51_port, A_neg(50) => 
                           negative_inputs_14_50_port, A_neg(49) => 
                           negative_inputs_14_49_port, A_neg(48) => 
                           negative_inputs_14_48_port, A_neg(47) => n109, 
                           A_neg(46) => negative_inputs_14_46_port, A_neg(45) 
                           => negative_inputs_14_45_port, A_neg(44) => 
                           negative_inputs_14_44_port, A_neg(43) => 
                           negative_inputs_14_43_port, A_neg(42) => 
                           negative_inputs_14_42_port, A_neg(41) => 
                           negative_inputs_14_41_port, A_neg(40) => 
                           negative_inputs_14_40_port, A_neg(39) => 
                           negative_inputs_14_39_port, A_neg(38) => 
                           negative_inputs_14_38_port, A_neg(37) => 
                           negative_inputs_14_37_port, A_neg(36) => 
                           negative_inputs_14_36_port, A_neg(35) => 
                           negative_inputs_14_35_port, A_neg(34) => 
                           negative_inputs_14_34_port, A_neg(33) => 
                           negative_inputs_14_33_port, A_neg(32) => 
                           negative_inputs_14_32_port, A_neg(31) => 
                           negative_inputs_14_31_port, A_neg(30) => 
                           negative_inputs_14_30_port, A_neg(29) => 
                           negative_inputs_14_29_port, A_neg(28) => 
                           negative_inputs_14_28_port, A_neg(27) => 
                           negative_inputs_14_27_port, A_neg(26) => 
                           negative_inputs_14_26_port, A_neg(25) => 
                           negative_inputs_14_25_port, A_neg(24) => 
                           negative_inputs_14_24_port, A_neg(23) => 
                           negative_inputs_14_23_port, A_neg(22) => 
                           negative_inputs_14_22_port, A_neg(21) => 
                           negative_inputs_14_21_port, A_neg(20) => 
                           negative_inputs_14_20_port, A_neg(19) => 
                           negative_inputs_14_19_port, A_neg(18) => 
                           negative_inputs_14_18_port, A_neg(17) => 
                           negative_inputs_14_17_port, A_neg(16) => 
                           negative_inputs_14_16_port, A_neg(15) => 
                           negative_inputs_14_15_port, A_neg(14) => 
                           negative_inputs_14_14_port, A_neg(13) => 
                           negative_inputs_14_13_port, A_neg(12) => 
                           negative_inputs_14_12_port, A_neg(11) => 
                           negative_inputs_14_11_port, A_neg(10) => 
                           negative_inputs_14_10_port, A_neg(9) => 
                           negative_inputs_14_9_port, A_neg(8) => 
                           negative_inputs_14_8_port, A_neg(7) => 
                           negative_inputs_14_7_port, A_neg(6) => 
                           negative_inputs_14_6_port, A_neg(5) => 
                           negative_inputs_14_5_port, A_neg(4) => 
                           negative_inputs_14_4_port, A_neg(3) => 
                           negative_inputs_14_3_port, A_neg(2) => 
                           negative_inputs_14_2_port, A_neg(1) => 
                           negative_inputs_14_1_port, A_neg(0) => n8, 
                           A_shifted(63) => positive_inputs_15_63_port, 
                           A_shifted(62) => positive_inputs_15_62_port, 
                           A_shifted(61) => positive_inputs_15_61_port, 
                           A_shifted(60) => positive_inputs_15_60_port, 
                           A_shifted(59) => positive_inputs_15_59_port, 
                           A_shifted(58) => positive_inputs_15_58_port, 
                           A_shifted(57) => positive_inputs_15_57_port, 
                           A_shifted(56) => positive_inputs_15_56_port, 
                           A_shifted(55) => positive_inputs_15_55_port, 
                           A_shifted(54) => positive_inputs_15_54_port, 
                           A_shifted(53) => positive_inputs_15_53_port, 
                           A_shifted(52) => positive_inputs_15_52_port, 
                           A_shifted(51) => positive_inputs_15_51_port, 
                           A_shifted(50) => positive_inputs_15_50_port, 
                           A_shifted(49) => positive_inputs_15_49_port, 
                           A_shifted(48) => positive_inputs_15_48_port, 
                           A_shifted(47) => n26, A_shifted(46) => n25, 
                           A_shifted(45) => n181, A_shifted(44) => n179, 
                           A_shifted(43) => n177, A_shifted(42) => n175, 
                           A_shifted(41) => n173, A_shifted(40) => n171, 
                           A_shifted(39) => n169, A_shifted(38) => n167, 
                           A_shifted(37) => n165, A_shifted(36) => n163, 
                           A_shifted(35) => n161, A_shifted(34) => n159, 
                           A_shifted(33) => n157, A_shifted(32) => n155, 
                           A_shifted(31) => n153, A_shifted(30) => n151, 
                           A_shifted(29) => n149, A_shifted(28) => n147, 
                           A_shifted(27) => n145, A_shifted(26) => n143, 
                           A_shifted(25) => n141, A_shifted(24) => n139, 
                           A_shifted(23) => n137, A_shifted(22) => n135, 
                           A_shifted(21) => n133, A_shifted(20) => n131, 
                           A_shifted(19) => n129, A_shifted(18) => n127, 
                           A_shifted(17) => n125, A_shifted(16) => n123, 
                           A_shifted(15) => n121, A_shifted(14) => 
                           positive_inputs_15_14_port, A_shifted(13) => 
                           positive_inputs_15_13_port, A_shifted(12) => 
                           positive_inputs_15_12_port, A_shifted(11) => 
                           positive_inputs_15_11_port, A_shifted(10) => 
                           positive_inputs_15_10_port, A_shifted(9) => 
                           positive_inputs_15_9_port, A_shifted(8) => 
                           positive_inputs_15_8_port, A_shifted(7) => 
                           positive_inputs_15_7_port, A_shifted(6) => 
                           positive_inputs_15_6_port, A_shifted(5) => 
                           positive_inputs_15_5_port, A_shifted(4) => 
                           positive_inputs_15_4_port, A_shifted(3) => 
                           positive_inputs_15_3_port, A_shifted(2) => 
                           positive_inputs_15_2_port, A_shifted(1) => 
                           positive_inputs_15_1_port, A_shifted(0) => n8, 
                           A_neg_shifted(63) => negative_inputs_15_63_port, 
                           A_neg_shifted(62) => negative_inputs_15_62_port, 
                           A_neg_shifted(61) => negative_inputs_15_61_port, 
                           A_neg_shifted(60) => negative_inputs_15_60_port, 
                           A_neg_shifted(59) => negative_inputs_15_59_port, 
                           A_neg_shifted(58) => negative_inputs_15_58_port, 
                           A_neg_shifted(57) => negative_inputs_15_57_port, 
                           A_neg_shifted(56) => negative_inputs_15_56_port, 
                           A_neg_shifted(55) => negative_inputs_15_55_port, 
                           A_neg_shifted(54) => negative_inputs_15_54_port, 
                           A_neg_shifted(53) => negative_inputs_15_53_port, 
                           A_neg_shifted(52) => negative_inputs_15_52_port, 
                           A_neg_shifted(51) => negative_inputs_15_51_port, 
                           A_neg_shifted(50) => negative_inputs_15_50_port, 
                           A_neg_shifted(49) => negative_inputs_15_49_port, 
                           A_neg_shifted(48) => negative_inputs_15_48_port, 
                           A_neg_shifted(47) => n107, A_neg_shifted(46) => n105
                           , A_neg_shifted(45) => n103, A_neg_shifted(44) => 
                           n101, A_neg_shifted(43) => n99, A_neg_shifted(42) =>
                           n97, A_neg_shifted(41) => n95, A_neg_shifted(40) => 
                           n93, A_neg_shifted(39) => n91, A_neg_shifted(38) => 
                           n89, A_neg_shifted(37) => n87, A_neg_shifted(36) => 
                           n85, A_neg_shifted(35) => n83, A_neg_shifted(34) => 
                           n81, A_neg_shifted(33) => n79, A_neg_shifted(32) => 
                           n77, A_neg_shifted(31) => n75, A_neg_shifted(30) => 
                           n73, A_neg_shifted(29) => n71, A_neg_shifted(28) => 
                           n69, A_neg_shifted(27) => n67, A_neg_shifted(26) => 
                           n65, A_neg_shifted(25) => n63, A_neg_shifted(24) => 
                           n61, A_neg_shifted(23) => n59, A_neg_shifted(22) => 
                           n57, A_neg_shifted(21) => n55, A_neg_shifted(20) => 
                           n53, A_neg_shifted(19) => n51, A_neg_shifted(18) => 
                           n49, A_neg_shifted(17) => n47, A_neg_shifted(16) => 
                           n45, A_neg_shifted(15) => n43, A_neg_shifted(14) => 
                           negative_inputs_15_14_port, A_neg_shifted(13) => 
                           negative_inputs_15_13_port, A_neg_shifted(12) => 
                           negative_inputs_15_12_port, A_neg_shifted(11) => 
                           negative_inputs_15_11_port, A_neg_shifted(10) => 
                           negative_inputs_15_10_port, A_neg_shifted(9) => 
                           negative_inputs_15_9_port, A_neg_shifted(8) => 
                           negative_inputs_15_8_port, A_neg_shifted(7) => 
                           negative_inputs_15_7_port, A_neg_shifted(6) => 
                           negative_inputs_15_6_port, A_neg_shifted(5) => 
                           negative_inputs_15_5_port, A_neg_shifted(4) => 
                           negative_inputs_15_4_port, A_neg_shifted(3) => 
                           negative_inputs_15_3_port, A_neg_shifted(2) => 
                           negative_inputs_15_2_port, A_neg_shifted(1) => 
                           negative_inputs_15_1_port, A_neg_shifted(0) => n8, 
                           Sel(2) => sel_7_2_port, Sel(1) => sel_7_1_port, 
                           Sel(0) => sel_7_0_port, Y(63) => 
                           MuxOutputs_7_63_port, Y(62) => MuxOutputs_7_62_port,
                           Y(61) => MuxOutputs_7_61_port, Y(60) => 
                           MuxOutputs_7_60_port, Y(59) => MuxOutputs_7_59_port,
                           Y(58) => MuxOutputs_7_58_port, Y(57) => 
                           MuxOutputs_7_57_port, Y(56) => MuxOutputs_7_56_port,
                           Y(55) => MuxOutputs_7_55_port, Y(54) => 
                           MuxOutputs_7_54_port, Y(53) => MuxOutputs_7_53_port,
                           Y(52) => MuxOutputs_7_52_port, Y(51) => 
                           MuxOutputs_7_51_port, Y(50) => MuxOutputs_7_50_port,
                           Y(49) => MuxOutputs_7_49_port, Y(48) => 
                           MuxOutputs_7_48_port, Y(47) => MuxOutputs_7_47_port,
                           Y(46) => MuxOutputs_7_46_port, Y(45) => 
                           MuxOutputs_7_45_port, Y(44) => MuxOutputs_7_44_port,
                           Y(43) => MuxOutputs_7_43_port, Y(42) => 
                           MuxOutputs_7_42_port, Y(41) => MuxOutputs_7_41_port,
                           Y(40) => MuxOutputs_7_40_port, Y(39) => 
                           MuxOutputs_7_39_port, Y(38) => MuxOutputs_7_38_port,
                           Y(37) => MuxOutputs_7_37_port, Y(36) => 
                           MuxOutputs_7_36_port, Y(35) => MuxOutputs_7_35_port,
                           Y(34) => MuxOutputs_7_34_port, Y(33) => 
                           MuxOutputs_7_33_port, Y(32) => MuxOutputs_7_32_port,
                           Y(31) => MuxOutputs_7_31_port, Y(30) => 
                           MuxOutputs_7_30_port, Y(29) => MuxOutputs_7_29_port,
                           Y(28) => MuxOutputs_7_28_port, Y(27) => 
                           MuxOutputs_7_27_port, Y(26) => MuxOutputs_7_26_port,
                           Y(25) => MuxOutputs_7_25_port, Y(24) => 
                           MuxOutputs_7_24_port, Y(23) => MuxOutputs_7_23_port,
                           Y(22) => MuxOutputs_7_22_port, Y(21) => 
                           MuxOutputs_7_21_port, Y(20) => MuxOutputs_7_20_port,
                           Y(19) => MuxOutputs_7_19_port, Y(18) => 
                           MuxOutputs_7_18_port, Y(17) => MuxOutputs_7_17_port,
                           Y(16) => MuxOutputs_7_16_port, Y(15) => 
                           MuxOutputs_7_15_port, Y(14) => MuxOutputs_7_14_port,
                           Y(13) => MuxOutputs_7_13_port, Y(12) => 
                           MuxOutputs_7_12_port, Y(11) => MuxOutputs_7_11_port,
                           Y(10) => MuxOutputs_7_10_port, Y(9) => 
                           MuxOutputs_7_9_port, Y(8) => MuxOutputs_7_8_port, 
                           Y(7) => MuxOutputs_7_7_port, Y(6) => 
                           MuxOutputs_7_6_port, Y(5) => MuxOutputs_7_5_port, 
                           Y(4) => MuxOutputs_7_4_port, Y(3) => 
                           MuxOutputs_7_3_port, Y(2) => MuxOutputs_7_2_port, 
                           Y(1) => MuxOutputs_7_1_port, Y(0) => 
                           MuxOutputs_7_0_port);
   encoderI_8 : encoder_24 port map( pieceofB(2) => B(17), pieceofB(1) => B(16)
                           , pieceofB(0) => B(15), sel(2) => sel_8_2_port, 
                           sel(1) => sel_8_1_port, sel(0) => sel_8_0_port);
   MUXI_8 : MUX51_MuxNbit64_24 port map( zeroSignal(63) => X_Logic0_port, 
                           zeroSignal(62) => X_Logic0_port, zeroSignal(61) => 
                           X_Logic0_port, zeroSignal(60) => X_Logic0_port, 
                           zeroSignal(59) => X_Logic0_port, zeroSignal(58) => 
                           X_Logic0_port, zeroSignal(57) => X_Logic0_port, 
                           zeroSignal(56) => X_Logic0_port, zeroSignal(55) => 
                           X_Logic0_port, zeroSignal(54) => X_Logic0_port, 
                           zeroSignal(53) => X_Logic0_port, zeroSignal(52) => 
                           X_Logic0_port, zeroSignal(51) => X_Logic0_port, 
                           zeroSignal(50) => X_Logic0_port, zeroSignal(49) => 
                           X_Logic0_port, zeroSignal(48) => X_Logic0_port, 
                           zeroSignal(47) => X_Logic0_port, zeroSignal(46) => 
                           X_Logic0_port, zeroSignal(45) => X_Logic0_port, 
                           zeroSignal(44) => X_Logic0_port, zeroSignal(43) => 
                           X_Logic0_port, zeroSignal(42) => X_Logic0_port, 
                           zeroSignal(41) => X_Logic0_port, zeroSignal(40) => 
                           X_Logic0_port, zeroSignal(39) => X_Logic0_port, 
                           zeroSignal(38) => X_Logic0_port, zeroSignal(37) => 
                           X_Logic0_port, zeroSignal(36) => X_Logic0_port, 
                           zeroSignal(35) => X_Logic0_port, zeroSignal(34) => 
                           X_Logic0_port, zeroSignal(33) => X_Logic0_port, 
                           zeroSignal(32) => X_Logic0_port, zeroSignal(31) => 
                           X_Logic0_port, zeroSignal(30) => X_Logic0_port, 
                           zeroSignal(29) => X_Logic0_port, zeroSignal(28) => 
                           X_Logic0_port, zeroSignal(27) => X_Logic0_port, 
                           zeroSignal(26) => X_Logic0_port, zeroSignal(25) => 
                           X_Logic0_port, zeroSignal(24) => X_Logic0_port, 
                           zeroSignal(23) => X_Logic0_port, zeroSignal(22) => 
                           X_Logic0_port, zeroSignal(21) => X_Logic0_port, 
                           zeroSignal(20) => X_Logic0_port, zeroSignal(19) => 
                           X_Logic0_port, zeroSignal(18) => X_Logic0_port, 
                           zeroSignal(17) => X_Logic0_port, zeroSignal(16) => 
                           X_Logic0_port, zeroSignal(15) => X_Logic0_port, 
                           zeroSignal(14) => X_Logic0_port, zeroSignal(13) => 
                           X_Logic0_port, zeroSignal(12) => X_Logic0_port, 
                           zeroSignal(11) => X_Logic0_port, zeroSignal(10) => 
                           X_Logic0_port, zeroSignal(9) => X_Logic0_port, 
                           zeroSignal(8) => X_Logic0_port, zeroSignal(7) => 
                           X_Logic0_port, zeroSignal(6) => X_Logic0_port, 
                           zeroSignal(5) => X_Logic0_port, zeroSignal(4) => 
                           X_Logic0_port, zeroSignal(3) => X_Logic0_port, 
                           zeroSignal(2) => X_Logic0_port, zeroSignal(1) => 
                           X_Logic0_port, zeroSignal(0) => X_Logic0_port, 
                           A_signal(63) => positive_inputs_16_63_port, 
                           A_signal(62) => positive_inputs_16_62_port, 
                           A_signal(61) => positive_inputs_16_61_port, 
                           A_signal(60) => positive_inputs_16_60_port, 
                           A_signal(59) => positive_inputs_16_59_port, 
                           A_signal(58) => positive_inputs_16_58_port, 
                           A_signal(57) => positive_inputs_16_57_port, 
                           A_signal(56) => positive_inputs_16_56_port, 
                           A_signal(55) => positive_inputs_16_55_port, 
                           A_signal(54) => positive_inputs_16_54_port, 
                           A_signal(53) => positive_inputs_16_53_port, 
                           A_signal(52) => positive_inputs_16_52_port, 
                           A_signal(51) => positive_inputs_16_51_port, 
                           A_signal(50) => positive_inputs_16_50_port, 
                           A_signal(49) => positive_inputs_16_49_port, 
                           A_signal(48) => positive_inputs_16_48_port, 
                           A_signal(47) => positive_inputs_16_47_port, 
                           A_signal(46) => positive_inputs_16_46_port, 
                           A_signal(45) => positive_inputs_16_45_port, 
                           A_signal(44) => positive_inputs_16_44_port, 
                           A_signal(43) => positive_inputs_16_43_port, 
                           A_signal(42) => positive_inputs_16_42_port, 
                           A_signal(41) => positive_inputs_16_41_port, 
                           A_signal(40) => positive_inputs_16_40_port, 
                           A_signal(39) => positive_inputs_16_39_port, 
                           A_signal(38) => positive_inputs_16_38_port, 
                           A_signal(37) => positive_inputs_16_37_port, 
                           A_signal(36) => positive_inputs_16_36_port, 
                           A_signal(35) => positive_inputs_16_35_port, 
                           A_signal(34) => positive_inputs_16_34_port, 
                           A_signal(33) => positive_inputs_16_33_port, 
                           A_signal(32) => positive_inputs_16_32_port, 
                           A_signal(31) => positive_inputs_16_31_port, 
                           A_signal(30) => positive_inputs_16_30_port, 
                           A_signal(29) => positive_inputs_16_29_port, 
                           A_signal(28) => positive_inputs_16_28_port, 
                           A_signal(27) => positive_inputs_16_27_port, 
                           A_signal(26) => positive_inputs_16_26_port, 
                           A_signal(25) => positive_inputs_16_25_port, 
                           A_signal(24) => positive_inputs_16_24_port, 
                           A_signal(23) => positive_inputs_16_23_port, 
                           A_signal(22) => positive_inputs_16_22_port, 
                           A_signal(21) => positive_inputs_16_21_port, 
                           A_signal(20) => positive_inputs_16_20_port, 
                           A_signal(19) => positive_inputs_16_19_port, 
                           A_signal(18) => positive_inputs_16_18_port, 
                           A_signal(17) => positive_inputs_16_17_port, 
                           A_signal(16) => positive_inputs_16_16_port, 
                           A_signal(15) => positive_inputs_16_15_port, 
                           A_signal(14) => positive_inputs_16_14_port, 
                           A_signal(13) => positive_inputs_16_13_port, 
                           A_signal(12) => positive_inputs_16_12_port, 
                           A_signal(11) => positive_inputs_16_11_port, 
                           A_signal(10) => positive_inputs_16_10_port, 
                           A_signal(9) => positive_inputs_16_9_port, 
                           A_signal(8) => positive_inputs_16_8_port, 
                           A_signal(7) => positive_inputs_16_7_port, 
                           A_signal(6) => positive_inputs_16_6_port, 
                           A_signal(5) => positive_inputs_16_5_port, 
                           A_signal(4) => positive_inputs_16_4_port, 
                           A_signal(3) => positive_inputs_16_3_port, 
                           A_signal(2) => positive_inputs_16_2_port, 
                           A_signal(1) => positive_inputs_16_1_port, 
                           A_signal(0) => n8, A_neg(63) => 
                           negative_inputs_16_63_port, A_neg(62) => 
                           negative_inputs_16_62_port, A_neg(61) => 
                           negative_inputs_16_61_port, A_neg(60) => 
                           negative_inputs_16_60_port, A_neg(59) => 
                           negative_inputs_16_59_port, A_neg(58) => 
                           negative_inputs_16_58_port, A_neg(57) => 
                           negative_inputs_16_57_port, A_neg(56) => 
                           negative_inputs_16_56_port, A_neg(55) => 
                           negative_inputs_16_55_port, A_neg(54) => 
                           negative_inputs_16_54_port, A_neg(53) => 
                           negative_inputs_16_53_port, A_neg(52) => 
                           negative_inputs_16_52_port, A_neg(51) => 
                           negative_inputs_16_51_port, A_neg(50) => 
                           negative_inputs_16_50_port, A_neg(49) => 
                           negative_inputs_16_49_port, A_neg(48) => 
                           negative_inputs_16_48_port, A_neg(47) => 
                           negative_inputs_16_47_port, A_neg(46) => 
                           negative_inputs_16_46_port, A_neg(45) => 
                           negative_inputs_16_45_port, A_neg(44) => 
                           negative_inputs_16_44_port, A_neg(43) => 
                           negative_inputs_16_43_port, A_neg(42) => 
                           negative_inputs_16_42_port, A_neg(41) => 
                           negative_inputs_16_41_port, A_neg(40) => 
                           negative_inputs_16_40_port, A_neg(39) => 
                           negative_inputs_16_39_port, A_neg(38) => 
                           negative_inputs_16_38_port, A_neg(37) => 
                           negative_inputs_16_37_port, A_neg(36) => 
                           negative_inputs_16_36_port, A_neg(35) => 
                           negative_inputs_16_35_port, A_neg(34) => 
                           negative_inputs_16_34_port, A_neg(33) => 
                           negative_inputs_16_33_port, A_neg(32) => 
                           negative_inputs_16_32_port, A_neg(31) => 
                           negative_inputs_16_31_port, A_neg(30) => 
                           negative_inputs_16_30_port, A_neg(29) => 
                           negative_inputs_16_29_port, A_neg(28) => 
                           negative_inputs_16_28_port, A_neg(27) => 
                           negative_inputs_16_27_port, A_neg(26) => 
                           negative_inputs_16_26_port, A_neg(25) => 
                           negative_inputs_16_25_port, A_neg(24) => 
                           negative_inputs_16_24_port, A_neg(23) => 
                           negative_inputs_16_23_port, A_neg(22) => 
                           negative_inputs_16_22_port, A_neg(21) => 
                           negative_inputs_16_21_port, A_neg(20) => 
                           negative_inputs_16_20_port, A_neg(19) => 
                           negative_inputs_16_19_port, A_neg(18) => 
                           negative_inputs_16_18_port, A_neg(17) => 
                           negative_inputs_16_17_port, A_neg(16) => 
                           negative_inputs_16_16_port, A_neg(15) => 
                           negative_inputs_16_15_port, A_neg(14) => 
                           negative_inputs_16_14_port, A_neg(13) => 
                           negative_inputs_16_13_port, A_neg(12) => 
                           negative_inputs_16_12_port, A_neg(11) => 
                           negative_inputs_16_11_port, A_neg(10) => 
                           negative_inputs_16_10_port, A_neg(9) => 
                           negative_inputs_16_9_port, A_neg(8) => 
                           negative_inputs_16_8_port, A_neg(7) => 
                           negative_inputs_16_7_port, A_neg(6) => 
                           negative_inputs_16_6_port, A_neg(5) => 
                           negative_inputs_16_5_port, A_neg(4) => 
                           negative_inputs_16_4_port, A_neg(3) => 
                           negative_inputs_16_3_port, A_neg(2) => 
                           negative_inputs_16_2_port, A_neg(1) => 
                           negative_inputs_16_1_port, A_neg(0) => n8, 
                           A_shifted(63) => positive_inputs_17_63_port, 
                           A_shifted(62) => positive_inputs_17_62_port, 
                           A_shifted(61) => positive_inputs_17_61_port, 
                           A_shifted(60) => positive_inputs_17_60_port, 
                           A_shifted(59) => positive_inputs_17_59_port, 
                           A_shifted(58) => positive_inputs_17_58_port, 
                           A_shifted(57) => positive_inputs_17_57_port, 
                           A_shifted(56) => positive_inputs_17_56_port, 
                           A_shifted(55) => positive_inputs_17_55_port, 
                           A_shifted(54) => positive_inputs_17_54_port, 
                           A_shifted(53) => positive_inputs_17_53_port, 
                           A_shifted(52) => positive_inputs_17_52_port, 
                           A_shifted(51) => positive_inputs_17_51_port, 
                           A_shifted(50) => positive_inputs_17_50_port, 
                           A_shifted(49) => positive_inputs_17_49_port, 
                           A_shifted(48) => positive_inputs_17_48_port, 
                           A_shifted(47) => positive_inputs_17_47_port, 
                           A_shifted(46) => positive_inputs_17_46_port, 
                           A_shifted(45) => positive_inputs_17_45_port, 
                           A_shifted(44) => positive_inputs_17_44_port, 
                           A_shifted(43) => positive_inputs_17_43_port, 
                           A_shifted(42) => positive_inputs_17_42_port, 
                           A_shifted(41) => positive_inputs_17_41_port, 
                           A_shifted(40) => positive_inputs_17_40_port, 
                           A_shifted(39) => positive_inputs_17_39_port, 
                           A_shifted(38) => positive_inputs_17_38_port, 
                           A_shifted(37) => positive_inputs_17_37_port, 
                           A_shifted(36) => positive_inputs_17_36_port, 
                           A_shifted(35) => positive_inputs_17_35_port, 
                           A_shifted(34) => positive_inputs_17_34_port, 
                           A_shifted(33) => positive_inputs_17_33_port, 
                           A_shifted(32) => positive_inputs_17_32_port, 
                           A_shifted(31) => positive_inputs_17_31_port, 
                           A_shifted(30) => positive_inputs_17_30_port, 
                           A_shifted(29) => positive_inputs_17_29_port, 
                           A_shifted(28) => positive_inputs_17_28_port, 
                           A_shifted(27) => positive_inputs_17_27_port, 
                           A_shifted(26) => positive_inputs_17_26_port, 
                           A_shifted(25) => positive_inputs_17_25_port, 
                           A_shifted(24) => positive_inputs_17_24_port, 
                           A_shifted(23) => positive_inputs_17_23_port, 
                           A_shifted(22) => positive_inputs_17_22_port, 
                           A_shifted(21) => positive_inputs_17_21_port, 
                           A_shifted(20) => positive_inputs_17_20_port, 
                           A_shifted(19) => positive_inputs_17_19_port, 
                           A_shifted(18) => positive_inputs_17_18_port, 
                           A_shifted(17) => positive_inputs_17_17_port, 
                           A_shifted(16) => positive_inputs_17_16_port, 
                           A_shifted(15) => positive_inputs_17_15_port, 
                           A_shifted(14) => positive_inputs_17_14_port, 
                           A_shifted(13) => positive_inputs_17_13_port, 
                           A_shifted(12) => positive_inputs_17_12_port, 
                           A_shifted(11) => positive_inputs_17_11_port, 
                           A_shifted(10) => positive_inputs_17_10_port, 
                           A_shifted(9) => positive_inputs_17_9_port, 
                           A_shifted(8) => positive_inputs_17_8_port, 
                           A_shifted(7) => positive_inputs_17_7_port, 
                           A_shifted(6) => positive_inputs_17_6_port, 
                           A_shifted(5) => positive_inputs_17_5_port, 
                           A_shifted(4) => positive_inputs_17_4_port, 
                           A_shifted(3) => positive_inputs_17_3_port, 
                           A_shifted(2) => positive_inputs_17_2_port, 
                           A_shifted(1) => positive_inputs_17_1_port, 
                           A_shifted(0) => n8, A_neg_shifted(63) => 
                           negative_inputs_17_63_port, A_neg_shifted(62) => 
                           negative_inputs_17_62_port, A_neg_shifted(61) => 
                           negative_inputs_17_61_port, A_neg_shifted(60) => 
                           negative_inputs_17_60_port, A_neg_shifted(59) => 
                           negative_inputs_17_59_port, A_neg_shifted(58) => 
                           negative_inputs_17_58_port, A_neg_shifted(57) => 
                           negative_inputs_17_57_port, A_neg_shifted(56) => 
                           negative_inputs_17_56_port, A_neg_shifted(55) => 
                           negative_inputs_17_55_port, A_neg_shifted(54) => 
                           negative_inputs_17_54_port, A_neg_shifted(53) => 
                           negative_inputs_17_53_port, A_neg_shifted(52) => 
                           negative_inputs_17_52_port, A_neg_shifted(51) => 
                           negative_inputs_17_51_port, A_neg_shifted(50) => 
                           negative_inputs_17_50_port, A_neg_shifted(49) => 
                           negative_inputs_17_49_port, A_neg_shifted(48) => 
                           negative_inputs_17_48_port, A_neg_shifted(47) => 
                           negative_inputs_17_47_port, A_neg_shifted(46) => 
                           negative_inputs_17_46_port, A_neg_shifted(45) => 
                           negative_inputs_17_45_port, A_neg_shifted(44) => 
                           negative_inputs_17_44_port, A_neg_shifted(43) => 
                           negative_inputs_17_43_port, A_neg_shifted(42) => 
                           negative_inputs_17_42_port, A_neg_shifted(41) => 
                           negative_inputs_17_41_port, A_neg_shifted(40) => 
                           negative_inputs_17_40_port, A_neg_shifted(39) => 
                           negative_inputs_17_39_port, A_neg_shifted(38) => 
                           negative_inputs_17_38_port, A_neg_shifted(37) => 
                           negative_inputs_17_37_port, A_neg_shifted(36) => 
                           negative_inputs_17_36_port, A_neg_shifted(35) => 
                           negative_inputs_17_35_port, A_neg_shifted(34) => 
                           negative_inputs_17_34_port, A_neg_shifted(33) => 
                           negative_inputs_17_33_port, A_neg_shifted(32) => 
                           negative_inputs_17_32_port, A_neg_shifted(31) => 
                           negative_inputs_17_31_port, A_neg_shifted(30) => 
                           negative_inputs_17_30_port, A_neg_shifted(29) => 
                           negative_inputs_17_29_port, A_neg_shifted(28) => 
                           negative_inputs_17_28_port, A_neg_shifted(27) => 
                           negative_inputs_17_27_port, A_neg_shifted(26) => 
                           negative_inputs_17_26_port, A_neg_shifted(25) => 
                           negative_inputs_17_25_port, A_neg_shifted(24) => 
                           negative_inputs_17_24_port, A_neg_shifted(23) => 
                           negative_inputs_17_23_port, A_neg_shifted(22) => 
                           negative_inputs_17_22_port, A_neg_shifted(21) => 
                           negative_inputs_17_21_port, A_neg_shifted(20) => 
                           negative_inputs_17_20_port, A_neg_shifted(19) => 
                           negative_inputs_17_19_port, A_neg_shifted(18) => 
                           negative_inputs_17_18_port, A_neg_shifted(17) => 
                           negative_inputs_17_17_port, A_neg_shifted(16) => 
                           negative_inputs_17_16_port, A_neg_shifted(15) => 
                           negative_inputs_17_15_port, A_neg_shifted(14) => 
                           negative_inputs_17_14_port, A_neg_shifted(13) => 
                           negative_inputs_17_13_port, A_neg_shifted(12) => 
                           negative_inputs_17_12_port, A_neg_shifted(11) => 
                           negative_inputs_17_11_port, A_neg_shifted(10) => 
                           negative_inputs_17_10_port, A_neg_shifted(9) => 
                           negative_inputs_17_9_port, A_neg_shifted(8) => 
                           negative_inputs_17_8_port, A_neg_shifted(7) => 
                           negative_inputs_17_7_port, A_neg_shifted(6) => 
                           negative_inputs_17_6_port, A_neg_shifted(5) => 
                           negative_inputs_17_5_port, A_neg_shifted(4) => 
                           negative_inputs_17_4_port, A_neg_shifted(3) => 
                           negative_inputs_17_3_port, A_neg_shifted(2) => 
                           negative_inputs_17_2_port, A_neg_shifted(1) => 
                           negative_inputs_17_1_port, A_neg_shifted(0) => n8, 
                           Sel(2) => sel_8_2_port, Sel(1) => sel_8_1_port, 
                           Sel(0) => sel_8_0_port, Y(63) => 
                           MuxOutputs_8_63_port, Y(62) => MuxOutputs_8_62_port,
                           Y(61) => MuxOutputs_8_61_port, Y(60) => 
                           MuxOutputs_8_60_port, Y(59) => MuxOutputs_8_59_port,
                           Y(58) => MuxOutputs_8_58_port, Y(57) => 
                           MuxOutputs_8_57_port, Y(56) => MuxOutputs_8_56_port,
                           Y(55) => MuxOutputs_8_55_port, Y(54) => 
                           MuxOutputs_8_54_port, Y(53) => MuxOutputs_8_53_port,
                           Y(52) => MuxOutputs_8_52_port, Y(51) => 
                           MuxOutputs_8_51_port, Y(50) => MuxOutputs_8_50_port,
                           Y(49) => MuxOutputs_8_49_port, Y(48) => 
                           MuxOutputs_8_48_port, Y(47) => MuxOutputs_8_47_port,
                           Y(46) => MuxOutputs_8_46_port, Y(45) => 
                           MuxOutputs_8_45_port, Y(44) => MuxOutputs_8_44_port,
                           Y(43) => MuxOutputs_8_43_port, Y(42) => 
                           MuxOutputs_8_42_port, Y(41) => MuxOutputs_8_41_port,
                           Y(40) => MuxOutputs_8_40_port, Y(39) => 
                           MuxOutputs_8_39_port, Y(38) => MuxOutputs_8_38_port,
                           Y(37) => MuxOutputs_8_37_port, Y(36) => 
                           MuxOutputs_8_36_port, Y(35) => MuxOutputs_8_35_port,
                           Y(34) => MuxOutputs_8_34_port, Y(33) => 
                           MuxOutputs_8_33_port, Y(32) => MuxOutputs_8_32_port,
                           Y(31) => MuxOutputs_8_31_port, Y(30) => 
                           MuxOutputs_8_30_port, Y(29) => MuxOutputs_8_29_port,
                           Y(28) => MuxOutputs_8_28_port, Y(27) => 
                           MuxOutputs_8_27_port, Y(26) => MuxOutputs_8_26_port,
                           Y(25) => MuxOutputs_8_25_port, Y(24) => 
                           MuxOutputs_8_24_port, Y(23) => MuxOutputs_8_23_port,
                           Y(22) => MuxOutputs_8_22_port, Y(21) => 
                           MuxOutputs_8_21_port, Y(20) => MuxOutputs_8_20_port,
                           Y(19) => MuxOutputs_8_19_port, Y(18) => 
                           MuxOutputs_8_18_port, Y(17) => MuxOutputs_8_17_port,
                           Y(16) => MuxOutputs_8_16_port, Y(15) => 
                           MuxOutputs_8_15_port, Y(14) => MuxOutputs_8_14_port,
                           Y(13) => MuxOutputs_8_13_port, Y(12) => 
                           MuxOutputs_8_12_port, Y(11) => MuxOutputs_8_11_port,
                           Y(10) => MuxOutputs_8_10_port, Y(9) => 
                           MuxOutputs_8_9_port, Y(8) => MuxOutputs_8_8_port, 
                           Y(7) => MuxOutputs_8_7_port, Y(6) => 
                           MuxOutputs_8_6_port, Y(5) => MuxOutputs_8_5_port, 
                           Y(4) => MuxOutputs_8_4_port, Y(3) => 
                           MuxOutputs_8_3_port, Y(2) => MuxOutputs_8_2_port, 
                           Y(1) => MuxOutputs_8_1_port, Y(0) => 
                           MuxOutputs_8_0_port);
   encoderI_9 : encoder_23 port map( pieceofB(2) => B(19), pieceofB(1) => B(18)
                           , pieceofB(0) => B(17), sel(2) => sel_9_2_port, 
                           sel(1) => sel_9_1_port, sel(0) => sel_9_0_port);
   MUXI_9 : MUX51_MuxNbit64_23 port map( zeroSignal(63) => X_Logic0_port, 
                           zeroSignal(62) => X_Logic0_port, zeroSignal(61) => 
                           X_Logic0_port, zeroSignal(60) => X_Logic0_port, 
                           zeroSignal(59) => X_Logic0_port, zeroSignal(58) => 
                           X_Logic0_port, zeroSignal(57) => X_Logic0_port, 
                           zeroSignal(56) => X_Logic0_port, zeroSignal(55) => 
                           X_Logic0_port, zeroSignal(54) => X_Logic0_port, 
                           zeroSignal(53) => X_Logic0_port, zeroSignal(52) => 
                           X_Logic0_port, zeroSignal(51) => X_Logic0_port, 
                           zeroSignal(50) => X_Logic0_port, zeroSignal(49) => 
                           X_Logic0_port, zeroSignal(48) => X_Logic0_port, 
                           zeroSignal(47) => X_Logic0_port, zeroSignal(46) => 
                           X_Logic0_port, zeroSignal(45) => X_Logic0_port, 
                           zeroSignal(44) => X_Logic0_port, zeroSignal(43) => 
                           X_Logic0_port, zeroSignal(42) => X_Logic0_port, 
                           zeroSignal(41) => X_Logic0_port, zeroSignal(40) => 
                           X_Logic0_port, zeroSignal(39) => X_Logic0_port, 
                           zeroSignal(38) => X_Logic0_port, zeroSignal(37) => 
                           X_Logic0_port, zeroSignal(36) => X_Logic0_port, 
                           zeroSignal(35) => X_Logic0_port, zeroSignal(34) => 
                           X_Logic0_port, zeroSignal(33) => X_Logic0_port, 
                           zeroSignal(32) => X_Logic0_port, zeroSignal(31) => 
                           X_Logic0_port, zeroSignal(30) => X_Logic0_port, 
                           zeroSignal(29) => X_Logic0_port, zeroSignal(28) => 
                           X_Logic0_port, zeroSignal(27) => X_Logic0_port, 
                           zeroSignal(26) => X_Logic0_port, zeroSignal(25) => 
                           X_Logic0_port, zeroSignal(24) => X_Logic0_port, 
                           zeroSignal(23) => X_Logic0_port, zeroSignal(22) => 
                           X_Logic0_port, zeroSignal(21) => X_Logic0_port, 
                           zeroSignal(20) => X_Logic0_port, zeroSignal(19) => 
                           X_Logic0_port, zeroSignal(18) => X_Logic0_port, 
                           zeroSignal(17) => X_Logic0_port, zeroSignal(16) => 
                           X_Logic0_port, zeroSignal(15) => X_Logic0_port, 
                           zeroSignal(14) => X_Logic0_port, zeroSignal(13) => 
                           X_Logic0_port, zeroSignal(12) => X_Logic0_port, 
                           zeroSignal(11) => X_Logic0_port, zeroSignal(10) => 
                           X_Logic0_port, zeroSignal(9) => X_Logic0_port, 
                           zeroSignal(8) => X_Logic0_port, zeroSignal(7) => 
                           X_Logic0_port, zeroSignal(6) => X_Logic0_port, 
                           zeroSignal(5) => X_Logic0_port, zeroSignal(4) => 
                           X_Logic0_port, zeroSignal(3) => X_Logic0_port, 
                           zeroSignal(2) => X_Logic0_port, zeroSignal(1) => 
                           X_Logic0_port, zeroSignal(0) => X_Logic0_port, 
                           A_signal(63) => positive_inputs_18_63_port, 
                           A_signal(62) => positive_inputs_18_62_port, 
                           A_signal(61) => positive_inputs_18_61_port, 
                           A_signal(60) => positive_inputs_18_60_port, 
                           A_signal(59) => positive_inputs_18_59_port, 
                           A_signal(58) => positive_inputs_18_58_port, 
                           A_signal(57) => positive_inputs_18_57_port, 
                           A_signal(56) => positive_inputs_18_56_port, 
                           A_signal(55) => positive_inputs_18_55_port, 
                           A_signal(54) => positive_inputs_18_54_port, 
                           A_signal(53) => positive_inputs_18_53_port, 
                           A_signal(52) => positive_inputs_18_52_port, 
                           A_signal(51) => positive_inputs_18_51_port, 
                           A_signal(50) => positive_inputs_18_50_port, 
                           A_signal(49) => positive_inputs_18_49_port, 
                           A_signal(48) => positive_inputs_18_48_port, 
                           A_signal(47) => positive_inputs_18_47_port, 
                           A_signal(46) => positive_inputs_18_46_port, 
                           A_signal(45) => positive_inputs_18_45_port, 
                           A_signal(44) => positive_inputs_18_44_port, 
                           A_signal(43) => positive_inputs_18_43_port, 
                           A_signal(42) => positive_inputs_18_42_port, 
                           A_signal(41) => positive_inputs_18_41_port, 
                           A_signal(40) => positive_inputs_18_40_port, 
                           A_signal(39) => positive_inputs_18_39_port, 
                           A_signal(38) => positive_inputs_18_38_port, 
                           A_signal(37) => positive_inputs_18_37_port, 
                           A_signal(36) => positive_inputs_18_36_port, 
                           A_signal(35) => positive_inputs_18_35_port, 
                           A_signal(34) => positive_inputs_18_34_port, 
                           A_signal(33) => positive_inputs_18_33_port, 
                           A_signal(32) => positive_inputs_18_32_port, 
                           A_signal(31) => positive_inputs_18_31_port, 
                           A_signal(30) => positive_inputs_18_30_port, 
                           A_signal(29) => positive_inputs_18_29_port, 
                           A_signal(28) => positive_inputs_18_28_port, 
                           A_signal(27) => positive_inputs_18_27_port, 
                           A_signal(26) => positive_inputs_18_26_port, 
                           A_signal(25) => positive_inputs_18_25_port, 
                           A_signal(24) => positive_inputs_18_24_port, 
                           A_signal(23) => positive_inputs_18_23_port, 
                           A_signal(22) => positive_inputs_18_22_port, 
                           A_signal(21) => positive_inputs_18_21_port, 
                           A_signal(20) => positive_inputs_18_20_port, 
                           A_signal(19) => positive_inputs_18_19_port, 
                           A_signal(18) => positive_inputs_18_18_port, 
                           A_signal(17) => positive_inputs_18_17_port, 
                           A_signal(16) => positive_inputs_18_16_port, 
                           A_signal(15) => positive_inputs_18_15_port, 
                           A_signal(14) => positive_inputs_18_14_port, 
                           A_signal(13) => positive_inputs_18_13_port, 
                           A_signal(12) => positive_inputs_18_12_port, 
                           A_signal(11) => positive_inputs_18_11_port, 
                           A_signal(10) => positive_inputs_18_10_port, 
                           A_signal(9) => positive_inputs_18_9_port, 
                           A_signal(8) => positive_inputs_18_8_port, 
                           A_signal(7) => positive_inputs_18_7_port, 
                           A_signal(6) => positive_inputs_18_6_port, 
                           A_signal(5) => positive_inputs_18_5_port, 
                           A_signal(4) => positive_inputs_18_4_port, 
                           A_signal(3) => positive_inputs_18_3_port, 
                           A_signal(2) => positive_inputs_18_2_port, 
                           A_signal(1) => positive_inputs_18_1_port, 
                           A_signal(0) => n8, A_neg(63) => 
                           negative_inputs_18_63_port, A_neg(62) => 
                           negative_inputs_18_62_port, A_neg(61) => 
                           negative_inputs_18_61_port, A_neg(60) => 
                           negative_inputs_18_60_port, A_neg(59) => 
                           negative_inputs_18_59_port, A_neg(58) => 
                           negative_inputs_18_58_port, A_neg(57) => 
                           negative_inputs_18_57_port, A_neg(56) => 
                           negative_inputs_18_56_port, A_neg(55) => 
                           negative_inputs_18_55_port, A_neg(54) => 
                           negative_inputs_18_54_port, A_neg(53) => 
                           negative_inputs_18_53_port, A_neg(52) => 
                           negative_inputs_18_52_port, A_neg(51) => 
                           negative_inputs_18_51_port, A_neg(50) => 
                           negative_inputs_18_50_port, A_neg(49) => 
                           negative_inputs_18_49_port, A_neg(48) => 
                           negative_inputs_18_48_port, A_neg(47) => 
                           negative_inputs_18_47_port, A_neg(46) => 
                           negative_inputs_18_46_port, A_neg(45) => 
                           negative_inputs_18_45_port, A_neg(44) => 
                           negative_inputs_18_44_port, A_neg(43) => 
                           negative_inputs_18_43_port, A_neg(42) => 
                           negative_inputs_18_42_port, A_neg(41) => 
                           negative_inputs_18_41_port, A_neg(40) => 
                           negative_inputs_18_40_port, A_neg(39) => 
                           negative_inputs_18_39_port, A_neg(38) => 
                           negative_inputs_18_38_port, A_neg(37) => 
                           negative_inputs_18_37_port, A_neg(36) => 
                           negative_inputs_18_36_port, A_neg(35) => 
                           negative_inputs_18_35_port, A_neg(34) => 
                           negative_inputs_18_34_port, A_neg(33) => 
                           negative_inputs_18_33_port, A_neg(32) => 
                           negative_inputs_18_32_port, A_neg(31) => 
                           negative_inputs_18_31_port, A_neg(30) => 
                           negative_inputs_18_30_port, A_neg(29) => 
                           negative_inputs_18_29_port, A_neg(28) => 
                           negative_inputs_18_28_port, A_neg(27) => 
                           negative_inputs_18_27_port, A_neg(26) => 
                           negative_inputs_18_26_port, A_neg(25) => 
                           negative_inputs_18_25_port, A_neg(24) => 
                           negative_inputs_18_24_port, A_neg(23) => 
                           negative_inputs_18_23_port, A_neg(22) => 
                           negative_inputs_18_22_port, A_neg(21) => 
                           negative_inputs_18_21_port, A_neg(20) => 
                           negative_inputs_18_20_port, A_neg(19) => 
                           negative_inputs_18_19_port, A_neg(18) => 
                           negative_inputs_18_18_port, A_neg(17) => 
                           negative_inputs_18_17_port, A_neg(16) => 
                           negative_inputs_18_16_port, A_neg(15) => 
                           negative_inputs_18_15_port, A_neg(14) => 
                           negative_inputs_18_14_port, A_neg(13) => 
                           negative_inputs_18_13_port, A_neg(12) => 
                           negative_inputs_18_12_port, A_neg(11) => 
                           negative_inputs_18_11_port, A_neg(10) => 
                           negative_inputs_18_10_port, A_neg(9) => 
                           negative_inputs_18_9_port, A_neg(8) => 
                           negative_inputs_18_8_port, A_neg(7) => 
                           negative_inputs_18_7_port, A_neg(6) => 
                           negative_inputs_18_6_port, A_neg(5) => 
                           negative_inputs_18_5_port, A_neg(4) => 
                           negative_inputs_18_4_port, A_neg(3) => 
                           negative_inputs_18_3_port, A_neg(2) => 
                           negative_inputs_18_2_port, A_neg(1) => 
                           negative_inputs_18_1_port, A_neg(0) => n8, 
                           A_shifted(63) => positive_inputs_19_63_port, 
                           A_shifted(62) => positive_inputs_19_62_port, 
                           A_shifted(61) => positive_inputs_19_61_port, 
                           A_shifted(60) => positive_inputs_19_60_port, 
                           A_shifted(59) => positive_inputs_19_59_port, 
                           A_shifted(58) => positive_inputs_19_58_port, 
                           A_shifted(57) => positive_inputs_19_57_port, 
                           A_shifted(56) => positive_inputs_19_56_port, 
                           A_shifted(55) => positive_inputs_19_55_port, 
                           A_shifted(54) => positive_inputs_19_54_port, 
                           A_shifted(53) => positive_inputs_19_53_port, 
                           A_shifted(52) => positive_inputs_19_52_port, 
                           A_shifted(51) => positive_inputs_19_51_port, 
                           A_shifted(50) => positive_inputs_19_50_port, 
                           A_shifted(49) => positive_inputs_19_49_port, 
                           A_shifted(48) => positive_inputs_19_48_port, 
                           A_shifted(47) => positive_inputs_19_47_port, 
                           A_shifted(46) => positive_inputs_19_46_port, 
                           A_shifted(45) => positive_inputs_19_45_port, 
                           A_shifted(44) => positive_inputs_19_44_port, 
                           A_shifted(43) => positive_inputs_19_43_port, 
                           A_shifted(42) => positive_inputs_19_42_port, 
                           A_shifted(41) => positive_inputs_19_41_port, 
                           A_shifted(40) => positive_inputs_19_40_port, 
                           A_shifted(39) => positive_inputs_19_39_port, 
                           A_shifted(38) => positive_inputs_19_38_port, 
                           A_shifted(37) => positive_inputs_19_37_port, 
                           A_shifted(36) => positive_inputs_19_36_port, 
                           A_shifted(35) => positive_inputs_19_35_port, 
                           A_shifted(34) => positive_inputs_19_34_port, 
                           A_shifted(33) => positive_inputs_19_33_port, 
                           A_shifted(32) => positive_inputs_19_32_port, 
                           A_shifted(31) => positive_inputs_19_31_port, 
                           A_shifted(30) => positive_inputs_19_30_port, 
                           A_shifted(29) => positive_inputs_19_29_port, 
                           A_shifted(28) => positive_inputs_19_28_port, 
                           A_shifted(27) => positive_inputs_19_27_port, 
                           A_shifted(26) => positive_inputs_19_26_port, 
                           A_shifted(25) => positive_inputs_19_25_port, 
                           A_shifted(24) => positive_inputs_19_24_port, 
                           A_shifted(23) => positive_inputs_19_23_port, 
                           A_shifted(22) => positive_inputs_19_22_port, 
                           A_shifted(21) => positive_inputs_19_21_port, 
                           A_shifted(20) => positive_inputs_19_20_port, 
                           A_shifted(19) => positive_inputs_19_19_port, 
                           A_shifted(18) => positive_inputs_19_18_port, 
                           A_shifted(17) => positive_inputs_19_17_port, 
                           A_shifted(16) => positive_inputs_19_16_port, 
                           A_shifted(15) => positive_inputs_19_15_port, 
                           A_shifted(14) => positive_inputs_19_14_port, 
                           A_shifted(13) => positive_inputs_19_13_port, 
                           A_shifted(12) => positive_inputs_19_12_port, 
                           A_shifted(11) => positive_inputs_19_11_port, 
                           A_shifted(10) => positive_inputs_19_10_port, 
                           A_shifted(9) => positive_inputs_19_9_port, 
                           A_shifted(8) => positive_inputs_19_8_port, 
                           A_shifted(7) => positive_inputs_19_7_port, 
                           A_shifted(6) => positive_inputs_19_6_port, 
                           A_shifted(5) => positive_inputs_19_5_port, 
                           A_shifted(4) => positive_inputs_19_4_port, 
                           A_shifted(3) => positive_inputs_19_3_port, 
                           A_shifted(2) => positive_inputs_19_2_port, 
                           A_shifted(1) => positive_inputs_19_1_port, 
                           A_shifted(0) => n8, A_neg_shifted(63) => 
                           negative_inputs_19_63_port, A_neg_shifted(62) => 
                           negative_inputs_19_62_port, A_neg_shifted(61) => 
                           negative_inputs_19_61_port, A_neg_shifted(60) => 
                           negative_inputs_19_60_port, A_neg_shifted(59) => 
                           negative_inputs_19_59_port, A_neg_shifted(58) => 
                           negative_inputs_19_58_port, A_neg_shifted(57) => 
                           negative_inputs_19_57_port, A_neg_shifted(56) => 
                           negative_inputs_19_56_port, A_neg_shifted(55) => 
                           negative_inputs_19_55_port, A_neg_shifted(54) => 
                           negative_inputs_19_54_port, A_neg_shifted(53) => 
                           negative_inputs_19_53_port, A_neg_shifted(52) => 
                           negative_inputs_19_52_port, A_neg_shifted(51) => 
                           negative_inputs_19_51_port, A_neg_shifted(50) => 
                           negative_inputs_19_50_port, A_neg_shifted(49) => 
                           negative_inputs_19_49_port, A_neg_shifted(48) => 
                           negative_inputs_19_48_port, A_neg_shifted(47) => 
                           negative_inputs_19_47_port, A_neg_shifted(46) => 
                           negative_inputs_19_46_port, A_neg_shifted(45) => 
                           negative_inputs_19_45_port, A_neg_shifted(44) => 
                           negative_inputs_19_44_port, A_neg_shifted(43) => 
                           negative_inputs_19_43_port, A_neg_shifted(42) => 
                           negative_inputs_19_42_port, A_neg_shifted(41) => 
                           negative_inputs_19_41_port, A_neg_shifted(40) => 
                           negative_inputs_19_40_port, A_neg_shifted(39) => 
                           negative_inputs_19_39_port, A_neg_shifted(38) => 
                           negative_inputs_19_38_port, A_neg_shifted(37) => 
                           negative_inputs_19_37_port, A_neg_shifted(36) => 
                           negative_inputs_19_36_port, A_neg_shifted(35) => 
                           negative_inputs_19_35_port, A_neg_shifted(34) => 
                           negative_inputs_19_34_port, A_neg_shifted(33) => 
                           negative_inputs_19_33_port, A_neg_shifted(32) => 
                           negative_inputs_19_32_port, A_neg_shifted(31) => 
                           negative_inputs_19_31_port, A_neg_shifted(30) => 
                           negative_inputs_19_30_port, A_neg_shifted(29) => 
                           negative_inputs_19_29_port, A_neg_shifted(28) => 
                           negative_inputs_19_28_port, A_neg_shifted(27) => 
                           negative_inputs_19_27_port, A_neg_shifted(26) => 
                           negative_inputs_19_26_port, A_neg_shifted(25) => 
                           negative_inputs_19_25_port, A_neg_shifted(24) => 
                           negative_inputs_19_24_port, A_neg_shifted(23) => 
                           negative_inputs_19_23_port, A_neg_shifted(22) => 
                           negative_inputs_19_22_port, A_neg_shifted(21) => 
                           negative_inputs_19_21_port, A_neg_shifted(20) => 
                           negative_inputs_19_20_port, A_neg_shifted(19) => 
                           negative_inputs_19_19_port, A_neg_shifted(18) => 
                           negative_inputs_19_18_port, A_neg_shifted(17) => 
                           negative_inputs_19_17_port, A_neg_shifted(16) => 
                           negative_inputs_19_16_port, A_neg_shifted(15) => 
                           negative_inputs_19_15_port, A_neg_shifted(14) => 
                           negative_inputs_19_14_port, A_neg_shifted(13) => 
                           negative_inputs_19_13_port, A_neg_shifted(12) => 
                           negative_inputs_19_12_port, A_neg_shifted(11) => 
                           negative_inputs_19_11_port, A_neg_shifted(10) => 
                           negative_inputs_19_10_port, A_neg_shifted(9) => 
                           negative_inputs_19_9_port, A_neg_shifted(8) => 
                           negative_inputs_19_8_port, A_neg_shifted(7) => 
                           negative_inputs_19_7_port, A_neg_shifted(6) => 
                           negative_inputs_19_6_port, A_neg_shifted(5) => 
                           negative_inputs_19_5_port, A_neg_shifted(4) => 
                           negative_inputs_19_4_port, A_neg_shifted(3) => 
                           negative_inputs_19_3_port, A_neg_shifted(2) => 
                           negative_inputs_19_2_port, A_neg_shifted(1) => 
                           negative_inputs_19_1_port, A_neg_shifted(0) => n8, 
                           Sel(2) => sel_9_2_port, Sel(1) => sel_9_1_port, 
                           Sel(0) => sel_9_0_port, Y(63) => 
                           MuxOutputs_9_63_port, Y(62) => MuxOutputs_9_62_port,
                           Y(61) => MuxOutputs_9_61_port, Y(60) => 
                           MuxOutputs_9_60_port, Y(59) => MuxOutputs_9_59_port,
                           Y(58) => MuxOutputs_9_58_port, Y(57) => 
                           MuxOutputs_9_57_port, Y(56) => MuxOutputs_9_56_port,
                           Y(55) => MuxOutputs_9_55_port, Y(54) => 
                           MuxOutputs_9_54_port, Y(53) => MuxOutputs_9_53_port,
                           Y(52) => MuxOutputs_9_52_port, Y(51) => 
                           MuxOutputs_9_51_port, Y(50) => MuxOutputs_9_50_port,
                           Y(49) => MuxOutputs_9_49_port, Y(48) => 
                           MuxOutputs_9_48_port, Y(47) => MuxOutputs_9_47_port,
                           Y(46) => MuxOutputs_9_46_port, Y(45) => 
                           MuxOutputs_9_45_port, Y(44) => MuxOutputs_9_44_port,
                           Y(43) => MuxOutputs_9_43_port, Y(42) => 
                           MuxOutputs_9_42_port, Y(41) => MuxOutputs_9_41_port,
                           Y(40) => MuxOutputs_9_40_port, Y(39) => 
                           MuxOutputs_9_39_port, Y(38) => MuxOutputs_9_38_port,
                           Y(37) => MuxOutputs_9_37_port, Y(36) => 
                           MuxOutputs_9_36_port, Y(35) => MuxOutputs_9_35_port,
                           Y(34) => MuxOutputs_9_34_port, Y(33) => 
                           MuxOutputs_9_33_port, Y(32) => MuxOutputs_9_32_port,
                           Y(31) => MuxOutputs_9_31_port, Y(30) => 
                           MuxOutputs_9_30_port, Y(29) => MuxOutputs_9_29_port,
                           Y(28) => MuxOutputs_9_28_port, Y(27) => 
                           MuxOutputs_9_27_port, Y(26) => MuxOutputs_9_26_port,
                           Y(25) => MuxOutputs_9_25_port, Y(24) => 
                           MuxOutputs_9_24_port, Y(23) => MuxOutputs_9_23_port,
                           Y(22) => MuxOutputs_9_22_port, Y(21) => 
                           MuxOutputs_9_21_port, Y(20) => MuxOutputs_9_20_port,
                           Y(19) => MuxOutputs_9_19_port, Y(18) => 
                           MuxOutputs_9_18_port, Y(17) => MuxOutputs_9_17_port,
                           Y(16) => MuxOutputs_9_16_port, Y(15) => 
                           MuxOutputs_9_15_port, Y(14) => MuxOutputs_9_14_port,
                           Y(13) => MuxOutputs_9_13_port, Y(12) => 
                           MuxOutputs_9_12_port, Y(11) => MuxOutputs_9_11_port,
                           Y(10) => MuxOutputs_9_10_port, Y(9) => 
                           MuxOutputs_9_9_port, Y(8) => MuxOutputs_9_8_port, 
                           Y(7) => MuxOutputs_9_7_port, Y(6) => 
                           MuxOutputs_9_6_port, Y(5) => MuxOutputs_9_5_port, 
                           Y(4) => MuxOutputs_9_4_port, Y(3) => 
                           MuxOutputs_9_3_port, Y(2) => MuxOutputs_9_2_port, 
                           Y(1) => MuxOutputs_9_1_port, Y(0) => 
                           MuxOutputs_9_0_port);
   encoderI_10 : encoder_22 port map( pieceofB(2) => B(21), pieceofB(1) => 
                           B(20), pieceofB(0) => B(19), sel(2) => sel_10_2_port
                           , sel(1) => sel_10_1_port, sel(0) => sel_10_0_port);
   MUXI_10 : MUX51_MuxNbit64_22 port map( zeroSignal(63) => X_Logic0_port, 
                           zeroSignal(62) => X_Logic0_port, zeroSignal(61) => 
                           X_Logic0_port, zeroSignal(60) => X_Logic0_port, 
                           zeroSignal(59) => X_Logic0_port, zeroSignal(58) => 
                           X_Logic0_port, zeroSignal(57) => X_Logic0_port, 
                           zeroSignal(56) => X_Logic0_port, zeroSignal(55) => 
                           X_Logic0_port, zeroSignal(54) => X_Logic0_port, 
                           zeroSignal(53) => X_Logic0_port, zeroSignal(52) => 
                           X_Logic0_port, zeroSignal(51) => X_Logic0_port, 
                           zeroSignal(50) => X_Logic0_port, zeroSignal(49) => 
                           X_Logic0_port, zeroSignal(48) => X_Logic0_port, 
                           zeroSignal(47) => X_Logic0_port, zeroSignal(46) => 
                           X_Logic0_port, zeroSignal(45) => X_Logic0_port, 
                           zeroSignal(44) => X_Logic0_port, zeroSignal(43) => 
                           X_Logic0_port, zeroSignal(42) => X_Logic0_port, 
                           zeroSignal(41) => X_Logic0_port, zeroSignal(40) => 
                           X_Logic0_port, zeroSignal(39) => X_Logic0_port, 
                           zeroSignal(38) => X_Logic0_port, zeroSignal(37) => 
                           X_Logic0_port, zeroSignal(36) => X_Logic0_port, 
                           zeroSignal(35) => X_Logic0_port, zeroSignal(34) => 
                           X_Logic0_port, zeroSignal(33) => X_Logic0_port, 
                           zeroSignal(32) => X_Logic0_port, zeroSignal(31) => 
                           X_Logic0_port, zeroSignal(30) => X_Logic0_port, 
                           zeroSignal(29) => X_Logic0_port, zeroSignal(28) => 
                           X_Logic0_port, zeroSignal(27) => X_Logic0_port, 
                           zeroSignal(26) => X_Logic0_port, zeroSignal(25) => 
                           X_Logic0_port, zeroSignal(24) => X_Logic0_port, 
                           zeroSignal(23) => X_Logic0_port, zeroSignal(22) => 
                           X_Logic0_port, zeroSignal(21) => X_Logic0_port, 
                           zeroSignal(20) => X_Logic0_port, zeroSignal(19) => 
                           X_Logic0_port, zeroSignal(18) => X_Logic0_port, 
                           zeroSignal(17) => X_Logic0_port, zeroSignal(16) => 
                           X_Logic0_port, zeroSignal(15) => X_Logic0_port, 
                           zeroSignal(14) => X_Logic0_port, zeroSignal(13) => 
                           X_Logic0_port, zeroSignal(12) => X_Logic0_port, 
                           zeroSignal(11) => X_Logic0_port, zeroSignal(10) => 
                           X_Logic0_port, zeroSignal(9) => X_Logic0_port, 
                           zeroSignal(8) => X_Logic0_port, zeroSignal(7) => 
                           X_Logic0_port, zeroSignal(6) => X_Logic0_port, 
                           zeroSignal(5) => X_Logic0_port, zeroSignal(4) => 
                           X_Logic0_port, zeroSignal(3) => X_Logic0_port, 
                           zeroSignal(2) => X_Logic0_port, zeroSignal(1) => 
                           X_Logic0_port, zeroSignal(0) => X_Logic0_port, 
                           A_signal(63) => positive_inputs_20_63_port, 
                           A_signal(62) => positive_inputs_20_62_port, 
                           A_signal(61) => positive_inputs_20_61_port, 
                           A_signal(60) => positive_inputs_20_60_port, 
                           A_signal(59) => positive_inputs_20_59_port, 
                           A_signal(58) => positive_inputs_20_58_port, 
                           A_signal(57) => positive_inputs_20_57_port, 
                           A_signal(56) => positive_inputs_20_56_port, 
                           A_signal(55) => positive_inputs_20_55_port, 
                           A_signal(54) => positive_inputs_20_54_port, 
                           A_signal(53) => positive_inputs_20_53_port, 
                           A_signal(52) => positive_inputs_20_52_port, 
                           A_signal(51) => positive_inputs_20_51_port, 
                           A_signal(50) => positive_inputs_20_50_port, 
                           A_signal(49) => positive_inputs_20_49_port, 
                           A_signal(48) => positive_inputs_20_48_port, 
                           A_signal(47) => positive_inputs_20_47_port, 
                           A_signal(46) => positive_inputs_20_46_port, 
                           A_signal(45) => positive_inputs_20_45_port, 
                           A_signal(44) => positive_inputs_20_44_port, 
                           A_signal(43) => positive_inputs_20_43_port, 
                           A_signal(42) => positive_inputs_20_42_port, 
                           A_signal(41) => positive_inputs_20_41_port, 
                           A_signal(40) => positive_inputs_20_40_port, 
                           A_signal(39) => positive_inputs_20_39_port, 
                           A_signal(38) => positive_inputs_20_38_port, 
                           A_signal(37) => positive_inputs_20_37_port, 
                           A_signal(36) => positive_inputs_20_36_port, 
                           A_signal(35) => positive_inputs_20_35_port, 
                           A_signal(34) => positive_inputs_20_34_port, 
                           A_signal(33) => positive_inputs_20_33_port, 
                           A_signal(32) => positive_inputs_20_32_port, 
                           A_signal(31) => positive_inputs_20_31_port, 
                           A_signal(30) => positive_inputs_20_30_port, 
                           A_signal(29) => positive_inputs_20_29_port, 
                           A_signal(28) => positive_inputs_20_28_port, 
                           A_signal(27) => positive_inputs_20_27_port, 
                           A_signal(26) => positive_inputs_20_26_port, 
                           A_signal(25) => positive_inputs_20_25_port, 
                           A_signal(24) => positive_inputs_20_24_port, 
                           A_signal(23) => positive_inputs_20_23_port, 
                           A_signal(22) => positive_inputs_20_22_port, 
                           A_signal(21) => positive_inputs_20_21_port, 
                           A_signal(20) => positive_inputs_20_20_port, 
                           A_signal(19) => positive_inputs_20_19_port, 
                           A_signal(18) => positive_inputs_20_18_port, 
                           A_signal(17) => positive_inputs_20_17_port, 
                           A_signal(16) => positive_inputs_20_16_port, 
                           A_signal(15) => positive_inputs_20_15_port, 
                           A_signal(14) => positive_inputs_20_14_port, 
                           A_signal(13) => positive_inputs_20_13_port, 
                           A_signal(12) => positive_inputs_20_12_port, 
                           A_signal(11) => positive_inputs_20_11_port, 
                           A_signal(10) => positive_inputs_20_10_port, 
                           A_signal(9) => positive_inputs_20_9_port, 
                           A_signal(8) => positive_inputs_20_8_port, 
                           A_signal(7) => positive_inputs_20_7_port, 
                           A_signal(6) => positive_inputs_20_6_port, 
                           A_signal(5) => positive_inputs_20_5_port, 
                           A_signal(4) => positive_inputs_20_4_port, 
                           A_signal(3) => positive_inputs_20_3_port, 
                           A_signal(2) => positive_inputs_20_2_port, 
                           A_signal(1) => positive_inputs_20_1_port, 
                           A_signal(0) => n8, A_neg(63) => 
                           negative_inputs_20_63_port, A_neg(62) => 
                           negative_inputs_20_62_port, A_neg(61) => 
                           negative_inputs_20_61_port, A_neg(60) => 
                           negative_inputs_20_60_port, A_neg(59) => 
                           negative_inputs_20_59_port, A_neg(58) => 
                           negative_inputs_20_58_port, A_neg(57) => 
                           negative_inputs_20_57_port, A_neg(56) => 
                           negative_inputs_20_56_port, A_neg(55) => 
                           negative_inputs_20_55_port, A_neg(54) => 
                           negative_inputs_20_54_port, A_neg(53) => 
                           negative_inputs_20_53_port, A_neg(52) => 
                           negative_inputs_20_52_port, A_neg(51) => 
                           negative_inputs_20_51_port, A_neg(50) => 
                           negative_inputs_20_50_port, A_neg(49) => 
                           negative_inputs_20_49_port, A_neg(48) => 
                           negative_inputs_20_48_port, A_neg(47) => 
                           negative_inputs_20_47_port, A_neg(46) => 
                           negative_inputs_20_46_port, A_neg(45) => 
                           negative_inputs_20_45_port, A_neg(44) => 
                           negative_inputs_20_44_port, A_neg(43) => 
                           negative_inputs_20_43_port, A_neg(42) => 
                           negative_inputs_20_42_port, A_neg(41) => 
                           negative_inputs_20_41_port, A_neg(40) => 
                           negative_inputs_20_40_port, A_neg(39) => 
                           negative_inputs_20_39_port, A_neg(38) => 
                           negative_inputs_20_38_port, A_neg(37) => 
                           negative_inputs_20_37_port, A_neg(36) => 
                           negative_inputs_20_36_port, A_neg(35) => 
                           negative_inputs_20_35_port, A_neg(34) => 
                           negative_inputs_20_34_port, A_neg(33) => 
                           negative_inputs_20_33_port, A_neg(32) => 
                           negative_inputs_20_32_port, A_neg(31) => 
                           negative_inputs_20_31_port, A_neg(30) => 
                           negative_inputs_20_30_port, A_neg(29) => 
                           negative_inputs_20_29_port, A_neg(28) => 
                           negative_inputs_20_28_port, A_neg(27) => 
                           negative_inputs_20_27_port, A_neg(26) => 
                           negative_inputs_20_26_port, A_neg(25) => 
                           negative_inputs_20_25_port, A_neg(24) => 
                           negative_inputs_20_24_port, A_neg(23) => 
                           negative_inputs_20_23_port, A_neg(22) => 
                           negative_inputs_20_22_port, A_neg(21) => 
                           negative_inputs_20_21_port, A_neg(20) => 
                           negative_inputs_20_20_port, A_neg(19) => 
                           negative_inputs_20_19_port, A_neg(18) => 
                           negative_inputs_20_18_port, A_neg(17) => 
                           negative_inputs_20_17_port, A_neg(16) => 
                           negative_inputs_20_16_port, A_neg(15) => 
                           negative_inputs_20_15_port, A_neg(14) => 
                           negative_inputs_20_14_port, A_neg(13) => 
                           negative_inputs_20_13_port, A_neg(12) => 
                           negative_inputs_20_12_port, A_neg(11) => 
                           negative_inputs_20_11_port, A_neg(10) => 
                           negative_inputs_20_10_port, A_neg(9) => 
                           negative_inputs_20_9_port, A_neg(8) => 
                           negative_inputs_20_8_port, A_neg(7) => 
                           negative_inputs_20_7_port, A_neg(6) => 
                           negative_inputs_20_6_port, A_neg(5) => 
                           negative_inputs_20_5_port, A_neg(4) => 
                           negative_inputs_20_4_port, A_neg(3) => 
                           negative_inputs_20_3_port, A_neg(2) => 
                           negative_inputs_20_2_port, A_neg(1) => 
                           negative_inputs_20_1_port, A_neg(0) => n8, 
                           A_shifted(63) => positive_inputs_21_63_port, 
                           A_shifted(62) => positive_inputs_21_62_port, 
                           A_shifted(61) => positive_inputs_21_61_port, 
                           A_shifted(60) => positive_inputs_21_60_port, 
                           A_shifted(59) => positive_inputs_21_59_port, 
                           A_shifted(58) => positive_inputs_21_58_port, 
                           A_shifted(57) => positive_inputs_21_57_port, 
                           A_shifted(56) => positive_inputs_21_56_port, 
                           A_shifted(55) => positive_inputs_21_55_port, 
                           A_shifted(54) => positive_inputs_21_54_port, 
                           A_shifted(53) => positive_inputs_21_53_port, 
                           A_shifted(52) => positive_inputs_21_52_port, 
                           A_shifted(51) => positive_inputs_21_51_port, 
                           A_shifted(50) => positive_inputs_21_50_port, 
                           A_shifted(49) => positive_inputs_21_49_port, 
                           A_shifted(48) => positive_inputs_21_48_port, 
                           A_shifted(47) => positive_inputs_21_47_port, 
                           A_shifted(46) => positive_inputs_21_46_port, 
                           A_shifted(45) => positive_inputs_21_45_port, 
                           A_shifted(44) => positive_inputs_21_44_port, 
                           A_shifted(43) => positive_inputs_21_43_port, 
                           A_shifted(42) => positive_inputs_21_42_port, 
                           A_shifted(41) => positive_inputs_21_41_port, 
                           A_shifted(40) => positive_inputs_21_40_port, 
                           A_shifted(39) => positive_inputs_21_39_port, 
                           A_shifted(38) => positive_inputs_21_38_port, 
                           A_shifted(37) => positive_inputs_21_37_port, 
                           A_shifted(36) => positive_inputs_21_36_port, 
                           A_shifted(35) => positive_inputs_21_35_port, 
                           A_shifted(34) => positive_inputs_21_34_port, 
                           A_shifted(33) => positive_inputs_21_33_port, 
                           A_shifted(32) => positive_inputs_21_32_port, 
                           A_shifted(31) => positive_inputs_21_31_port, 
                           A_shifted(30) => positive_inputs_21_30_port, 
                           A_shifted(29) => positive_inputs_21_29_port, 
                           A_shifted(28) => positive_inputs_21_28_port, 
                           A_shifted(27) => positive_inputs_21_27_port, 
                           A_shifted(26) => positive_inputs_21_26_port, 
                           A_shifted(25) => positive_inputs_21_25_port, 
                           A_shifted(24) => positive_inputs_21_24_port, 
                           A_shifted(23) => positive_inputs_21_23_port, 
                           A_shifted(22) => positive_inputs_21_22_port, 
                           A_shifted(21) => positive_inputs_21_21_port, 
                           A_shifted(20) => positive_inputs_21_20_port, 
                           A_shifted(19) => positive_inputs_21_19_port, 
                           A_shifted(18) => positive_inputs_21_18_port, 
                           A_shifted(17) => positive_inputs_21_17_port, 
                           A_shifted(16) => positive_inputs_21_16_port, 
                           A_shifted(15) => positive_inputs_21_15_port, 
                           A_shifted(14) => positive_inputs_21_14_port, 
                           A_shifted(13) => positive_inputs_21_13_port, 
                           A_shifted(12) => positive_inputs_21_12_port, 
                           A_shifted(11) => positive_inputs_21_11_port, 
                           A_shifted(10) => positive_inputs_21_10_port, 
                           A_shifted(9) => positive_inputs_21_9_port, 
                           A_shifted(8) => positive_inputs_21_8_port, 
                           A_shifted(7) => positive_inputs_21_7_port, 
                           A_shifted(6) => positive_inputs_21_6_port, 
                           A_shifted(5) => positive_inputs_21_5_port, 
                           A_shifted(4) => positive_inputs_21_4_port, 
                           A_shifted(3) => positive_inputs_21_3_port, 
                           A_shifted(2) => positive_inputs_21_2_port, 
                           A_shifted(1) => positive_inputs_21_1_port, 
                           A_shifted(0) => n8, A_neg_shifted(63) => 
                           negative_inputs_21_63_port, A_neg_shifted(62) => 
                           negative_inputs_21_62_port, A_neg_shifted(61) => 
                           negative_inputs_21_61_port, A_neg_shifted(60) => 
                           negative_inputs_21_60_port, A_neg_shifted(59) => 
                           negative_inputs_21_59_port, A_neg_shifted(58) => 
                           negative_inputs_21_58_port, A_neg_shifted(57) => 
                           negative_inputs_21_57_port, A_neg_shifted(56) => 
                           negative_inputs_21_56_port, A_neg_shifted(55) => 
                           negative_inputs_21_55_port, A_neg_shifted(54) => 
                           negative_inputs_21_54_port, A_neg_shifted(53) => 
                           negative_inputs_21_53_port, A_neg_shifted(52) => 
                           negative_inputs_21_52_port, A_neg_shifted(51) => 
                           negative_inputs_21_51_port, A_neg_shifted(50) => 
                           negative_inputs_21_50_port, A_neg_shifted(49) => 
                           negative_inputs_21_49_port, A_neg_shifted(48) => 
                           negative_inputs_21_48_port, A_neg_shifted(47) => 
                           negative_inputs_21_47_port, A_neg_shifted(46) => 
                           negative_inputs_21_46_port, A_neg_shifted(45) => 
                           negative_inputs_21_45_port, A_neg_shifted(44) => 
                           negative_inputs_21_44_port, A_neg_shifted(43) => 
                           negative_inputs_21_43_port, A_neg_shifted(42) => 
                           negative_inputs_21_42_port, A_neg_shifted(41) => 
                           negative_inputs_21_41_port, A_neg_shifted(40) => 
                           negative_inputs_21_40_port, A_neg_shifted(39) => 
                           negative_inputs_21_39_port, A_neg_shifted(38) => 
                           negative_inputs_21_38_port, A_neg_shifted(37) => 
                           negative_inputs_21_37_port, A_neg_shifted(36) => 
                           negative_inputs_21_36_port, A_neg_shifted(35) => 
                           negative_inputs_21_35_port, A_neg_shifted(34) => 
                           negative_inputs_21_34_port, A_neg_shifted(33) => 
                           negative_inputs_21_33_port, A_neg_shifted(32) => 
                           negative_inputs_21_32_port, A_neg_shifted(31) => 
                           negative_inputs_21_31_port, A_neg_shifted(30) => 
                           negative_inputs_21_30_port, A_neg_shifted(29) => 
                           negative_inputs_21_29_port, A_neg_shifted(28) => 
                           negative_inputs_21_28_port, A_neg_shifted(27) => 
                           negative_inputs_21_27_port, A_neg_shifted(26) => 
                           negative_inputs_21_26_port, A_neg_shifted(25) => 
                           negative_inputs_21_25_port, A_neg_shifted(24) => 
                           negative_inputs_21_24_port, A_neg_shifted(23) => 
                           negative_inputs_21_23_port, A_neg_shifted(22) => 
                           negative_inputs_21_22_port, A_neg_shifted(21) => 
                           negative_inputs_21_21_port, A_neg_shifted(20) => 
                           negative_inputs_21_20_port, A_neg_shifted(19) => 
                           negative_inputs_21_19_port, A_neg_shifted(18) => 
                           negative_inputs_21_18_port, A_neg_shifted(17) => 
                           negative_inputs_21_17_port, A_neg_shifted(16) => 
                           negative_inputs_21_16_port, A_neg_shifted(15) => 
                           negative_inputs_21_15_port, A_neg_shifted(14) => 
                           negative_inputs_21_14_port, A_neg_shifted(13) => 
                           negative_inputs_21_13_port, A_neg_shifted(12) => 
                           negative_inputs_21_12_port, A_neg_shifted(11) => 
                           negative_inputs_21_11_port, A_neg_shifted(10) => 
                           negative_inputs_21_10_port, A_neg_shifted(9) => 
                           negative_inputs_21_9_port, A_neg_shifted(8) => 
                           negative_inputs_21_8_port, A_neg_shifted(7) => 
                           negative_inputs_21_7_port, A_neg_shifted(6) => 
                           negative_inputs_21_6_port, A_neg_shifted(5) => 
                           negative_inputs_21_5_port, A_neg_shifted(4) => 
                           negative_inputs_21_4_port, A_neg_shifted(3) => 
                           negative_inputs_21_3_port, A_neg_shifted(2) => 
                           negative_inputs_21_2_port, A_neg_shifted(1) => 
                           negative_inputs_21_1_port, A_neg_shifted(0) => n8, 
                           Sel(2) => sel_10_2_port, Sel(1) => sel_10_1_port, 
                           Sel(0) => sel_10_0_port, Y(63) => 
                           MuxOutputs_10_63_port, Y(62) => 
                           MuxOutputs_10_62_port, Y(61) => 
                           MuxOutputs_10_61_port, Y(60) => 
                           MuxOutputs_10_60_port, Y(59) => 
                           MuxOutputs_10_59_port, Y(58) => 
                           MuxOutputs_10_58_port, Y(57) => 
                           MuxOutputs_10_57_port, Y(56) => 
                           MuxOutputs_10_56_port, Y(55) => 
                           MuxOutputs_10_55_port, Y(54) => 
                           MuxOutputs_10_54_port, Y(53) => 
                           MuxOutputs_10_53_port, Y(52) => 
                           MuxOutputs_10_52_port, Y(51) => 
                           MuxOutputs_10_51_port, Y(50) => 
                           MuxOutputs_10_50_port, Y(49) => 
                           MuxOutputs_10_49_port, Y(48) => 
                           MuxOutputs_10_48_port, Y(47) => 
                           MuxOutputs_10_47_port, Y(46) => 
                           MuxOutputs_10_46_port, Y(45) => 
                           MuxOutputs_10_45_port, Y(44) => 
                           MuxOutputs_10_44_port, Y(43) => 
                           MuxOutputs_10_43_port, Y(42) => 
                           MuxOutputs_10_42_port, Y(41) => 
                           MuxOutputs_10_41_port, Y(40) => 
                           MuxOutputs_10_40_port, Y(39) => 
                           MuxOutputs_10_39_port, Y(38) => 
                           MuxOutputs_10_38_port, Y(37) => 
                           MuxOutputs_10_37_port, Y(36) => 
                           MuxOutputs_10_36_port, Y(35) => 
                           MuxOutputs_10_35_port, Y(34) => 
                           MuxOutputs_10_34_port, Y(33) => 
                           MuxOutputs_10_33_port, Y(32) => 
                           MuxOutputs_10_32_port, Y(31) => 
                           MuxOutputs_10_31_port, Y(30) => 
                           MuxOutputs_10_30_port, Y(29) => 
                           MuxOutputs_10_29_port, Y(28) => 
                           MuxOutputs_10_28_port, Y(27) => 
                           MuxOutputs_10_27_port, Y(26) => 
                           MuxOutputs_10_26_port, Y(25) => 
                           MuxOutputs_10_25_port, Y(24) => 
                           MuxOutputs_10_24_port, Y(23) => 
                           MuxOutputs_10_23_port, Y(22) => 
                           MuxOutputs_10_22_port, Y(21) => 
                           MuxOutputs_10_21_port, Y(20) => 
                           MuxOutputs_10_20_port, Y(19) => 
                           MuxOutputs_10_19_port, Y(18) => 
                           MuxOutputs_10_18_port, Y(17) => 
                           MuxOutputs_10_17_port, Y(16) => 
                           MuxOutputs_10_16_port, Y(15) => 
                           MuxOutputs_10_15_port, Y(14) => 
                           MuxOutputs_10_14_port, Y(13) => 
                           MuxOutputs_10_13_port, Y(12) => 
                           MuxOutputs_10_12_port, Y(11) => 
                           MuxOutputs_10_11_port, Y(10) => 
                           MuxOutputs_10_10_port, Y(9) => MuxOutputs_10_9_port,
                           Y(8) => MuxOutputs_10_8_port, Y(7) => 
                           MuxOutputs_10_7_port, Y(6) => MuxOutputs_10_6_port, 
                           Y(5) => MuxOutputs_10_5_port, Y(4) => 
                           MuxOutputs_10_4_port, Y(3) => MuxOutputs_10_3_port, 
                           Y(2) => MuxOutputs_10_2_port, Y(1) => 
                           MuxOutputs_10_1_port, Y(0) => MuxOutputs_10_0_port);
   encoderI_11 : encoder_21 port map( pieceofB(2) => B(23), pieceofB(1) => 
                           B(22), pieceofB(0) => B(21), sel(2) => sel_11_2_port
                           , sel(1) => sel_11_1_port, sel(0) => sel_11_0_port);
   MUXI_11 : MUX51_MuxNbit64_21 port map( zeroSignal(63) => X_Logic0_port, 
                           zeroSignal(62) => X_Logic0_port, zeroSignal(61) => 
                           X_Logic0_port, zeroSignal(60) => X_Logic0_port, 
                           zeroSignal(59) => X_Logic0_port, zeroSignal(58) => 
                           X_Logic0_port, zeroSignal(57) => X_Logic0_port, 
                           zeroSignal(56) => X_Logic0_port, zeroSignal(55) => 
                           X_Logic0_port, zeroSignal(54) => X_Logic0_port, 
                           zeroSignal(53) => X_Logic0_port, zeroSignal(52) => 
                           X_Logic0_port, zeroSignal(51) => X_Logic0_port, 
                           zeroSignal(50) => X_Logic0_port, zeroSignal(49) => 
                           X_Logic0_port, zeroSignal(48) => X_Logic0_port, 
                           zeroSignal(47) => X_Logic0_port, zeroSignal(46) => 
                           X_Logic0_port, zeroSignal(45) => X_Logic0_port, 
                           zeroSignal(44) => X_Logic0_port, zeroSignal(43) => 
                           X_Logic0_port, zeroSignal(42) => X_Logic0_port, 
                           zeroSignal(41) => X_Logic0_port, zeroSignal(40) => 
                           X_Logic0_port, zeroSignal(39) => X_Logic0_port, 
                           zeroSignal(38) => X_Logic0_port, zeroSignal(37) => 
                           X_Logic0_port, zeroSignal(36) => X_Logic0_port, 
                           zeroSignal(35) => X_Logic0_port, zeroSignal(34) => 
                           X_Logic0_port, zeroSignal(33) => X_Logic0_port, 
                           zeroSignal(32) => X_Logic0_port, zeroSignal(31) => 
                           X_Logic0_port, zeroSignal(30) => X_Logic0_port, 
                           zeroSignal(29) => X_Logic0_port, zeroSignal(28) => 
                           X_Logic0_port, zeroSignal(27) => X_Logic0_port, 
                           zeroSignal(26) => X_Logic0_port, zeroSignal(25) => 
                           X_Logic0_port, zeroSignal(24) => X_Logic0_port, 
                           zeroSignal(23) => X_Logic0_port, zeroSignal(22) => 
                           X_Logic0_port, zeroSignal(21) => X_Logic0_port, 
                           zeroSignal(20) => X_Logic0_port, zeroSignal(19) => 
                           X_Logic0_port, zeroSignal(18) => X_Logic0_port, 
                           zeroSignal(17) => X_Logic0_port, zeroSignal(16) => 
                           X_Logic0_port, zeroSignal(15) => X_Logic0_port, 
                           zeroSignal(14) => X_Logic0_port, zeroSignal(13) => 
                           X_Logic0_port, zeroSignal(12) => X_Logic0_port, 
                           zeroSignal(11) => X_Logic0_port, zeroSignal(10) => 
                           X_Logic0_port, zeroSignal(9) => X_Logic0_port, 
                           zeroSignal(8) => X_Logic0_port, zeroSignal(7) => 
                           X_Logic0_port, zeroSignal(6) => X_Logic0_port, 
                           zeroSignal(5) => X_Logic0_port, zeroSignal(4) => 
                           X_Logic0_port, zeroSignal(3) => X_Logic0_port, 
                           zeroSignal(2) => X_Logic0_port, zeroSignal(1) => 
                           X_Logic0_port, zeroSignal(0) => X_Logic0_port, 
                           A_signal(63) => positive_inputs_22_63_port, 
                           A_signal(62) => positive_inputs_22_62_port, 
                           A_signal(61) => positive_inputs_22_61_port, 
                           A_signal(60) => positive_inputs_22_60_port, 
                           A_signal(59) => positive_inputs_22_59_port, 
                           A_signal(58) => positive_inputs_22_58_port, 
                           A_signal(57) => positive_inputs_22_57_port, 
                           A_signal(56) => positive_inputs_22_56_port, 
                           A_signal(55) => positive_inputs_22_55_port, 
                           A_signal(54) => positive_inputs_22_54_port, 
                           A_signal(53) => positive_inputs_22_53_port, 
                           A_signal(52) => positive_inputs_22_52_port, 
                           A_signal(51) => positive_inputs_22_51_port, 
                           A_signal(50) => positive_inputs_22_50_port, 
                           A_signal(49) => positive_inputs_22_49_port, 
                           A_signal(48) => positive_inputs_22_48_port, 
                           A_signal(47) => positive_inputs_22_47_port, 
                           A_signal(46) => positive_inputs_22_46_port, 
                           A_signal(45) => positive_inputs_22_45_port, 
                           A_signal(44) => positive_inputs_22_44_port, 
                           A_signal(43) => positive_inputs_22_43_port, 
                           A_signal(42) => positive_inputs_22_42_port, 
                           A_signal(41) => positive_inputs_22_41_port, 
                           A_signal(40) => positive_inputs_22_40_port, 
                           A_signal(39) => positive_inputs_22_39_port, 
                           A_signal(38) => positive_inputs_22_38_port, 
                           A_signal(37) => positive_inputs_22_37_port, 
                           A_signal(36) => positive_inputs_22_36_port, 
                           A_signal(35) => positive_inputs_22_35_port, 
                           A_signal(34) => positive_inputs_22_34_port, 
                           A_signal(33) => positive_inputs_22_33_port, 
                           A_signal(32) => positive_inputs_22_32_port, 
                           A_signal(31) => positive_inputs_22_31_port, 
                           A_signal(30) => positive_inputs_22_30_port, 
                           A_signal(29) => positive_inputs_22_29_port, 
                           A_signal(28) => positive_inputs_22_28_port, 
                           A_signal(27) => positive_inputs_22_27_port, 
                           A_signal(26) => positive_inputs_22_26_port, 
                           A_signal(25) => positive_inputs_22_25_port, 
                           A_signal(24) => positive_inputs_22_24_port, 
                           A_signal(23) => positive_inputs_22_23_port, 
                           A_signal(22) => positive_inputs_22_22_port, 
                           A_signal(21) => positive_inputs_22_21_port, 
                           A_signal(20) => positive_inputs_22_20_port, 
                           A_signal(19) => positive_inputs_22_19_port, 
                           A_signal(18) => positive_inputs_22_18_port, 
                           A_signal(17) => positive_inputs_22_17_port, 
                           A_signal(16) => positive_inputs_22_16_port, 
                           A_signal(15) => positive_inputs_22_15_port, 
                           A_signal(14) => positive_inputs_22_14_port, 
                           A_signal(13) => positive_inputs_22_13_port, 
                           A_signal(12) => positive_inputs_22_12_port, 
                           A_signal(11) => positive_inputs_22_11_port, 
                           A_signal(10) => positive_inputs_22_10_port, 
                           A_signal(9) => positive_inputs_22_9_port, 
                           A_signal(8) => positive_inputs_22_8_port, 
                           A_signal(7) => positive_inputs_22_7_port, 
                           A_signal(6) => positive_inputs_22_6_port, 
                           A_signal(5) => positive_inputs_22_5_port, 
                           A_signal(4) => positive_inputs_22_4_port, 
                           A_signal(3) => positive_inputs_22_3_port, 
                           A_signal(2) => positive_inputs_22_2_port, 
                           A_signal(1) => positive_inputs_22_1_port, 
                           A_signal(0) => n8, A_neg(63) => 
                           negative_inputs_22_63_port, A_neg(62) => 
                           negative_inputs_22_62_port, A_neg(61) => 
                           negative_inputs_22_61_port, A_neg(60) => 
                           negative_inputs_22_60_port, A_neg(59) => 
                           negative_inputs_22_59_port, A_neg(58) => 
                           negative_inputs_22_58_port, A_neg(57) => 
                           negative_inputs_22_57_port, A_neg(56) => 
                           negative_inputs_22_56_port, A_neg(55) => 
                           negative_inputs_22_55_port, A_neg(54) => 
                           negative_inputs_22_54_port, A_neg(53) => 
                           negative_inputs_22_53_port, A_neg(52) => 
                           negative_inputs_22_52_port, A_neg(51) => 
                           negative_inputs_22_51_port, A_neg(50) => 
                           negative_inputs_22_50_port, A_neg(49) => 
                           negative_inputs_22_49_port, A_neg(48) => 
                           negative_inputs_22_48_port, A_neg(47) => 
                           negative_inputs_22_47_port, A_neg(46) => 
                           negative_inputs_22_46_port, A_neg(45) => 
                           negative_inputs_22_45_port, A_neg(44) => 
                           negative_inputs_22_44_port, A_neg(43) => 
                           negative_inputs_22_43_port, A_neg(42) => 
                           negative_inputs_22_42_port, A_neg(41) => 
                           negative_inputs_22_41_port, A_neg(40) => 
                           negative_inputs_22_40_port, A_neg(39) => 
                           negative_inputs_22_39_port, A_neg(38) => 
                           negative_inputs_22_38_port, A_neg(37) => 
                           negative_inputs_22_37_port, A_neg(36) => 
                           negative_inputs_22_36_port, A_neg(35) => 
                           negative_inputs_22_35_port, A_neg(34) => 
                           negative_inputs_22_34_port, A_neg(33) => 
                           negative_inputs_22_33_port, A_neg(32) => 
                           negative_inputs_22_32_port, A_neg(31) => 
                           negative_inputs_22_31_port, A_neg(30) => 
                           negative_inputs_22_30_port, A_neg(29) => 
                           negative_inputs_22_29_port, A_neg(28) => 
                           negative_inputs_22_28_port, A_neg(27) => 
                           negative_inputs_22_27_port, A_neg(26) => 
                           negative_inputs_22_26_port, A_neg(25) => 
                           negative_inputs_22_25_port, A_neg(24) => 
                           negative_inputs_22_24_port, A_neg(23) => 
                           negative_inputs_22_23_port, A_neg(22) => 
                           negative_inputs_22_22_port, A_neg(21) => 
                           negative_inputs_22_21_port, A_neg(20) => 
                           negative_inputs_22_20_port, A_neg(19) => 
                           negative_inputs_22_19_port, A_neg(18) => 
                           negative_inputs_22_18_port, A_neg(17) => 
                           negative_inputs_22_17_port, A_neg(16) => 
                           negative_inputs_22_16_port, A_neg(15) => 
                           negative_inputs_22_15_port, A_neg(14) => 
                           negative_inputs_22_14_port, A_neg(13) => 
                           negative_inputs_22_13_port, A_neg(12) => 
                           negative_inputs_22_12_port, A_neg(11) => 
                           negative_inputs_22_11_port, A_neg(10) => 
                           negative_inputs_22_10_port, A_neg(9) => 
                           negative_inputs_22_9_port, A_neg(8) => 
                           negative_inputs_22_8_port, A_neg(7) => 
                           negative_inputs_22_7_port, A_neg(6) => 
                           negative_inputs_22_6_port, A_neg(5) => 
                           negative_inputs_22_5_port, A_neg(4) => 
                           negative_inputs_22_4_port, A_neg(3) => 
                           negative_inputs_22_3_port, A_neg(2) => 
                           negative_inputs_22_2_port, A_neg(1) => 
                           negative_inputs_22_1_port, A_neg(0) => n8, 
                           A_shifted(63) => positive_inputs_23_63_port, 
                           A_shifted(62) => positive_inputs_23_62_port, 
                           A_shifted(61) => positive_inputs_23_61_port, 
                           A_shifted(60) => positive_inputs_23_60_port, 
                           A_shifted(59) => positive_inputs_23_59_port, 
                           A_shifted(58) => positive_inputs_23_58_port, 
                           A_shifted(57) => positive_inputs_23_57_port, 
                           A_shifted(56) => positive_inputs_23_56_port, 
                           A_shifted(55) => positive_inputs_23_55_port, 
                           A_shifted(54) => positive_inputs_23_54_port, 
                           A_shifted(53) => positive_inputs_23_53_port, 
                           A_shifted(52) => positive_inputs_23_52_port, 
                           A_shifted(51) => positive_inputs_23_51_port, 
                           A_shifted(50) => positive_inputs_23_50_port, 
                           A_shifted(49) => positive_inputs_23_49_port, 
                           A_shifted(48) => positive_inputs_23_48_port, 
                           A_shifted(47) => positive_inputs_23_47_port, 
                           A_shifted(46) => positive_inputs_23_46_port, 
                           A_shifted(45) => positive_inputs_23_45_port, 
                           A_shifted(44) => positive_inputs_23_44_port, 
                           A_shifted(43) => positive_inputs_23_43_port, 
                           A_shifted(42) => positive_inputs_23_42_port, 
                           A_shifted(41) => positive_inputs_23_41_port, 
                           A_shifted(40) => positive_inputs_23_40_port, 
                           A_shifted(39) => positive_inputs_23_39_port, 
                           A_shifted(38) => positive_inputs_23_38_port, 
                           A_shifted(37) => positive_inputs_23_37_port, 
                           A_shifted(36) => positive_inputs_23_36_port, 
                           A_shifted(35) => positive_inputs_23_35_port, 
                           A_shifted(34) => positive_inputs_23_34_port, 
                           A_shifted(33) => positive_inputs_23_33_port, 
                           A_shifted(32) => positive_inputs_23_32_port, 
                           A_shifted(31) => positive_inputs_23_31_port, 
                           A_shifted(30) => positive_inputs_23_30_port, 
                           A_shifted(29) => positive_inputs_23_29_port, 
                           A_shifted(28) => positive_inputs_23_28_port, 
                           A_shifted(27) => positive_inputs_23_27_port, 
                           A_shifted(26) => positive_inputs_23_26_port, 
                           A_shifted(25) => positive_inputs_23_25_port, 
                           A_shifted(24) => positive_inputs_23_24_port, 
                           A_shifted(23) => positive_inputs_23_23_port, 
                           A_shifted(22) => positive_inputs_23_22_port, 
                           A_shifted(21) => positive_inputs_23_21_port, 
                           A_shifted(20) => positive_inputs_23_20_port, 
                           A_shifted(19) => positive_inputs_23_19_port, 
                           A_shifted(18) => positive_inputs_23_18_port, 
                           A_shifted(17) => positive_inputs_23_17_port, 
                           A_shifted(16) => positive_inputs_23_16_port, 
                           A_shifted(15) => positive_inputs_23_15_port, 
                           A_shifted(14) => positive_inputs_23_14_port, 
                           A_shifted(13) => positive_inputs_23_13_port, 
                           A_shifted(12) => positive_inputs_23_12_port, 
                           A_shifted(11) => positive_inputs_23_11_port, 
                           A_shifted(10) => positive_inputs_23_10_port, 
                           A_shifted(9) => positive_inputs_23_9_port, 
                           A_shifted(8) => positive_inputs_23_8_port, 
                           A_shifted(7) => positive_inputs_23_7_port, 
                           A_shifted(6) => positive_inputs_23_6_port, 
                           A_shifted(5) => positive_inputs_23_5_port, 
                           A_shifted(4) => positive_inputs_23_4_port, 
                           A_shifted(3) => positive_inputs_23_3_port, 
                           A_shifted(2) => positive_inputs_23_2_port, 
                           A_shifted(1) => positive_inputs_23_1_port, 
                           A_shifted(0) => n8, A_neg_shifted(63) => 
                           negative_inputs_23_63_port, A_neg_shifted(62) => 
                           negative_inputs_23_62_port, A_neg_shifted(61) => 
                           negative_inputs_23_61_port, A_neg_shifted(60) => 
                           negative_inputs_23_60_port, A_neg_shifted(59) => 
                           negative_inputs_23_59_port, A_neg_shifted(58) => 
                           negative_inputs_23_58_port, A_neg_shifted(57) => 
                           negative_inputs_23_57_port, A_neg_shifted(56) => 
                           negative_inputs_23_56_port, A_neg_shifted(55) => 
                           negative_inputs_23_55_port, A_neg_shifted(54) => 
                           negative_inputs_23_54_port, A_neg_shifted(53) => 
                           negative_inputs_23_53_port, A_neg_shifted(52) => 
                           negative_inputs_23_52_port, A_neg_shifted(51) => 
                           negative_inputs_23_51_port, A_neg_shifted(50) => 
                           negative_inputs_23_50_port, A_neg_shifted(49) => 
                           negative_inputs_23_49_port, A_neg_shifted(48) => 
                           negative_inputs_23_48_port, A_neg_shifted(47) => 
                           negative_inputs_23_47_port, A_neg_shifted(46) => 
                           negative_inputs_23_46_port, A_neg_shifted(45) => 
                           negative_inputs_23_45_port, A_neg_shifted(44) => 
                           negative_inputs_23_44_port, A_neg_shifted(43) => 
                           negative_inputs_23_43_port, A_neg_shifted(42) => 
                           negative_inputs_23_42_port, A_neg_shifted(41) => 
                           negative_inputs_23_41_port, A_neg_shifted(40) => 
                           negative_inputs_23_40_port, A_neg_shifted(39) => 
                           negative_inputs_23_39_port, A_neg_shifted(38) => 
                           negative_inputs_23_38_port, A_neg_shifted(37) => 
                           negative_inputs_23_37_port, A_neg_shifted(36) => 
                           negative_inputs_23_36_port, A_neg_shifted(35) => 
                           negative_inputs_23_35_port, A_neg_shifted(34) => 
                           negative_inputs_23_34_port, A_neg_shifted(33) => 
                           negative_inputs_23_33_port, A_neg_shifted(32) => 
                           negative_inputs_23_32_port, A_neg_shifted(31) => 
                           negative_inputs_23_31_port, A_neg_shifted(30) => 
                           negative_inputs_23_30_port, A_neg_shifted(29) => 
                           negative_inputs_23_29_port, A_neg_shifted(28) => 
                           negative_inputs_23_28_port, A_neg_shifted(27) => 
                           negative_inputs_23_27_port, A_neg_shifted(26) => 
                           negative_inputs_23_26_port, A_neg_shifted(25) => 
                           negative_inputs_23_25_port, A_neg_shifted(24) => 
                           negative_inputs_23_24_port, A_neg_shifted(23) => 
                           negative_inputs_23_23_port, A_neg_shifted(22) => 
                           negative_inputs_23_22_port, A_neg_shifted(21) => 
                           negative_inputs_23_21_port, A_neg_shifted(20) => 
                           negative_inputs_23_20_port, A_neg_shifted(19) => 
                           negative_inputs_23_19_port, A_neg_shifted(18) => 
                           negative_inputs_23_18_port, A_neg_shifted(17) => 
                           negative_inputs_23_17_port, A_neg_shifted(16) => 
                           negative_inputs_23_16_port, A_neg_shifted(15) => 
                           negative_inputs_23_15_port, A_neg_shifted(14) => 
                           negative_inputs_23_14_port, A_neg_shifted(13) => 
                           negative_inputs_23_13_port, A_neg_shifted(12) => 
                           negative_inputs_23_12_port, A_neg_shifted(11) => 
                           negative_inputs_23_11_port, A_neg_shifted(10) => 
                           negative_inputs_23_10_port, A_neg_shifted(9) => 
                           negative_inputs_23_9_port, A_neg_shifted(8) => 
                           negative_inputs_23_8_port, A_neg_shifted(7) => 
                           negative_inputs_23_7_port, A_neg_shifted(6) => 
                           negative_inputs_23_6_port, A_neg_shifted(5) => 
                           negative_inputs_23_5_port, A_neg_shifted(4) => 
                           negative_inputs_23_4_port, A_neg_shifted(3) => 
                           negative_inputs_23_3_port, A_neg_shifted(2) => 
                           negative_inputs_23_2_port, A_neg_shifted(1) => 
                           negative_inputs_23_1_port, A_neg_shifted(0) => n8, 
                           Sel(2) => sel_11_2_port, Sel(1) => sel_11_1_port, 
                           Sel(0) => sel_11_0_port, Y(63) => 
                           MuxOutputs_11_63_port, Y(62) => 
                           MuxOutputs_11_62_port, Y(61) => 
                           MuxOutputs_11_61_port, Y(60) => 
                           MuxOutputs_11_60_port, Y(59) => 
                           MuxOutputs_11_59_port, Y(58) => 
                           MuxOutputs_11_58_port, Y(57) => 
                           MuxOutputs_11_57_port, Y(56) => 
                           MuxOutputs_11_56_port, Y(55) => 
                           MuxOutputs_11_55_port, Y(54) => 
                           MuxOutputs_11_54_port, Y(53) => 
                           MuxOutputs_11_53_port, Y(52) => 
                           MuxOutputs_11_52_port, Y(51) => 
                           MuxOutputs_11_51_port, Y(50) => 
                           MuxOutputs_11_50_port, Y(49) => 
                           MuxOutputs_11_49_port, Y(48) => 
                           MuxOutputs_11_48_port, Y(47) => 
                           MuxOutputs_11_47_port, Y(46) => 
                           MuxOutputs_11_46_port, Y(45) => 
                           MuxOutputs_11_45_port, Y(44) => 
                           MuxOutputs_11_44_port, Y(43) => 
                           MuxOutputs_11_43_port, Y(42) => 
                           MuxOutputs_11_42_port, Y(41) => 
                           MuxOutputs_11_41_port, Y(40) => 
                           MuxOutputs_11_40_port, Y(39) => 
                           MuxOutputs_11_39_port, Y(38) => 
                           MuxOutputs_11_38_port, Y(37) => 
                           MuxOutputs_11_37_port, Y(36) => 
                           MuxOutputs_11_36_port, Y(35) => 
                           MuxOutputs_11_35_port, Y(34) => 
                           MuxOutputs_11_34_port, Y(33) => 
                           MuxOutputs_11_33_port, Y(32) => 
                           MuxOutputs_11_32_port, Y(31) => 
                           MuxOutputs_11_31_port, Y(30) => 
                           MuxOutputs_11_30_port, Y(29) => 
                           MuxOutputs_11_29_port, Y(28) => 
                           MuxOutputs_11_28_port, Y(27) => 
                           MuxOutputs_11_27_port, Y(26) => 
                           MuxOutputs_11_26_port, Y(25) => 
                           MuxOutputs_11_25_port, Y(24) => 
                           MuxOutputs_11_24_port, Y(23) => 
                           MuxOutputs_11_23_port, Y(22) => 
                           MuxOutputs_11_22_port, Y(21) => 
                           MuxOutputs_11_21_port, Y(20) => 
                           MuxOutputs_11_20_port, Y(19) => 
                           MuxOutputs_11_19_port, Y(18) => 
                           MuxOutputs_11_18_port, Y(17) => 
                           MuxOutputs_11_17_port, Y(16) => 
                           MuxOutputs_11_16_port, Y(15) => 
                           MuxOutputs_11_15_port, Y(14) => 
                           MuxOutputs_11_14_port, Y(13) => 
                           MuxOutputs_11_13_port, Y(12) => 
                           MuxOutputs_11_12_port, Y(11) => 
                           MuxOutputs_11_11_port, Y(10) => 
                           MuxOutputs_11_10_port, Y(9) => MuxOutputs_11_9_port,
                           Y(8) => MuxOutputs_11_8_port, Y(7) => 
                           MuxOutputs_11_7_port, Y(6) => MuxOutputs_11_6_port, 
                           Y(5) => MuxOutputs_11_5_port, Y(4) => 
                           MuxOutputs_11_4_port, Y(3) => MuxOutputs_11_3_port, 
                           Y(2) => MuxOutputs_11_2_port, Y(1) => 
                           MuxOutputs_11_1_port, Y(0) => MuxOutputs_11_0_port);
   encoderI_12 : encoder_20 port map( pieceofB(2) => B(25), pieceofB(1) => 
                           B(24), pieceofB(0) => B(23), sel(2) => sel_12_2_port
                           , sel(1) => sel_12_1_port, sel(0) => sel_12_0_port);
   MUXI_12 : MUX51_MuxNbit64_20 port map( zeroSignal(63) => X_Logic0_port, 
                           zeroSignal(62) => X_Logic0_port, zeroSignal(61) => 
                           X_Logic0_port, zeroSignal(60) => X_Logic0_port, 
                           zeroSignal(59) => X_Logic0_port, zeroSignal(58) => 
                           X_Logic0_port, zeroSignal(57) => X_Logic0_port, 
                           zeroSignal(56) => X_Logic0_port, zeroSignal(55) => 
                           X_Logic0_port, zeroSignal(54) => X_Logic0_port, 
                           zeroSignal(53) => X_Logic0_port, zeroSignal(52) => 
                           X_Logic0_port, zeroSignal(51) => X_Logic0_port, 
                           zeroSignal(50) => X_Logic0_port, zeroSignal(49) => 
                           X_Logic0_port, zeroSignal(48) => X_Logic0_port, 
                           zeroSignal(47) => X_Logic0_port, zeroSignal(46) => 
                           X_Logic0_port, zeroSignal(45) => X_Logic0_port, 
                           zeroSignal(44) => X_Logic0_port, zeroSignal(43) => 
                           X_Logic0_port, zeroSignal(42) => X_Logic0_port, 
                           zeroSignal(41) => X_Logic0_port, zeroSignal(40) => 
                           X_Logic0_port, zeroSignal(39) => X_Logic0_port, 
                           zeroSignal(38) => X_Logic0_port, zeroSignal(37) => 
                           X_Logic0_port, zeroSignal(36) => X_Logic0_port, 
                           zeroSignal(35) => X_Logic0_port, zeroSignal(34) => 
                           X_Logic0_port, zeroSignal(33) => X_Logic0_port, 
                           zeroSignal(32) => X_Logic0_port, zeroSignal(31) => 
                           X_Logic0_port, zeroSignal(30) => X_Logic0_port, 
                           zeroSignal(29) => X_Logic0_port, zeroSignal(28) => 
                           X_Logic0_port, zeroSignal(27) => X_Logic0_port, 
                           zeroSignal(26) => X_Logic0_port, zeroSignal(25) => 
                           X_Logic0_port, zeroSignal(24) => X_Logic0_port, 
                           zeroSignal(23) => X_Logic0_port, zeroSignal(22) => 
                           X_Logic0_port, zeroSignal(21) => X_Logic0_port, 
                           zeroSignal(20) => X_Logic0_port, zeroSignal(19) => 
                           X_Logic0_port, zeroSignal(18) => X_Logic0_port, 
                           zeroSignal(17) => X_Logic0_port, zeroSignal(16) => 
                           X_Logic0_port, zeroSignal(15) => X_Logic0_port, 
                           zeroSignal(14) => X_Logic0_port, zeroSignal(13) => 
                           X_Logic0_port, zeroSignal(12) => X_Logic0_port, 
                           zeroSignal(11) => X_Logic0_port, zeroSignal(10) => 
                           X_Logic0_port, zeroSignal(9) => X_Logic0_port, 
                           zeroSignal(8) => X_Logic0_port, zeroSignal(7) => 
                           X_Logic0_port, zeroSignal(6) => X_Logic0_port, 
                           zeroSignal(5) => X_Logic0_port, zeroSignal(4) => 
                           X_Logic0_port, zeroSignal(3) => X_Logic0_port, 
                           zeroSignal(2) => X_Logic0_port, zeroSignal(1) => 
                           X_Logic0_port, zeroSignal(0) => X_Logic0_port, 
                           A_signal(63) => positive_inputs_24_63_port, 
                           A_signal(62) => positive_inputs_24_62_port, 
                           A_signal(61) => positive_inputs_24_61_port, 
                           A_signal(60) => positive_inputs_24_60_port, 
                           A_signal(59) => positive_inputs_24_59_port, 
                           A_signal(58) => positive_inputs_24_58_port, 
                           A_signal(57) => positive_inputs_24_57_port, 
                           A_signal(56) => positive_inputs_24_56_port, 
                           A_signal(55) => positive_inputs_24_55_port, 
                           A_signal(54) => positive_inputs_24_54_port, 
                           A_signal(53) => positive_inputs_24_53_port, 
                           A_signal(52) => positive_inputs_24_52_port, 
                           A_signal(51) => positive_inputs_24_51_port, 
                           A_signal(50) => positive_inputs_24_50_port, 
                           A_signal(49) => positive_inputs_24_49_port, 
                           A_signal(48) => positive_inputs_24_48_port, 
                           A_signal(47) => positive_inputs_24_47_port, 
                           A_signal(46) => positive_inputs_24_46_port, 
                           A_signal(45) => positive_inputs_24_45_port, 
                           A_signal(44) => positive_inputs_24_44_port, 
                           A_signal(43) => positive_inputs_24_43_port, 
                           A_signal(42) => positive_inputs_24_42_port, 
                           A_signal(41) => positive_inputs_24_41_port, 
                           A_signal(40) => positive_inputs_24_40_port, 
                           A_signal(39) => positive_inputs_24_39_port, 
                           A_signal(38) => positive_inputs_24_38_port, 
                           A_signal(37) => positive_inputs_24_37_port, 
                           A_signal(36) => positive_inputs_24_36_port, 
                           A_signal(35) => positive_inputs_24_35_port, 
                           A_signal(34) => positive_inputs_24_34_port, 
                           A_signal(33) => positive_inputs_24_33_port, 
                           A_signal(32) => positive_inputs_24_32_port, 
                           A_signal(31) => positive_inputs_24_31_port, 
                           A_signal(30) => positive_inputs_24_30_port, 
                           A_signal(29) => positive_inputs_24_29_port, 
                           A_signal(28) => positive_inputs_24_28_port, 
                           A_signal(27) => positive_inputs_24_27_port, 
                           A_signal(26) => positive_inputs_24_26_port, 
                           A_signal(25) => positive_inputs_24_25_port, 
                           A_signal(24) => positive_inputs_24_24_port, 
                           A_signal(23) => positive_inputs_24_23_port, 
                           A_signal(22) => positive_inputs_24_22_port, 
                           A_signal(21) => positive_inputs_24_21_port, 
                           A_signal(20) => positive_inputs_24_20_port, 
                           A_signal(19) => positive_inputs_24_19_port, 
                           A_signal(18) => positive_inputs_24_18_port, 
                           A_signal(17) => positive_inputs_24_17_port, 
                           A_signal(16) => positive_inputs_24_16_port, 
                           A_signal(15) => positive_inputs_24_15_port, 
                           A_signal(14) => positive_inputs_24_14_port, 
                           A_signal(13) => positive_inputs_24_13_port, 
                           A_signal(12) => positive_inputs_24_12_port, 
                           A_signal(11) => positive_inputs_24_11_port, 
                           A_signal(10) => positive_inputs_24_10_port, 
                           A_signal(9) => positive_inputs_24_9_port, 
                           A_signal(8) => positive_inputs_24_8_port, 
                           A_signal(7) => positive_inputs_24_7_port, 
                           A_signal(6) => positive_inputs_24_6_port, 
                           A_signal(5) => positive_inputs_24_5_port, 
                           A_signal(4) => positive_inputs_24_4_port, 
                           A_signal(3) => positive_inputs_24_3_port, 
                           A_signal(2) => positive_inputs_24_2_port, 
                           A_signal(1) => positive_inputs_24_1_port, 
                           A_signal(0) => n8, A_neg(63) => 
                           negative_inputs_24_63_port, A_neg(62) => 
                           negative_inputs_24_62_port, A_neg(61) => 
                           negative_inputs_24_61_port, A_neg(60) => 
                           negative_inputs_24_60_port, A_neg(59) => 
                           negative_inputs_24_59_port, A_neg(58) => 
                           negative_inputs_24_58_port, A_neg(57) => 
                           negative_inputs_24_57_port, A_neg(56) => 
                           negative_inputs_24_56_port, A_neg(55) => 
                           negative_inputs_24_55_port, A_neg(54) => 
                           negative_inputs_24_54_port, A_neg(53) => 
                           negative_inputs_24_53_port, A_neg(52) => 
                           negative_inputs_24_52_port, A_neg(51) => 
                           negative_inputs_24_51_port, A_neg(50) => 
                           negative_inputs_24_50_port, A_neg(49) => 
                           negative_inputs_24_49_port, A_neg(48) => 
                           negative_inputs_24_48_port, A_neg(47) => 
                           negative_inputs_24_47_port, A_neg(46) => 
                           negative_inputs_24_46_port, A_neg(45) => 
                           negative_inputs_24_45_port, A_neg(44) => 
                           negative_inputs_24_44_port, A_neg(43) => 
                           negative_inputs_24_43_port, A_neg(42) => 
                           negative_inputs_24_42_port, A_neg(41) => 
                           negative_inputs_24_41_port, A_neg(40) => 
                           negative_inputs_24_40_port, A_neg(39) => 
                           negative_inputs_24_39_port, A_neg(38) => 
                           negative_inputs_24_38_port, A_neg(37) => 
                           negative_inputs_24_37_port, A_neg(36) => 
                           negative_inputs_24_36_port, A_neg(35) => 
                           negative_inputs_24_35_port, A_neg(34) => 
                           negative_inputs_24_34_port, A_neg(33) => 
                           negative_inputs_24_33_port, A_neg(32) => 
                           negative_inputs_24_32_port, A_neg(31) => 
                           negative_inputs_24_31_port, A_neg(30) => 
                           negative_inputs_24_30_port, A_neg(29) => 
                           negative_inputs_24_29_port, A_neg(28) => 
                           negative_inputs_24_28_port, A_neg(27) => 
                           negative_inputs_24_27_port, A_neg(26) => 
                           negative_inputs_24_26_port, A_neg(25) => 
                           negative_inputs_24_25_port, A_neg(24) => 
                           negative_inputs_24_24_port, A_neg(23) => 
                           negative_inputs_24_23_port, A_neg(22) => 
                           negative_inputs_24_22_port, A_neg(21) => 
                           negative_inputs_24_21_port, A_neg(20) => 
                           negative_inputs_24_20_port, A_neg(19) => 
                           negative_inputs_24_19_port, A_neg(18) => 
                           negative_inputs_24_18_port, A_neg(17) => 
                           negative_inputs_24_17_port, A_neg(16) => 
                           negative_inputs_24_16_port, A_neg(15) => 
                           negative_inputs_24_15_port, A_neg(14) => 
                           negative_inputs_24_14_port, A_neg(13) => 
                           negative_inputs_24_13_port, A_neg(12) => 
                           negative_inputs_24_12_port, A_neg(11) => 
                           negative_inputs_24_11_port, A_neg(10) => 
                           negative_inputs_24_10_port, A_neg(9) => 
                           negative_inputs_24_9_port, A_neg(8) => 
                           negative_inputs_24_8_port, A_neg(7) => 
                           negative_inputs_24_7_port, A_neg(6) => 
                           negative_inputs_24_6_port, A_neg(5) => 
                           negative_inputs_24_5_port, A_neg(4) => 
                           negative_inputs_24_4_port, A_neg(3) => 
                           negative_inputs_24_3_port, A_neg(2) => 
                           negative_inputs_24_2_port, A_neg(1) => 
                           negative_inputs_24_1_port, A_neg(0) => n8, 
                           A_shifted(63) => positive_inputs_25_63_port, 
                           A_shifted(62) => positive_inputs_25_62_port, 
                           A_shifted(61) => positive_inputs_25_61_port, 
                           A_shifted(60) => positive_inputs_25_60_port, 
                           A_shifted(59) => positive_inputs_25_59_port, 
                           A_shifted(58) => positive_inputs_25_58_port, 
                           A_shifted(57) => positive_inputs_25_57_port, 
                           A_shifted(56) => positive_inputs_25_56_port, 
                           A_shifted(55) => positive_inputs_25_55_port, 
                           A_shifted(54) => positive_inputs_25_54_port, 
                           A_shifted(53) => positive_inputs_25_53_port, 
                           A_shifted(52) => positive_inputs_25_52_port, 
                           A_shifted(51) => positive_inputs_25_51_port, 
                           A_shifted(50) => positive_inputs_25_50_port, 
                           A_shifted(49) => positive_inputs_25_49_port, 
                           A_shifted(48) => positive_inputs_25_48_port, 
                           A_shifted(47) => positive_inputs_25_47_port, 
                           A_shifted(46) => positive_inputs_25_46_port, 
                           A_shifted(45) => positive_inputs_25_45_port, 
                           A_shifted(44) => positive_inputs_25_44_port, 
                           A_shifted(43) => positive_inputs_25_43_port, 
                           A_shifted(42) => positive_inputs_25_42_port, 
                           A_shifted(41) => positive_inputs_25_41_port, 
                           A_shifted(40) => positive_inputs_25_40_port, 
                           A_shifted(39) => positive_inputs_25_39_port, 
                           A_shifted(38) => positive_inputs_25_38_port, 
                           A_shifted(37) => positive_inputs_25_37_port, 
                           A_shifted(36) => positive_inputs_25_36_port, 
                           A_shifted(35) => positive_inputs_25_35_port, 
                           A_shifted(34) => positive_inputs_25_34_port, 
                           A_shifted(33) => positive_inputs_25_33_port, 
                           A_shifted(32) => positive_inputs_25_32_port, 
                           A_shifted(31) => positive_inputs_25_31_port, 
                           A_shifted(30) => positive_inputs_25_30_port, 
                           A_shifted(29) => positive_inputs_25_29_port, 
                           A_shifted(28) => positive_inputs_25_28_port, 
                           A_shifted(27) => positive_inputs_25_27_port, 
                           A_shifted(26) => positive_inputs_25_26_port, 
                           A_shifted(25) => positive_inputs_25_25_port, 
                           A_shifted(24) => positive_inputs_25_24_port, 
                           A_shifted(23) => positive_inputs_25_23_port, 
                           A_shifted(22) => positive_inputs_25_22_port, 
                           A_shifted(21) => positive_inputs_25_21_port, 
                           A_shifted(20) => positive_inputs_25_20_port, 
                           A_shifted(19) => positive_inputs_25_19_port, 
                           A_shifted(18) => positive_inputs_25_18_port, 
                           A_shifted(17) => positive_inputs_25_17_port, 
                           A_shifted(16) => positive_inputs_25_16_port, 
                           A_shifted(15) => positive_inputs_25_15_port, 
                           A_shifted(14) => positive_inputs_25_14_port, 
                           A_shifted(13) => positive_inputs_25_13_port, 
                           A_shifted(12) => positive_inputs_25_12_port, 
                           A_shifted(11) => positive_inputs_25_11_port, 
                           A_shifted(10) => positive_inputs_25_10_port, 
                           A_shifted(9) => positive_inputs_25_9_port, 
                           A_shifted(8) => positive_inputs_25_8_port, 
                           A_shifted(7) => positive_inputs_25_7_port, 
                           A_shifted(6) => positive_inputs_25_6_port, 
                           A_shifted(5) => positive_inputs_25_5_port, 
                           A_shifted(4) => positive_inputs_25_4_port, 
                           A_shifted(3) => positive_inputs_25_3_port, 
                           A_shifted(2) => positive_inputs_25_2_port, 
                           A_shifted(1) => positive_inputs_25_1_port, 
                           A_shifted(0) => n8, A_neg_shifted(63) => 
                           negative_inputs_25_63_port, A_neg_shifted(62) => 
                           negative_inputs_25_62_port, A_neg_shifted(61) => 
                           negative_inputs_25_61_port, A_neg_shifted(60) => 
                           negative_inputs_25_60_port, A_neg_shifted(59) => 
                           negative_inputs_25_59_port, A_neg_shifted(58) => 
                           negative_inputs_25_58_port, A_neg_shifted(57) => 
                           negative_inputs_25_57_port, A_neg_shifted(56) => 
                           negative_inputs_25_56_port, A_neg_shifted(55) => 
                           negative_inputs_25_55_port, A_neg_shifted(54) => 
                           negative_inputs_25_54_port, A_neg_shifted(53) => 
                           negative_inputs_25_53_port, A_neg_shifted(52) => 
                           negative_inputs_25_52_port, A_neg_shifted(51) => 
                           negative_inputs_25_51_port, A_neg_shifted(50) => 
                           negative_inputs_25_50_port, A_neg_shifted(49) => 
                           negative_inputs_25_49_port, A_neg_shifted(48) => 
                           negative_inputs_25_48_port, A_neg_shifted(47) => 
                           negative_inputs_25_47_port, A_neg_shifted(46) => 
                           negative_inputs_25_46_port, A_neg_shifted(45) => 
                           negative_inputs_25_45_port, A_neg_shifted(44) => 
                           negative_inputs_25_44_port, A_neg_shifted(43) => 
                           negative_inputs_25_43_port, A_neg_shifted(42) => 
                           negative_inputs_25_42_port, A_neg_shifted(41) => 
                           negative_inputs_25_41_port, A_neg_shifted(40) => 
                           negative_inputs_25_40_port, A_neg_shifted(39) => 
                           negative_inputs_25_39_port, A_neg_shifted(38) => 
                           negative_inputs_25_38_port, A_neg_shifted(37) => 
                           negative_inputs_25_37_port, A_neg_shifted(36) => 
                           negative_inputs_25_36_port, A_neg_shifted(35) => 
                           negative_inputs_25_35_port, A_neg_shifted(34) => 
                           negative_inputs_25_34_port, A_neg_shifted(33) => 
                           negative_inputs_25_33_port, A_neg_shifted(32) => 
                           negative_inputs_25_32_port, A_neg_shifted(31) => 
                           negative_inputs_25_31_port, A_neg_shifted(30) => 
                           negative_inputs_25_30_port, A_neg_shifted(29) => 
                           negative_inputs_25_29_port, A_neg_shifted(28) => 
                           negative_inputs_25_28_port, A_neg_shifted(27) => 
                           negative_inputs_25_27_port, A_neg_shifted(26) => 
                           negative_inputs_25_26_port, A_neg_shifted(25) => 
                           negative_inputs_25_25_port, A_neg_shifted(24) => 
                           negative_inputs_25_24_port, A_neg_shifted(23) => 
                           negative_inputs_25_23_port, A_neg_shifted(22) => 
                           negative_inputs_25_22_port, A_neg_shifted(21) => 
                           negative_inputs_25_21_port, A_neg_shifted(20) => 
                           negative_inputs_25_20_port, A_neg_shifted(19) => 
                           negative_inputs_25_19_port, A_neg_shifted(18) => 
                           negative_inputs_25_18_port, A_neg_shifted(17) => 
                           negative_inputs_25_17_port, A_neg_shifted(16) => 
                           negative_inputs_25_16_port, A_neg_shifted(15) => 
                           negative_inputs_25_15_port, A_neg_shifted(14) => 
                           negative_inputs_25_14_port, A_neg_shifted(13) => 
                           negative_inputs_25_13_port, A_neg_shifted(12) => 
                           negative_inputs_25_12_port, A_neg_shifted(11) => 
                           negative_inputs_25_11_port, A_neg_shifted(10) => 
                           negative_inputs_25_10_port, A_neg_shifted(9) => 
                           negative_inputs_25_9_port, A_neg_shifted(8) => 
                           negative_inputs_25_8_port, A_neg_shifted(7) => 
                           negative_inputs_25_7_port, A_neg_shifted(6) => 
                           negative_inputs_25_6_port, A_neg_shifted(5) => 
                           negative_inputs_25_5_port, A_neg_shifted(4) => 
                           negative_inputs_25_4_port, A_neg_shifted(3) => 
                           negative_inputs_25_3_port, A_neg_shifted(2) => 
                           negative_inputs_25_2_port, A_neg_shifted(1) => 
                           negative_inputs_25_1_port, A_neg_shifted(0) => n8, 
                           Sel(2) => sel_12_2_port, Sel(1) => sel_12_1_port, 
                           Sel(0) => sel_12_0_port, Y(63) => 
                           MuxOutputs_12_63_port, Y(62) => 
                           MuxOutputs_12_62_port, Y(61) => 
                           MuxOutputs_12_61_port, Y(60) => 
                           MuxOutputs_12_60_port, Y(59) => 
                           MuxOutputs_12_59_port, Y(58) => 
                           MuxOutputs_12_58_port, Y(57) => 
                           MuxOutputs_12_57_port, Y(56) => 
                           MuxOutputs_12_56_port, Y(55) => 
                           MuxOutputs_12_55_port, Y(54) => 
                           MuxOutputs_12_54_port, Y(53) => 
                           MuxOutputs_12_53_port, Y(52) => 
                           MuxOutputs_12_52_port, Y(51) => 
                           MuxOutputs_12_51_port, Y(50) => 
                           MuxOutputs_12_50_port, Y(49) => 
                           MuxOutputs_12_49_port, Y(48) => 
                           MuxOutputs_12_48_port, Y(47) => 
                           MuxOutputs_12_47_port, Y(46) => 
                           MuxOutputs_12_46_port, Y(45) => 
                           MuxOutputs_12_45_port, Y(44) => 
                           MuxOutputs_12_44_port, Y(43) => 
                           MuxOutputs_12_43_port, Y(42) => 
                           MuxOutputs_12_42_port, Y(41) => 
                           MuxOutputs_12_41_port, Y(40) => 
                           MuxOutputs_12_40_port, Y(39) => 
                           MuxOutputs_12_39_port, Y(38) => 
                           MuxOutputs_12_38_port, Y(37) => 
                           MuxOutputs_12_37_port, Y(36) => 
                           MuxOutputs_12_36_port, Y(35) => 
                           MuxOutputs_12_35_port, Y(34) => 
                           MuxOutputs_12_34_port, Y(33) => 
                           MuxOutputs_12_33_port, Y(32) => 
                           MuxOutputs_12_32_port, Y(31) => 
                           MuxOutputs_12_31_port, Y(30) => 
                           MuxOutputs_12_30_port, Y(29) => 
                           MuxOutputs_12_29_port, Y(28) => 
                           MuxOutputs_12_28_port, Y(27) => 
                           MuxOutputs_12_27_port, Y(26) => 
                           MuxOutputs_12_26_port, Y(25) => 
                           MuxOutputs_12_25_port, Y(24) => 
                           MuxOutputs_12_24_port, Y(23) => 
                           MuxOutputs_12_23_port, Y(22) => 
                           MuxOutputs_12_22_port, Y(21) => 
                           MuxOutputs_12_21_port, Y(20) => 
                           MuxOutputs_12_20_port, Y(19) => 
                           MuxOutputs_12_19_port, Y(18) => 
                           MuxOutputs_12_18_port, Y(17) => 
                           MuxOutputs_12_17_port, Y(16) => 
                           MuxOutputs_12_16_port, Y(15) => 
                           MuxOutputs_12_15_port, Y(14) => 
                           MuxOutputs_12_14_port, Y(13) => 
                           MuxOutputs_12_13_port, Y(12) => 
                           MuxOutputs_12_12_port, Y(11) => 
                           MuxOutputs_12_11_port, Y(10) => 
                           MuxOutputs_12_10_port, Y(9) => MuxOutputs_12_9_port,
                           Y(8) => MuxOutputs_12_8_port, Y(7) => 
                           MuxOutputs_12_7_port, Y(6) => MuxOutputs_12_6_port, 
                           Y(5) => MuxOutputs_12_5_port, Y(4) => 
                           MuxOutputs_12_4_port, Y(3) => MuxOutputs_12_3_port, 
                           Y(2) => MuxOutputs_12_2_port, Y(1) => 
                           MuxOutputs_12_1_port, Y(0) => MuxOutputs_12_0_port);
   encoderI_13 : encoder_19 port map( pieceofB(2) => B(27), pieceofB(1) => 
                           B(26), pieceofB(0) => B(25), sel(2) => sel_13_2_port
                           , sel(1) => sel_13_1_port, sel(0) => sel_13_0_port);
   MUXI_13 : MUX51_MuxNbit64_19 port map( zeroSignal(63) => X_Logic0_port, 
                           zeroSignal(62) => X_Logic0_port, zeroSignal(61) => 
                           X_Logic0_port, zeroSignal(60) => X_Logic0_port, 
                           zeroSignal(59) => X_Logic0_port, zeroSignal(58) => 
                           X_Logic0_port, zeroSignal(57) => X_Logic0_port, 
                           zeroSignal(56) => X_Logic0_port, zeroSignal(55) => 
                           X_Logic0_port, zeroSignal(54) => X_Logic0_port, 
                           zeroSignal(53) => X_Logic0_port, zeroSignal(52) => 
                           X_Logic0_port, zeroSignal(51) => X_Logic0_port, 
                           zeroSignal(50) => X_Logic0_port, zeroSignal(49) => 
                           X_Logic0_port, zeroSignal(48) => X_Logic0_port, 
                           zeroSignal(47) => X_Logic0_port, zeroSignal(46) => 
                           X_Logic0_port, zeroSignal(45) => X_Logic0_port, 
                           zeroSignal(44) => X_Logic0_port, zeroSignal(43) => 
                           X_Logic0_port, zeroSignal(42) => X_Logic0_port, 
                           zeroSignal(41) => X_Logic0_port, zeroSignal(40) => 
                           X_Logic0_port, zeroSignal(39) => X_Logic0_port, 
                           zeroSignal(38) => X_Logic0_port, zeroSignal(37) => 
                           X_Logic0_port, zeroSignal(36) => X_Logic0_port, 
                           zeroSignal(35) => X_Logic0_port, zeroSignal(34) => 
                           X_Logic0_port, zeroSignal(33) => X_Logic0_port, 
                           zeroSignal(32) => X_Logic0_port, zeroSignal(31) => 
                           X_Logic0_port, zeroSignal(30) => X_Logic0_port, 
                           zeroSignal(29) => X_Logic0_port, zeroSignal(28) => 
                           X_Logic0_port, zeroSignal(27) => X_Logic0_port, 
                           zeroSignal(26) => X_Logic0_port, zeroSignal(25) => 
                           X_Logic0_port, zeroSignal(24) => X_Logic0_port, 
                           zeroSignal(23) => X_Logic0_port, zeroSignal(22) => 
                           X_Logic0_port, zeroSignal(21) => X_Logic0_port, 
                           zeroSignal(20) => X_Logic0_port, zeroSignal(19) => 
                           X_Logic0_port, zeroSignal(18) => X_Logic0_port, 
                           zeroSignal(17) => X_Logic0_port, zeroSignal(16) => 
                           X_Logic0_port, zeroSignal(15) => X_Logic0_port, 
                           zeroSignal(14) => X_Logic0_port, zeroSignal(13) => 
                           X_Logic0_port, zeroSignal(12) => X_Logic0_port, 
                           zeroSignal(11) => X_Logic0_port, zeroSignal(10) => 
                           X_Logic0_port, zeroSignal(9) => X_Logic0_port, 
                           zeroSignal(8) => X_Logic0_port, zeroSignal(7) => 
                           X_Logic0_port, zeroSignal(6) => X_Logic0_port, 
                           zeroSignal(5) => X_Logic0_port, zeroSignal(4) => 
                           X_Logic0_port, zeroSignal(3) => X_Logic0_port, 
                           zeroSignal(2) => X_Logic0_port, zeroSignal(1) => 
                           X_Logic0_port, zeroSignal(0) => X_Logic0_port, 
                           A_signal(63) => positive_inputs_26_63_port, 
                           A_signal(62) => positive_inputs_26_62_port, 
                           A_signal(61) => positive_inputs_26_61_port, 
                           A_signal(60) => positive_inputs_26_60_port, 
                           A_signal(59) => positive_inputs_26_59_port, 
                           A_signal(58) => positive_inputs_26_58_port, 
                           A_signal(57) => positive_inputs_26_57_port, 
                           A_signal(56) => positive_inputs_26_56_port, 
                           A_signal(55) => positive_inputs_26_55_port, 
                           A_signal(54) => positive_inputs_26_54_port, 
                           A_signal(53) => positive_inputs_26_53_port, 
                           A_signal(52) => positive_inputs_26_52_port, 
                           A_signal(51) => positive_inputs_26_51_port, 
                           A_signal(50) => positive_inputs_26_50_port, 
                           A_signal(49) => positive_inputs_26_49_port, 
                           A_signal(48) => positive_inputs_26_48_port, 
                           A_signal(47) => positive_inputs_26_47_port, 
                           A_signal(46) => positive_inputs_26_46_port, 
                           A_signal(45) => positive_inputs_26_45_port, 
                           A_signal(44) => positive_inputs_26_44_port, 
                           A_signal(43) => positive_inputs_26_43_port, 
                           A_signal(42) => positive_inputs_26_42_port, 
                           A_signal(41) => positive_inputs_26_41_port, 
                           A_signal(40) => positive_inputs_26_40_port, 
                           A_signal(39) => positive_inputs_26_39_port, 
                           A_signal(38) => positive_inputs_26_38_port, 
                           A_signal(37) => positive_inputs_26_37_port, 
                           A_signal(36) => positive_inputs_26_36_port, 
                           A_signal(35) => positive_inputs_26_35_port, 
                           A_signal(34) => positive_inputs_26_34_port, 
                           A_signal(33) => positive_inputs_26_33_port, 
                           A_signal(32) => positive_inputs_26_32_port, 
                           A_signal(31) => positive_inputs_26_31_port, 
                           A_signal(30) => positive_inputs_26_30_port, 
                           A_signal(29) => positive_inputs_26_29_port, 
                           A_signal(28) => positive_inputs_26_28_port, 
                           A_signal(27) => positive_inputs_26_27_port, 
                           A_signal(26) => positive_inputs_26_26_port, 
                           A_signal(25) => positive_inputs_26_25_port, 
                           A_signal(24) => positive_inputs_26_24_port, 
                           A_signal(23) => positive_inputs_26_23_port, 
                           A_signal(22) => positive_inputs_26_22_port, 
                           A_signal(21) => positive_inputs_26_21_port, 
                           A_signal(20) => positive_inputs_26_20_port, 
                           A_signal(19) => positive_inputs_26_19_port, 
                           A_signal(18) => positive_inputs_26_18_port, 
                           A_signal(17) => positive_inputs_26_17_port, 
                           A_signal(16) => positive_inputs_26_16_port, 
                           A_signal(15) => positive_inputs_26_15_port, 
                           A_signal(14) => positive_inputs_26_14_port, 
                           A_signal(13) => positive_inputs_26_13_port, 
                           A_signal(12) => positive_inputs_26_12_port, 
                           A_signal(11) => positive_inputs_26_11_port, 
                           A_signal(10) => positive_inputs_26_10_port, 
                           A_signal(9) => positive_inputs_26_9_port, 
                           A_signal(8) => positive_inputs_26_8_port, 
                           A_signal(7) => positive_inputs_26_7_port, 
                           A_signal(6) => positive_inputs_26_6_port, 
                           A_signal(5) => positive_inputs_26_5_port, 
                           A_signal(4) => positive_inputs_26_4_port, 
                           A_signal(3) => positive_inputs_26_3_port, 
                           A_signal(2) => positive_inputs_26_2_port, 
                           A_signal(1) => positive_inputs_26_1_port, 
                           A_signal(0) => n8, A_neg(63) => 
                           negative_inputs_26_63_port, A_neg(62) => 
                           negative_inputs_26_62_port, A_neg(61) => 
                           negative_inputs_26_61_port, A_neg(60) => 
                           negative_inputs_26_60_port, A_neg(59) => 
                           negative_inputs_26_59_port, A_neg(58) => 
                           negative_inputs_26_58_port, A_neg(57) => 
                           negative_inputs_26_57_port, A_neg(56) => 
                           negative_inputs_26_56_port, A_neg(55) => 
                           negative_inputs_26_55_port, A_neg(54) => 
                           negative_inputs_26_54_port, A_neg(53) => 
                           negative_inputs_26_53_port, A_neg(52) => 
                           negative_inputs_26_52_port, A_neg(51) => 
                           negative_inputs_26_51_port, A_neg(50) => 
                           negative_inputs_26_50_port, A_neg(49) => 
                           negative_inputs_26_49_port, A_neg(48) => 
                           negative_inputs_26_48_port, A_neg(47) => 
                           negative_inputs_26_47_port, A_neg(46) => 
                           negative_inputs_26_46_port, A_neg(45) => 
                           negative_inputs_26_45_port, A_neg(44) => 
                           negative_inputs_26_44_port, A_neg(43) => 
                           negative_inputs_26_43_port, A_neg(42) => 
                           negative_inputs_26_42_port, A_neg(41) => 
                           negative_inputs_26_41_port, A_neg(40) => 
                           negative_inputs_26_40_port, A_neg(39) => 
                           negative_inputs_26_39_port, A_neg(38) => 
                           negative_inputs_26_38_port, A_neg(37) => 
                           negative_inputs_26_37_port, A_neg(36) => 
                           negative_inputs_26_36_port, A_neg(35) => 
                           negative_inputs_26_35_port, A_neg(34) => 
                           negative_inputs_26_34_port, A_neg(33) => 
                           negative_inputs_26_33_port, A_neg(32) => 
                           negative_inputs_26_32_port, A_neg(31) => 
                           negative_inputs_26_31_port, A_neg(30) => 
                           negative_inputs_26_30_port, A_neg(29) => 
                           negative_inputs_26_29_port, A_neg(28) => 
                           negative_inputs_26_28_port, A_neg(27) => 
                           negative_inputs_26_27_port, A_neg(26) => 
                           negative_inputs_26_26_port, A_neg(25) => 
                           negative_inputs_26_25_port, A_neg(24) => 
                           negative_inputs_26_24_port, A_neg(23) => 
                           negative_inputs_26_23_port, A_neg(22) => 
                           negative_inputs_26_22_port, A_neg(21) => 
                           negative_inputs_26_21_port, A_neg(20) => 
                           negative_inputs_26_20_port, A_neg(19) => 
                           negative_inputs_26_19_port, A_neg(18) => 
                           negative_inputs_26_18_port, A_neg(17) => 
                           negative_inputs_26_17_port, A_neg(16) => 
                           negative_inputs_26_16_port, A_neg(15) => 
                           negative_inputs_26_15_port, A_neg(14) => 
                           negative_inputs_26_14_port, A_neg(13) => 
                           negative_inputs_26_13_port, A_neg(12) => 
                           negative_inputs_26_12_port, A_neg(11) => 
                           negative_inputs_26_11_port, A_neg(10) => 
                           negative_inputs_26_10_port, A_neg(9) => 
                           negative_inputs_26_9_port, A_neg(8) => 
                           negative_inputs_26_8_port, A_neg(7) => 
                           negative_inputs_26_7_port, A_neg(6) => 
                           negative_inputs_26_6_port, A_neg(5) => 
                           negative_inputs_26_5_port, A_neg(4) => 
                           negative_inputs_26_4_port, A_neg(3) => 
                           negative_inputs_26_3_port, A_neg(2) => 
                           negative_inputs_26_2_port, A_neg(1) => 
                           negative_inputs_26_1_port, A_neg(0) => n8, 
                           A_shifted(63) => positive_inputs_27_63_port, 
                           A_shifted(62) => positive_inputs_27_62_port, 
                           A_shifted(61) => positive_inputs_27_61_port, 
                           A_shifted(60) => positive_inputs_27_60_port, 
                           A_shifted(59) => positive_inputs_27_59_port, 
                           A_shifted(58) => positive_inputs_27_58_port, 
                           A_shifted(57) => positive_inputs_27_57_port, 
                           A_shifted(56) => positive_inputs_27_56_port, 
                           A_shifted(55) => positive_inputs_27_55_port, 
                           A_shifted(54) => positive_inputs_27_54_port, 
                           A_shifted(53) => positive_inputs_27_53_port, 
                           A_shifted(52) => positive_inputs_27_52_port, 
                           A_shifted(51) => positive_inputs_27_51_port, 
                           A_shifted(50) => positive_inputs_27_50_port, 
                           A_shifted(49) => positive_inputs_27_49_port, 
                           A_shifted(48) => positive_inputs_27_48_port, 
                           A_shifted(47) => positive_inputs_27_47_port, 
                           A_shifted(46) => positive_inputs_27_46_port, 
                           A_shifted(45) => positive_inputs_27_45_port, 
                           A_shifted(44) => positive_inputs_27_44_port, 
                           A_shifted(43) => positive_inputs_27_43_port, 
                           A_shifted(42) => positive_inputs_27_42_port, 
                           A_shifted(41) => positive_inputs_27_41_port, 
                           A_shifted(40) => positive_inputs_27_40_port, 
                           A_shifted(39) => positive_inputs_27_39_port, 
                           A_shifted(38) => positive_inputs_27_38_port, 
                           A_shifted(37) => positive_inputs_27_37_port, 
                           A_shifted(36) => positive_inputs_27_36_port, 
                           A_shifted(35) => positive_inputs_27_35_port, 
                           A_shifted(34) => positive_inputs_27_34_port, 
                           A_shifted(33) => positive_inputs_27_33_port, 
                           A_shifted(32) => positive_inputs_27_32_port, 
                           A_shifted(31) => positive_inputs_27_31_port, 
                           A_shifted(30) => positive_inputs_27_30_port, 
                           A_shifted(29) => positive_inputs_27_29_port, 
                           A_shifted(28) => positive_inputs_27_28_port, 
                           A_shifted(27) => positive_inputs_27_27_port, 
                           A_shifted(26) => positive_inputs_27_26_port, 
                           A_shifted(25) => positive_inputs_27_25_port, 
                           A_shifted(24) => positive_inputs_27_24_port, 
                           A_shifted(23) => positive_inputs_27_23_port, 
                           A_shifted(22) => positive_inputs_27_22_port, 
                           A_shifted(21) => positive_inputs_27_21_port, 
                           A_shifted(20) => positive_inputs_27_20_port, 
                           A_shifted(19) => positive_inputs_27_19_port, 
                           A_shifted(18) => positive_inputs_27_18_port, 
                           A_shifted(17) => positive_inputs_27_17_port, 
                           A_shifted(16) => positive_inputs_27_16_port, 
                           A_shifted(15) => positive_inputs_27_15_port, 
                           A_shifted(14) => positive_inputs_27_14_port, 
                           A_shifted(13) => positive_inputs_27_13_port, 
                           A_shifted(12) => positive_inputs_27_12_port, 
                           A_shifted(11) => positive_inputs_27_11_port, 
                           A_shifted(10) => positive_inputs_27_10_port, 
                           A_shifted(9) => positive_inputs_27_9_port, 
                           A_shifted(8) => positive_inputs_27_8_port, 
                           A_shifted(7) => positive_inputs_27_7_port, 
                           A_shifted(6) => positive_inputs_27_6_port, 
                           A_shifted(5) => positive_inputs_27_5_port, 
                           A_shifted(4) => positive_inputs_27_4_port, 
                           A_shifted(3) => positive_inputs_27_3_port, 
                           A_shifted(2) => positive_inputs_27_2_port, 
                           A_shifted(1) => positive_inputs_27_1_port, 
                           A_shifted(0) => n8, A_neg_shifted(63) => 
                           negative_inputs_27_63_port, A_neg_shifted(62) => 
                           negative_inputs_27_62_port, A_neg_shifted(61) => 
                           negative_inputs_27_61_port, A_neg_shifted(60) => 
                           negative_inputs_27_60_port, A_neg_shifted(59) => 
                           negative_inputs_27_59_port, A_neg_shifted(58) => 
                           negative_inputs_27_58_port, A_neg_shifted(57) => 
                           negative_inputs_27_57_port, A_neg_shifted(56) => 
                           negative_inputs_27_56_port, A_neg_shifted(55) => 
                           negative_inputs_27_55_port, A_neg_shifted(54) => 
                           negative_inputs_27_54_port, A_neg_shifted(53) => 
                           negative_inputs_27_53_port, A_neg_shifted(52) => 
                           negative_inputs_27_52_port, A_neg_shifted(51) => 
                           negative_inputs_27_51_port, A_neg_shifted(50) => 
                           negative_inputs_27_50_port, A_neg_shifted(49) => 
                           negative_inputs_27_49_port, A_neg_shifted(48) => 
                           negative_inputs_27_48_port, A_neg_shifted(47) => 
                           negative_inputs_27_47_port, A_neg_shifted(46) => 
                           negative_inputs_27_46_port, A_neg_shifted(45) => 
                           negative_inputs_27_45_port, A_neg_shifted(44) => 
                           negative_inputs_27_44_port, A_neg_shifted(43) => 
                           negative_inputs_27_43_port, A_neg_shifted(42) => 
                           negative_inputs_27_42_port, A_neg_shifted(41) => 
                           negative_inputs_27_41_port, A_neg_shifted(40) => 
                           negative_inputs_27_40_port, A_neg_shifted(39) => 
                           negative_inputs_27_39_port, A_neg_shifted(38) => 
                           negative_inputs_27_38_port, A_neg_shifted(37) => 
                           negative_inputs_27_37_port, A_neg_shifted(36) => 
                           negative_inputs_27_36_port, A_neg_shifted(35) => 
                           negative_inputs_27_35_port, A_neg_shifted(34) => 
                           negative_inputs_27_34_port, A_neg_shifted(33) => 
                           negative_inputs_27_33_port, A_neg_shifted(32) => 
                           negative_inputs_27_32_port, A_neg_shifted(31) => 
                           negative_inputs_27_31_port, A_neg_shifted(30) => 
                           negative_inputs_27_30_port, A_neg_shifted(29) => 
                           negative_inputs_27_29_port, A_neg_shifted(28) => 
                           negative_inputs_27_28_port, A_neg_shifted(27) => 
                           negative_inputs_27_27_port, A_neg_shifted(26) => 
                           negative_inputs_27_26_port, A_neg_shifted(25) => 
                           negative_inputs_27_25_port, A_neg_shifted(24) => 
                           negative_inputs_27_24_port, A_neg_shifted(23) => 
                           negative_inputs_27_23_port, A_neg_shifted(22) => 
                           negative_inputs_27_22_port, A_neg_shifted(21) => 
                           negative_inputs_27_21_port, A_neg_shifted(20) => 
                           negative_inputs_27_20_port, A_neg_shifted(19) => 
                           negative_inputs_27_19_port, A_neg_shifted(18) => 
                           negative_inputs_27_18_port, A_neg_shifted(17) => 
                           negative_inputs_27_17_port, A_neg_shifted(16) => 
                           negative_inputs_27_16_port, A_neg_shifted(15) => 
                           negative_inputs_27_15_port, A_neg_shifted(14) => 
                           negative_inputs_27_14_port, A_neg_shifted(13) => 
                           negative_inputs_27_13_port, A_neg_shifted(12) => 
                           negative_inputs_27_12_port, A_neg_shifted(11) => 
                           negative_inputs_27_11_port, A_neg_shifted(10) => 
                           negative_inputs_27_10_port, A_neg_shifted(9) => 
                           negative_inputs_27_9_port, A_neg_shifted(8) => 
                           negative_inputs_27_8_port, A_neg_shifted(7) => 
                           negative_inputs_27_7_port, A_neg_shifted(6) => 
                           negative_inputs_27_6_port, A_neg_shifted(5) => 
                           negative_inputs_27_5_port, A_neg_shifted(4) => 
                           negative_inputs_27_4_port, A_neg_shifted(3) => 
                           negative_inputs_27_3_port, A_neg_shifted(2) => 
                           negative_inputs_27_2_port, A_neg_shifted(1) => 
                           negative_inputs_27_1_port, A_neg_shifted(0) => n8, 
                           Sel(2) => sel_13_2_port, Sel(1) => sel_13_1_port, 
                           Sel(0) => sel_13_0_port, Y(63) => 
                           MuxOutputs_13_63_port, Y(62) => 
                           MuxOutputs_13_62_port, Y(61) => 
                           MuxOutputs_13_61_port, Y(60) => 
                           MuxOutputs_13_60_port, Y(59) => 
                           MuxOutputs_13_59_port, Y(58) => 
                           MuxOutputs_13_58_port, Y(57) => 
                           MuxOutputs_13_57_port, Y(56) => 
                           MuxOutputs_13_56_port, Y(55) => 
                           MuxOutputs_13_55_port, Y(54) => 
                           MuxOutputs_13_54_port, Y(53) => 
                           MuxOutputs_13_53_port, Y(52) => 
                           MuxOutputs_13_52_port, Y(51) => 
                           MuxOutputs_13_51_port, Y(50) => 
                           MuxOutputs_13_50_port, Y(49) => 
                           MuxOutputs_13_49_port, Y(48) => 
                           MuxOutputs_13_48_port, Y(47) => 
                           MuxOutputs_13_47_port, Y(46) => 
                           MuxOutputs_13_46_port, Y(45) => 
                           MuxOutputs_13_45_port, Y(44) => 
                           MuxOutputs_13_44_port, Y(43) => 
                           MuxOutputs_13_43_port, Y(42) => 
                           MuxOutputs_13_42_port, Y(41) => 
                           MuxOutputs_13_41_port, Y(40) => 
                           MuxOutputs_13_40_port, Y(39) => 
                           MuxOutputs_13_39_port, Y(38) => 
                           MuxOutputs_13_38_port, Y(37) => 
                           MuxOutputs_13_37_port, Y(36) => 
                           MuxOutputs_13_36_port, Y(35) => 
                           MuxOutputs_13_35_port, Y(34) => 
                           MuxOutputs_13_34_port, Y(33) => 
                           MuxOutputs_13_33_port, Y(32) => 
                           MuxOutputs_13_32_port, Y(31) => 
                           MuxOutputs_13_31_port, Y(30) => 
                           MuxOutputs_13_30_port, Y(29) => 
                           MuxOutputs_13_29_port, Y(28) => 
                           MuxOutputs_13_28_port, Y(27) => 
                           MuxOutputs_13_27_port, Y(26) => 
                           MuxOutputs_13_26_port, Y(25) => 
                           MuxOutputs_13_25_port, Y(24) => 
                           MuxOutputs_13_24_port, Y(23) => 
                           MuxOutputs_13_23_port, Y(22) => 
                           MuxOutputs_13_22_port, Y(21) => 
                           MuxOutputs_13_21_port, Y(20) => 
                           MuxOutputs_13_20_port, Y(19) => 
                           MuxOutputs_13_19_port, Y(18) => 
                           MuxOutputs_13_18_port, Y(17) => 
                           MuxOutputs_13_17_port, Y(16) => 
                           MuxOutputs_13_16_port, Y(15) => 
                           MuxOutputs_13_15_port, Y(14) => 
                           MuxOutputs_13_14_port, Y(13) => 
                           MuxOutputs_13_13_port, Y(12) => 
                           MuxOutputs_13_12_port, Y(11) => 
                           MuxOutputs_13_11_port, Y(10) => 
                           MuxOutputs_13_10_port, Y(9) => MuxOutputs_13_9_port,
                           Y(8) => MuxOutputs_13_8_port, Y(7) => 
                           MuxOutputs_13_7_port, Y(6) => MuxOutputs_13_6_port, 
                           Y(5) => MuxOutputs_13_5_port, Y(4) => 
                           MuxOutputs_13_4_port, Y(3) => MuxOutputs_13_3_port, 
                           Y(2) => MuxOutputs_13_2_port, Y(1) => 
                           MuxOutputs_13_1_port, Y(0) => MuxOutputs_13_0_port);
   encoderI_14 : encoder_18 port map( pieceofB(2) => B(29), pieceofB(1) => 
                           B(28), pieceofB(0) => B(27), sel(2) => sel_14_2_port
                           , sel(1) => sel_14_1_port, sel(0) => sel_14_0_port);
   MUXI_14 : MUX51_MuxNbit64_18 port map( zeroSignal(63) => X_Logic0_port, 
                           zeroSignal(62) => X_Logic0_port, zeroSignal(61) => 
                           X_Logic0_port, zeroSignal(60) => X_Logic0_port, 
                           zeroSignal(59) => X_Logic0_port, zeroSignal(58) => 
                           X_Logic0_port, zeroSignal(57) => X_Logic0_port, 
                           zeroSignal(56) => X_Logic0_port, zeroSignal(55) => 
                           X_Logic0_port, zeroSignal(54) => X_Logic0_port, 
                           zeroSignal(53) => X_Logic0_port, zeroSignal(52) => 
                           X_Logic0_port, zeroSignal(51) => X_Logic0_port, 
                           zeroSignal(50) => X_Logic0_port, zeroSignal(49) => 
                           X_Logic0_port, zeroSignal(48) => X_Logic0_port, 
                           zeroSignal(47) => X_Logic0_port, zeroSignal(46) => 
                           X_Logic0_port, zeroSignal(45) => X_Logic0_port, 
                           zeroSignal(44) => X_Logic0_port, zeroSignal(43) => 
                           X_Logic0_port, zeroSignal(42) => X_Logic0_port, 
                           zeroSignal(41) => X_Logic0_port, zeroSignal(40) => 
                           X_Logic0_port, zeroSignal(39) => X_Logic0_port, 
                           zeroSignal(38) => X_Logic0_port, zeroSignal(37) => 
                           X_Logic0_port, zeroSignal(36) => X_Logic0_port, 
                           zeroSignal(35) => X_Logic0_port, zeroSignal(34) => 
                           X_Logic0_port, zeroSignal(33) => X_Logic0_port, 
                           zeroSignal(32) => X_Logic0_port, zeroSignal(31) => 
                           X_Logic0_port, zeroSignal(30) => X_Logic0_port, 
                           zeroSignal(29) => X_Logic0_port, zeroSignal(28) => 
                           X_Logic0_port, zeroSignal(27) => X_Logic0_port, 
                           zeroSignal(26) => X_Logic0_port, zeroSignal(25) => 
                           X_Logic0_port, zeroSignal(24) => X_Logic0_port, 
                           zeroSignal(23) => X_Logic0_port, zeroSignal(22) => 
                           X_Logic0_port, zeroSignal(21) => X_Logic0_port, 
                           zeroSignal(20) => X_Logic0_port, zeroSignal(19) => 
                           X_Logic0_port, zeroSignal(18) => X_Logic0_port, 
                           zeroSignal(17) => X_Logic0_port, zeroSignal(16) => 
                           X_Logic0_port, zeroSignal(15) => X_Logic0_port, 
                           zeroSignal(14) => X_Logic0_port, zeroSignal(13) => 
                           X_Logic0_port, zeroSignal(12) => X_Logic0_port, 
                           zeroSignal(11) => X_Logic0_port, zeroSignal(10) => 
                           X_Logic0_port, zeroSignal(9) => X_Logic0_port, 
                           zeroSignal(8) => X_Logic0_port, zeroSignal(7) => 
                           X_Logic0_port, zeroSignal(6) => X_Logic0_port, 
                           zeroSignal(5) => X_Logic0_port, zeroSignal(4) => 
                           X_Logic0_port, zeroSignal(3) => X_Logic0_port, 
                           zeroSignal(2) => X_Logic0_port, zeroSignal(1) => 
                           X_Logic0_port, zeroSignal(0) => X_Logic0_port, 
                           A_signal(63) => positive_inputs_28_63_port, 
                           A_signal(62) => positive_inputs_28_62_port, 
                           A_signal(61) => positive_inputs_28_61_port, 
                           A_signal(60) => positive_inputs_28_60_port, 
                           A_signal(59) => positive_inputs_28_59_port, 
                           A_signal(58) => positive_inputs_28_58_port, 
                           A_signal(57) => positive_inputs_28_57_port, 
                           A_signal(56) => positive_inputs_28_56_port, 
                           A_signal(55) => positive_inputs_28_55_port, 
                           A_signal(54) => positive_inputs_28_54_port, 
                           A_signal(53) => positive_inputs_28_53_port, 
                           A_signal(52) => positive_inputs_28_52_port, 
                           A_signal(51) => positive_inputs_28_51_port, 
                           A_signal(50) => positive_inputs_28_50_port, 
                           A_signal(49) => positive_inputs_28_49_port, 
                           A_signal(48) => positive_inputs_28_48_port, 
                           A_signal(47) => positive_inputs_28_47_port, 
                           A_signal(46) => positive_inputs_28_46_port, 
                           A_signal(45) => positive_inputs_28_45_port, 
                           A_signal(44) => positive_inputs_28_44_port, 
                           A_signal(43) => positive_inputs_28_43_port, 
                           A_signal(42) => positive_inputs_28_42_port, 
                           A_signal(41) => positive_inputs_28_41_port, 
                           A_signal(40) => positive_inputs_28_40_port, 
                           A_signal(39) => positive_inputs_28_39_port, 
                           A_signal(38) => positive_inputs_28_38_port, 
                           A_signal(37) => positive_inputs_28_37_port, 
                           A_signal(36) => positive_inputs_28_36_port, 
                           A_signal(35) => positive_inputs_28_35_port, 
                           A_signal(34) => positive_inputs_28_34_port, 
                           A_signal(33) => positive_inputs_28_33_port, 
                           A_signal(32) => positive_inputs_28_32_port, 
                           A_signal(31) => positive_inputs_28_31_port, 
                           A_signal(30) => positive_inputs_28_30_port, 
                           A_signal(29) => positive_inputs_28_29_port, 
                           A_signal(28) => positive_inputs_28_28_port, 
                           A_signal(27) => positive_inputs_28_27_port, 
                           A_signal(26) => positive_inputs_28_26_port, 
                           A_signal(25) => positive_inputs_28_25_port, 
                           A_signal(24) => positive_inputs_28_24_port, 
                           A_signal(23) => positive_inputs_28_23_port, 
                           A_signal(22) => positive_inputs_28_22_port, 
                           A_signal(21) => positive_inputs_28_21_port, 
                           A_signal(20) => positive_inputs_28_20_port, 
                           A_signal(19) => positive_inputs_28_19_port, 
                           A_signal(18) => positive_inputs_28_18_port, 
                           A_signal(17) => positive_inputs_28_17_port, 
                           A_signal(16) => positive_inputs_28_16_port, 
                           A_signal(15) => positive_inputs_28_15_port, 
                           A_signal(14) => positive_inputs_28_14_port, 
                           A_signal(13) => positive_inputs_28_13_port, 
                           A_signal(12) => positive_inputs_28_12_port, 
                           A_signal(11) => positive_inputs_28_11_port, 
                           A_signal(10) => positive_inputs_28_10_port, 
                           A_signal(9) => positive_inputs_28_9_port, 
                           A_signal(8) => positive_inputs_28_8_port, 
                           A_signal(7) => positive_inputs_28_7_port, 
                           A_signal(6) => positive_inputs_28_6_port, 
                           A_signal(5) => positive_inputs_28_5_port, 
                           A_signal(4) => positive_inputs_28_4_port, 
                           A_signal(3) => positive_inputs_28_3_port, 
                           A_signal(2) => positive_inputs_28_2_port, 
                           A_signal(1) => positive_inputs_28_1_port, 
                           A_signal(0) => n8, A_neg(63) => 
                           negative_inputs_28_63_port, A_neg(62) => 
                           negative_inputs_28_62_port, A_neg(61) => 
                           negative_inputs_28_61_port, A_neg(60) => 
                           negative_inputs_28_60_port, A_neg(59) => 
                           negative_inputs_28_59_port, A_neg(58) => 
                           negative_inputs_28_58_port, A_neg(57) => 
                           negative_inputs_28_57_port, A_neg(56) => 
                           negative_inputs_28_56_port, A_neg(55) => 
                           negative_inputs_28_55_port, A_neg(54) => 
                           negative_inputs_28_54_port, A_neg(53) => 
                           negative_inputs_28_53_port, A_neg(52) => 
                           negative_inputs_28_52_port, A_neg(51) => 
                           negative_inputs_28_51_port, A_neg(50) => 
                           negative_inputs_28_50_port, A_neg(49) => 
                           negative_inputs_28_49_port, A_neg(48) => 
                           negative_inputs_28_48_port, A_neg(47) => 
                           negative_inputs_28_47_port, A_neg(46) => 
                           negative_inputs_28_46_port, A_neg(45) => 
                           negative_inputs_28_45_port, A_neg(44) => 
                           negative_inputs_28_44_port, A_neg(43) => 
                           negative_inputs_28_43_port, A_neg(42) => 
                           negative_inputs_28_42_port, A_neg(41) => 
                           negative_inputs_28_41_port, A_neg(40) => 
                           negative_inputs_28_40_port, A_neg(39) => 
                           negative_inputs_28_39_port, A_neg(38) => 
                           negative_inputs_28_38_port, A_neg(37) => 
                           negative_inputs_28_37_port, A_neg(36) => 
                           negative_inputs_28_36_port, A_neg(35) => 
                           negative_inputs_28_35_port, A_neg(34) => 
                           negative_inputs_28_34_port, A_neg(33) => 
                           negative_inputs_28_33_port, A_neg(32) => 
                           negative_inputs_28_32_port, A_neg(31) => 
                           negative_inputs_28_31_port, A_neg(30) => 
                           negative_inputs_28_30_port, A_neg(29) => 
                           negative_inputs_28_29_port, A_neg(28) => 
                           negative_inputs_28_28_port, A_neg(27) => 
                           negative_inputs_28_27_port, A_neg(26) => 
                           negative_inputs_28_26_port, A_neg(25) => 
                           negative_inputs_28_25_port, A_neg(24) => 
                           negative_inputs_28_24_port, A_neg(23) => 
                           negative_inputs_28_23_port, A_neg(22) => 
                           negative_inputs_28_22_port, A_neg(21) => 
                           negative_inputs_28_21_port, A_neg(20) => 
                           negative_inputs_28_20_port, A_neg(19) => 
                           negative_inputs_28_19_port, A_neg(18) => 
                           negative_inputs_28_18_port, A_neg(17) => 
                           negative_inputs_28_17_port, A_neg(16) => 
                           negative_inputs_28_16_port, A_neg(15) => 
                           negative_inputs_28_15_port, A_neg(14) => 
                           negative_inputs_28_14_port, A_neg(13) => 
                           negative_inputs_28_13_port, A_neg(12) => 
                           negative_inputs_28_12_port, A_neg(11) => 
                           negative_inputs_28_11_port, A_neg(10) => 
                           negative_inputs_28_10_port, A_neg(9) => 
                           negative_inputs_28_9_port, A_neg(8) => 
                           negative_inputs_28_8_port, A_neg(7) => 
                           negative_inputs_28_7_port, A_neg(6) => 
                           negative_inputs_28_6_port, A_neg(5) => 
                           negative_inputs_28_5_port, A_neg(4) => 
                           negative_inputs_28_4_port, A_neg(3) => 
                           negative_inputs_28_3_port, A_neg(2) => 
                           negative_inputs_28_2_port, A_neg(1) => 
                           negative_inputs_28_1_port, A_neg(0) => n8, 
                           A_shifted(63) => positive_inputs_29_63_port, 
                           A_shifted(62) => positive_inputs_29_62_port, 
                           A_shifted(61) => positive_inputs_29_61_port, 
                           A_shifted(60) => positive_inputs_29_60_port, 
                           A_shifted(59) => positive_inputs_29_59_port, 
                           A_shifted(58) => positive_inputs_29_58_port, 
                           A_shifted(57) => positive_inputs_29_57_port, 
                           A_shifted(56) => positive_inputs_29_56_port, 
                           A_shifted(55) => positive_inputs_29_55_port, 
                           A_shifted(54) => positive_inputs_29_54_port, 
                           A_shifted(53) => positive_inputs_29_53_port, 
                           A_shifted(52) => positive_inputs_29_52_port, 
                           A_shifted(51) => positive_inputs_29_51_port, 
                           A_shifted(50) => positive_inputs_29_50_port, 
                           A_shifted(49) => positive_inputs_29_49_port, 
                           A_shifted(48) => positive_inputs_29_48_port, 
                           A_shifted(47) => positive_inputs_29_47_port, 
                           A_shifted(46) => positive_inputs_29_46_port, 
                           A_shifted(45) => positive_inputs_29_45_port, 
                           A_shifted(44) => positive_inputs_29_44_port, 
                           A_shifted(43) => positive_inputs_29_43_port, 
                           A_shifted(42) => positive_inputs_29_42_port, 
                           A_shifted(41) => positive_inputs_29_41_port, 
                           A_shifted(40) => positive_inputs_29_40_port, 
                           A_shifted(39) => positive_inputs_29_39_port, 
                           A_shifted(38) => positive_inputs_29_38_port, 
                           A_shifted(37) => positive_inputs_29_37_port, 
                           A_shifted(36) => positive_inputs_29_36_port, 
                           A_shifted(35) => positive_inputs_29_35_port, 
                           A_shifted(34) => positive_inputs_29_34_port, 
                           A_shifted(33) => positive_inputs_29_33_port, 
                           A_shifted(32) => positive_inputs_29_32_port, 
                           A_shifted(31) => positive_inputs_29_31_port, 
                           A_shifted(30) => positive_inputs_29_30_port, 
                           A_shifted(29) => positive_inputs_29_29_port, 
                           A_shifted(28) => positive_inputs_29_28_port, 
                           A_shifted(27) => positive_inputs_29_27_port, 
                           A_shifted(26) => positive_inputs_29_26_port, 
                           A_shifted(25) => positive_inputs_29_25_port, 
                           A_shifted(24) => positive_inputs_29_24_port, 
                           A_shifted(23) => positive_inputs_29_23_port, 
                           A_shifted(22) => positive_inputs_29_22_port, 
                           A_shifted(21) => positive_inputs_29_21_port, 
                           A_shifted(20) => positive_inputs_29_20_port, 
                           A_shifted(19) => positive_inputs_29_19_port, 
                           A_shifted(18) => positive_inputs_29_18_port, 
                           A_shifted(17) => positive_inputs_29_17_port, 
                           A_shifted(16) => positive_inputs_29_16_port, 
                           A_shifted(15) => positive_inputs_29_15_port, 
                           A_shifted(14) => positive_inputs_29_14_port, 
                           A_shifted(13) => positive_inputs_29_13_port, 
                           A_shifted(12) => positive_inputs_29_12_port, 
                           A_shifted(11) => positive_inputs_29_11_port, 
                           A_shifted(10) => positive_inputs_29_10_port, 
                           A_shifted(9) => positive_inputs_29_9_port, 
                           A_shifted(8) => positive_inputs_29_8_port, 
                           A_shifted(7) => positive_inputs_29_7_port, 
                           A_shifted(6) => positive_inputs_29_6_port, 
                           A_shifted(5) => positive_inputs_29_5_port, 
                           A_shifted(4) => positive_inputs_29_4_port, 
                           A_shifted(3) => positive_inputs_29_3_port, 
                           A_shifted(2) => positive_inputs_29_2_port, 
                           A_shifted(1) => positive_inputs_29_1_port, 
                           A_shifted(0) => n8, A_neg_shifted(63) => 
                           negative_inputs_29_63_port, A_neg_shifted(62) => 
                           negative_inputs_29_62_port, A_neg_shifted(61) => 
                           negative_inputs_29_61_port, A_neg_shifted(60) => 
                           negative_inputs_29_60_port, A_neg_shifted(59) => 
                           negative_inputs_29_59_port, A_neg_shifted(58) => 
                           negative_inputs_29_58_port, A_neg_shifted(57) => 
                           negative_inputs_29_57_port, A_neg_shifted(56) => 
                           negative_inputs_29_56_port, A_neg_shifted(55) => 
                           negative_inputs_29_55_port, A_neg_shifted(54) => 
                           negative_inputs_29_54_port, A_neg_shifted(53) => 
                           negative_inputs_29_53_port, A_neg_shifted(52) => 
                           negative_inputs_29_52_port, A_neg_shifted(51) => 
                           negative_inputs_29_51_port, A_neg_shifted(50) => 
                           negative_inputs_29_50_port, A_neg_shifted(49) => 
                           negative_inputs_29_49_port, A_neg_shifted(48) => 
                           negative_inputs_29_48_port, A_neg_shifted(47) => 
                           negative_inputs_29_47_port, A_neg_shifted(46) => 
                           negative_inputs_29_46_port, A_neg_shifted(45) => 
                           negative_inputs_29_45_port, A_neg_shifted(44) => 
                           negative_inputs_29_44_port, A_neg_shifted(43) => 
                           negative_inputs_29_43_port, A_neg_shifted(42) => 
                           negative_inputs_29_42_port, A_neg_shifted(41) => 
                           negative_inputs_29_41_port, A_neg_shifted(40) => 
                           negative_inputs_29_40_port, A_neg_shifted(39) => 
                           negative_inputs_29_39_port, A_neg_shifted(38) => 
                           negative_inputs_29_38_port, A_neg_shifted(37) => 
                           negative_inputs_29_37_port, A_neg_shifted(36) => 
                           negative_inputs_29_36_port, A_neg_shifted(35) => 
                           negative_inputs_29_35_port, A_neg_shifted(34) => 
                           negative_inputs_29_34_port, A_neg_shifted(33) => 
                           negative_inputs_29_33_port, A_neg_shifted(32) => 
                           negative_inputs_29_32_port, A_neg_shifted(31) => 
                           negative_inputs_29_31_port, A_neg_shifted(30) => 
                           negative_inputs_29_30_port, A_neg_shifted(29) => 
                           negative_inputs_29_29_port, A_neg_shifted(28) => 
                           negative_inputs_29_28_port, A_neg_shifted(27) => 
                           negative_inputs_29_27_port, A_neg_shifted(26) => 
                           negative_inputs_29_26_port, A_neg_shifted(25) => 
                           negative_inputs_29_25_port, A_neg_shifted(24) => 
                           negative_inputs_29_24_port, A_neg_shifted(23) => 
                           negative_inputs_29_23_port, A_neg_shifted(22) => 
                           negative_inputs_29_22_port, A_neg_shifted(21) => 
                           negative_inputs_29_21_port, A_neg_shifted(20) => 
                           negative_inputs_29_20_port, A_neg_shifted(19) => 
                           negative_inputs_29_19_port, A_neg_shifted(18) => 
                           negative_inputs_29_18_port, A_neg_shifted(17) => 
                           negative_inputs_29_17_port, A_neg_shifted(16) => 
                           negative_inputs_29_16_port, A_neg_shifted(15) => 
                           negative_inputs_29_15_port, A_neg_shifted(14) => 
                           negative_inputs_29_14_port, A_neg_shifted(13) => 
                           negative_inputs_29_13_port, A_neg_shifted(12) => 
                           negative_inputs_29_12_port, A_neg_shifted(11) => 
                           negative_inputs_29_11_port, A_neg_shifted(10) => 
                           negative_inputs_29_10_port, A_neg_shifted(9) => 
                           negative_inputs_29_9_port, A_neg_shifted(8) => 
                           negative_inputs_29_8_port, A_neg_shifted(7) => 
                           negative_inputs_29_7_port, A_neg_shifted(6) => 
                           negative_inputs_29_6_port, A_neg_shifted(5) => 
                           negative_inputs_29_5_port, A_neg_shifted(4) => 
                           negative_inputs_29_4_port, A_neg_shifted(3) => 
                           negative_inputs_29_3_port, A_neg_shifted(2) => 
                           negative_inputs_29_2_port, A_neg_shifted(1) => 
                           negative_inputs_29_1_port, A_neg_shifted(0) => n8, 
                           Sel(2) => sel_14_2_port, Sel(1) => sel_14_1_port, 
                           Sel(0) => sel_14_0_port, Y(63) => 
                           MuxOutputs_14_63_port, Y(62) => 
                           MuxOutputs_14_62_port, Y(61) => 
                           MuxOutputs_14_61_port, Y(60) => 
                           MuxOutputs_14_60_port, Y(59) => 
                           MuxOutputs_14_59_port, Y(58) => 
                           MuxOutputs_14_58_port, Y(57) => 
                           MuxOutputs_14_57_port, Y(56) => 
                           MuxOutputs_14_56_port, Y(55) => 
                           MuxOutputs_14_55_port, Y(54) => 
                           MuxOutputs_14_54_port, Y(53) => 
                           MuxOutputs_14_53_port, Y(52) => 
                           MuxOutputs_14_52_port, Y(51) => 
                           MuxOutputs_14_51_port, Y(50) => 
                           MuxOutputs_14_50_port, Y(49) => 
                           MuxOutputs_14_49_port, Y(48) => 
                           MuxOutputs_14_48_port, Y(47) => 
                           MuxOutputs_14_47_port, Y(46) => 
                           MuxOutputs_14_46_port, Y(45) => 
                           MuxOutputs_14_45_port, Y(44) => 
                           MuxOutputs_14_44_port, Y(43) => 
                           MuxOutputs_14_43_port, Y(42) => 
                           MuxOutputs_14_42_port, Y(41) => 
                           MuxOutputs_14_41_port, Y(40) => 
                           MuxOutputs_14_40_port, Y(39) => 
                           MuxOutputs_14_39_port, Y(38) => 
                           MuxOutputs_14_38_port, Y(37) => 
                           MuxOutputs_14_37_port, Y(36) => 
                           MuxOutputs_14_36_port, Y(35) => 
                           MuxOutputs_14_35_port, Y(34) => 
                           MuxOutputs_14_34_port, Y(33) => 
                           MuxOutputs_14_33_port, Y(32) => 
                           MuxOutputs_14_32_port, Y(31) => 
                           MuxOutputs_14_31_port, Y(30) => 
                           MuxOutputs_14_30_port, Y(29) => 
                           MuxOutputs_14_29_port, Y(28) => 
                           MuxOutputs_14_28_port, Y(27) => 
                           MuxOutputs_14_27_port, Y(26) => 
                           MuxOutputs_14_26_port, Y(25) => 
                           MuxOutputs_14_25_port, Y(24) => 
                           MuxOutputs_14_24_port, Y(23) => 
                           MuxOutputs_14_23_port, Y(22) => 
                           MuxOutputs_14_22_port, Y(21) => 
                           MuxOutputs_14_21_port, Y(20) => 
                           MuxOutputs_14_20_port, Y(19) => 
                           MuxOutputs_14_19_port, Y(18) => 
                           MuxOutputs_14_18_port, Y(17) => 
                           MuxOutputs_14_17_port, Y(16) => 
                           MuxOutputs_14_16_port, Y(15) => 
                           MuxOutputs_14_15_port, Y(14) => 
                           MuxOutputs_14_14_port, Y(13) => 
                           MuxOutputs_14_13_port, Y(12) => 
                           MuxOutputs_14_12_port, Y(11) => 
                           MuxOutputs_14_11_port, Y(10) => 
                           MuxOutputs_14_10_port, Y(9) => MuxOutputs_14_9_port,
                           Y(8) => MuxOutputs_14_8_port, Y(7) => 
                           MuxOutputs_14_7_port, Y(6) => MuxOutputs_14_6_port, 
                           Y(5) => MuxOutputs_14_5_port, Y(4) => 
                           MuxOutputs_14_4_port, Y(3) => MuxOutputs_14_3_port, 
                           Y(2) => MuxOutputs_14_2_port, Y(1) => 
                           MuxOutputs_14_1_port, Y(0) => MuxOutputs_14_0_port);
   encoderI_15 : encoder_17 port map( pieceofB(2) => B(31), pieceofB(1) => 
                           B(30), pieceofB(0) => B(29), sel(2) => sel_15_2_port
                           , sel(1) => sel_15_1_port, sel(0) => sel_15_0_port);
   MUXI_15 : MUX51_MuxNbit64_17 port map( zeroSignal(63) => X_Logic0_port, 
                           zeroSignal(62) => X_Logic0_port, zeroSignal(61) => 
                           X_Logic0_port, zeroSignal(60) => X_Logic0_port, 
                           zeroSignal(59) => X_Logic0_port, zeroSignal(58) => 
                           X_Logic0_port, zeroSignal(57) => X_Logic0_port, 
                           zeroSignal(56) => X_Logic0_port, zeroSignal(55) => 
                           X_Logic0_port, zeroSignal(54) => X_Logic0_port, 
                           zeroSignal(53) => X_Logic0_port, zeroSignal(52) => 
                           X_Logic0_port, zeroSignal(51) => X_Logic0_port, 
                           zeroSignal(50) => X_Logic0_port, zeroSignal(49) => 
                           X_Logic0_port, zeroSignal(48) => X_Logic0_port, 
                           zeroSignal(47) => X_Logic0_port, zeroSignal(46) => 
                           X_Logic0_port, zeroSignal(45) => X_Logic0_port, 
                           zeroSignal(44) => X_Logic0_port, zeroSignal(43) => 
                           X_Logic0_port, zeroSignal(42) => X_Logic0_port, 
                           zeroSignal(41) => X_Logic0_port, zeroSignal(40) => 
                           X_Logic0_port, zeroSignal(39) => X_Logic0_port, 
                           zeroSignal(38) => X_Logic0_port, zeroSignal(37) => 
                           X_Logic0_port, zeroSignal(36) => X_Logic0_port, 
                           zeroSignal(35) => X_Logic0_port, zeroSignal(34) => 
                           X_Logic0_port, zeroSignal(33) => X_Logic0_port, 
                           zeroSignal(32) => X_Logic0_port, zeroSignal(31) => 
                           X_Logic0_port, zeroSignal(30) => X_Logic0_port, 
                           zeroSignal(29) => X_Logic0_port, zeroSignal(28) => 
                           X_Logic0_port, zeroSignal(27) => X_Logic0_port, 
                           zeroSignal(26) => X_Logic0_port, zeroSignal(25) => 
                           X_Logic0_port, zeroSignal(24) => X_Logic0_port, 
                           zeroSignal(23) => X_Logic0_port, zeroSignal(22) => 
                           X_Logic0_port, zeroSignal(21) => X_Logic0_port, 
                           zeroSignal(20) => X_Logic0_port, zeroSignal(19) => 
                           X_Logic0_port, zeroSignal(18) => X_Logic0_port, 
                           zeroSignal(17) => X_Logic0_port, zeroSignal(16) => 
                           X_Logic0_port, zeroSignal(15) => X_Logic0_port, 
                           zeroSignal(14) => X_Logic0_port, zeroSignal(13) => 
                           X_Logic0_port, zeroSignal(12) => X_Logic0_port, 
                           zeroSignal(11) => X_Logic0_port, zeroSignal(10) => 
                           X_Logic0_port, zeroSignal(9) => X_Logic0_port, 
                           zeroSignal(8) => X_Logic0_port, zeroSignal(7) => 
                           X_Logic0_port, zeroSignal(6) => X_Logic0_port, 
                           zeroSignal(5) => X_Logic0_port, zeroSignal(4) => 
                           X_Logic0_port, zeroSignal(3) => X_Logic0_port, 
                           zeroSignal(2) => X_Logic0_port, zeroSignal(1) => 
                           X_Logic0_port, zeroSignal(0) => X_Logic0_port, 
                           A_signal(63) => positive_inputs_30_63_port, 
                           A_signal(62) => positive_inputs_30_62_port, 
                           A_signal(61) => positive_inputs_30_61_port, 
                           A_signal(60) => positive_inputs_30_60_port, 
                           A_signal(59) => positive_inputs_30_59_port, 
                           A_signal(58) => positive_inputs_30_58_port, 
                           A_signal(57) => positive_inputs_30_57_port, 
                           A_signal(56) => positive_inputs_30_56_port, 
                           A_signal(55) => positive_inputs_30_55_port, 
                           A_signal(54) => positive_inputs_30_54_port, 
                           A_signal(53) => positive_inputs_30_53_port, 
                           A_signal(52) => positive_inputs_30_52_port, 
                           A_signal(51) => positive_inputs_30_51_port, 
                           A_signal(50) => positive_inputs_30_50_port, 
                           A_signal(49) => positive_inputs_30_49_port, 
                           A_signal(48) => positive_inputs_30_48_port, 
                           A_signal(47) => positive_inputs_30_47_port, 
                           A_signal(46) => positive_inputs_30_46_port, 
                           A_signal(45) => positive_inputs_30_45_port, 
                           A_signal(44) => positive_inputs_30_44_port, 
                           A_signal(43) => positive_inputs_30_43_port, 
                           A_signal(42) => positive_inputs_30_42_port, 
                           A_signal(41) => positive_inputs_30_41_port, 
                           A_signal(40) => positive_inputs_30_40_port, 
                           A_signal(39) => positive_inputs_30_39_port, 
                           A_signal(38) => positive_inputs_30_38_port, 
                           A_signal(37) => positive_inputs_30_37_port, 
                           A_signal(36) => positive_inputs_30_36_port, 
                           A_signal(35) => positive_inputs_30_35_port, 
                           A_signal(34) => positive_inputs_30_34_port, 
                           A_signal(33) => positive_inputs_30_33_port, 
                           A_signal(32) => positive_inputs_30_32_port, 
                           A_signal(31) => positive_inputs_30_31_port, 
                           A_signal(30) => positive_inputs_30_30_port, 
                           A_signal(29) => positive_inputs_30_29_port, 
                           A_signal(28) => positive_inputs_30_28_port, 
                           A_signal(27) => positive_inputs_30_27_port, 
                           A_signal(26) => positive_inputs_30_26_port, 
                           A_signal(25) => positive_inputs_30_25_port, 
                           A_signal(24) => positive_inputs_30_24_port, 
                           A_signal(23) => positive_inputs_30_23_port, 
                           A_signal(22) => positive_inputs_30_22_port, 
                           A_signal(21) => positive_inputs_30_21_port, 
                           A_signal(20) => positive_inputs_30_20_port, 
                           A_signal(19) => positive_inputs_30_19_port, 
                           A_signal(18) => positive_inputs_30_18_port, 
                           A_signal(17) => positive_inputs_30_17_port, 
                           A_signal(16) => positive_inputs_30_16_port, 
                           A_signal(15) => positive_inputs_30_15_port, 
                           A_signal(14) => positive_inputs_30_14_port, 
                           A_signal(13) => positive_inputs_30_13_port, 
                           A_signal(12) => positive_inputs_30_12_port, 
                           A_signal(11) => positive_inputs_30_11_port, 
                           A_signal(10) => positive_inputs_30_10_port, 
                           A_signal(9) => positive_inputs_30_9_port, 
                           A_signal(8) => positive_inputs_30_8_port, 
                           A_signal(7) => positive_inputs_30_7_port, 
                           A_signal(6) => positive_inputs_30_6_port, 
                           A_signal(5) => positive_inputs_30_5_port, 
                           A_signal(4) => positive_inputs_30_4_port, 
                           A_signal(3) => positive_inputs_30_3_port, 
                           A_signal(2) => positive_inputs_30_2_port, 
                           A_signal(1) => positive_inputs_30_1_port, 
                           A_signal(0) => n8, A_neg(63) => 
                           negative_inputs_30_63_port, A_neg(62) => 
                           negative_inputs_30_62_port, A_neg(61) => 
                           negative_inputs_30_61_port, A_neg(60) => 
                           negative_inputs_30_60_port, A_neg(59) => 
                           negative_inputs_30_59_port, A_neg(58) => 
                           negative_inputs_30_58_port, A_neg(57) => 
                           negative_inputs_30_57_port, A_neg(56) => 
                           negative_inputs_30_56_port, A_neg(55) => 
                           negative_inputs_30_55_port, A_neg(54) => 
                           negative_inputs_30_54_port, A_neg(53) => 
                           negative_inputs_30_53_port, A_neg(52) => 
                           negative_inputs_30_52_port, A_neg(51) => 
                           negative_inputs_30_51_port, A_neg(50) => 
                           negative_inputs_30_50_port, A_neg(49) => 
                           negative_inputs_30_49_port, A_neg(48) => 
                           negative_inputs_30_48_port, A_neg(47) => 
                           negative_inputs_30_47_port, A_neg(46) => 
                           negative_inputs_30_46_port, A_neg(45) => 
                           negative_inputs_30_45_port, A_neg(44) => 
                           negative_inputs_30_44_port, A_neg(43) => 
                           negative_inputs_30_43_port, A_neg(42) => 
                           negative_inputs_30_42_port, A_neg(41) => 
                           negative_inputs_30_41_port, A_neg(40) => 
                           negative_inputs_30_40_port, A_neg(39) => 
                           negative_inputs_30_39_port, A_neg(38) => 
                           negative_inputs_30_38_port, A_neg(37) => 
                           negative_inputs_30_37_port, A_neg(36) => 
                           negative_inputs_30_36_port, A_neg(35) => 
                           negative_inputs_30_35_port, A_neg(34) => 
                           negative_inputs_30_34_port, A_neg(33) => 
                           negative_inputs_30_33_port, A_neg(32) => 
                           negative_inputs_30_32_port, A_neg(31) => 
                           negative_inputs_30_31_port, A_neg(30) => 
                           negative_inputs_30_30_port, A_neg(29) => 
                           negative_inputs_30_29_port, A_neg(28) => 
                           negative_inputs_30_28_port, A_neg(27) => 
                           negative_inputs_30_27_port, A_neg(26) => 
                           negative_inputs_30_26_port, A_neg(25) => 
                           negative_inputs_30_25_port, A_neg(24) => 
                           negative_inputs_30_24_port, A_neg(23) => 
                           negative_inputs_30_23_port, A_neg(22) => 
                           negative_inputs_30_22_port, A_neg(21) => 
                           negative_inputs_30_21_port, A_neg(20) => 
                           negative_inputs_30_20_port, A_neg(19) => 
                           negative_inputs_30_19_port, A_neg(18) => 
                           negative_inputs_30_18_port, A_neg(17) => 
                           negative_inputs_30_17_port, A_neg(16) => 
                           negative_inputs_30_16_port, A_neg(15) => 
                           negative_inputs_30_15_port, A_neg(14) => 
                           negative_inputs_30_14_port, A_neg(13) => 
                           negative_inputs_30_13_port, A_neg(12) => 
                           negative_inputs_30_12_port, A_neg(11) => 
                           negative_inputs_30_11_port, A_neg(10) => 
                           negative_inputs_30_10_port, A_neg(9) => 
                           negative_inputs_30_9_port, A_neg(8) => 
                           negative_inputs_30_8_port, A_neg(7) => 
                           negative_inputs_30_7_port, A_neg(6) => 
                           negative_inputs_30_6_port, A_neg(5) => 
                           negative_inputs_30_5_port, A_neg(4) => 
                           negative_inputs_30_4_port, A_neg(3) => 
                           negative_inputs_30_3_port, A_neg(2) => 
                           negative_inputs_30_2_port, A_neg(1) => 
                           negative_inputs_30_1_port, A_neg(0) => n8, 
                           A_shifted(63) => positive_inputs_31_63_port, 
                           A_shifted(62) => positive_inputs_31_62_port, 
                           A_shifted(61) => positive_inputs_31_61_port, 
                           A_shifted(60) => positive_inputs_31_60_port, 
                           A_shifted(59) => positive_inputs_31_59_port, 
                           A_shifted(58) => positive_inputs_31_58_port, 
                           A_shifted(57) => positive_inputs_31_57_port, 
                           A_shifted(56) => positive_inputs_31_56_port, 
                           A_shifted(55) => positive_inputs_31_55_port, 
                           A_shifted(54) => positive_inputs_31_54_port, 
                           A_shifted(53) => positive_inputs_31_53_port, 
                           A_shifted(52) => positive_inputs_31_52_port, 
                           A_shifted(51) => positive_inputs_31_51_port, 
                           A_shifted(50) => positive_inputs_31_50_port, 
                           A_shifted(49) => positive_inputs_31_49_port, 
                           A_shifted(48) => positive_inputs_31_48_port, 
                           A_shifted(47) => positive_inputs_31_47_port, 
                           A_shifted(46) => positive_inputs_31_46_port, 
                           A_shifted(45) => positive_inputs_31_45_port, 
                           A_shifted(44) => positive_inputs_31_44_port, 
                           A_shifted(43) => positive_inputs_31_43_port, 
                           A_shifted(42) => positive_inputs_31_42_port, 
                           A_shifted(41) => positive_inputs_31_41_port, 
                           A_shifted(40) => positive_inputs_31_40_port, 
                           A_shifted(39) => positive_inputs_31_39_port, 
                           A_shifted(38) => positive_inputs_31_38_port, 
                           A_shifted(37) => positive_inputs_31_37_port, 
                           A_shifted(36) => positive_inputs_31_36_port, 
                           A_shifted(35) => positive_inputs_31_35_port, 
                           A_shifted(34) => positive_inputs_31_34_port, 
                           A_shifted(33) => positive_inputs_31_33_port, 
                           A_shifted(32) => positive_inputs_31_32_port, 
                           A_shifted(31) => positive_inputs_31_31_port, 
                           A_shifted(30) => positive_inputs_31_30_port, 
                           A_shifted(29) => positive_inputs_31_29_port, 
                           A_shifted(28) => positive_inputs_31_28_port, 
                           A_shifted(27) => positive_inputs_31_27_port, 
                           A_shifted(26) => positive_inputs_31_26_port, 
                           A_shifted(25) => positive_inputs_31_25_port, 
                           A_shifted(24) => positive_inputs_31_24_port, 
                           A_shifted(23) => positive_inputs_31_23_port, 
                           A_shifted(22) => positive_inputs_31_22_port, 
                           A_shifted(21) => positive_inputs_31_21_port, 
                           A_shifted(20) => positive_inputs_31_20_port, 
                           A_shifted(19) => positive_inputs_31_19_port, 
                           A_shifted(18) => positive_inputs_31_18_port, 
                           A_shifted(17) => positive_inputs_31_17_port, 
                           A_shifted(16) => positive_inputs_31_16_port, 
                           A_shifted(15) => positive_inputs_31_15_port, 
                           A_shifted(14) => positive_inputs_31_14_port, 
                           A_shifted(13) => positive_inputs_31_13_port, 
                           A_shifted(12) => positive_inputs_31_12_port, 
                           A_shifted(11) => positive_inputs_31_11_port, 
                           A_shifted(10) => positive_inputs_31_10_port, 
                           A_shifted(9) => positive_inputs_31_9_port, 
                           A_shifted(8) => positive_inputs_31_8_port, 
                           A_shifted(7) => positive_inputs_31_7_port, 
                           A_shifted(6) => positive_inputs_31_6_port, 
                           A_shifted(5) => positive_inputs_31_5_port, 
                           A_shifted(4) => positive_inputs_31_4_port, 
                           A_shifted(3) => positive_inputs_31_3_port, 
                           A_shifted(2) => positive_inputs_31_2_port, 
                           A_shifted(1) => positive_inputs_31_1_port, 
                           A_shifted(0) => n8, A_neg_shifted(63) => 
                           negative_inputs_31_63_port, A_neg_shifted(62) => 
                           negative_inputs_31_62_port, A_neg_shifted(61) => 
                           negative_inputs_31_61_port, A_neg_shifted(60) => 
                           negative_inputs_31_60_port, A_neg_shifted(59) => 
                           negative_inputs_31_59_port, A_neg_shifted(58) => 
                           negative_inputs_31_58_port, A_neg_shifted(57) => 
                           negative_inputs_31_57_port, A_neg_shifted(56) => 
                           negative_inputs_31_56_port, A_neg_shifted(55) => 
                           negative_inputs_31_55_port, A_neg_shifted(54) => 
                           negative_inputs_31_54_port, A_neg_shifted(53) => 
                           negative_inputs_31_53_port, A_neg_shifted(52) => 
                           negative_inputs_31_52_port, A_neg_shifted(51) => 
                           negative_inputs_31_51_port, A_neg_shifted(50) => 
                           negative_inputs_31_50_port, A_neg_shifted(49) => 
                           negative_inputs_31_49_port, A_neg_shifted(48) => 
                           negative_inputs_31_48_port, A_neg_shifted(47) => 
                           negative_inputs_31_47_port, A_neg_shifted(46) => 
                           negative_inputs_31_46_port, A_neg_shifted(45) => 
                           negative_inputs_31_45_port, A_neg_shifted(44) => 
                           negative_inputs_31_44_port, A_neg_shifted(43) => 
                           negative_inputs_31_43_port, A_neg_shifted(42) => 
                           negative_inputs_31_42_port, A_neg_shifted(41) => 
                           negative_inputs_31_41_port, A_neg_shifted(40) => 
                           negative_inputs_31_40_port, A_neg_shifted(39) => 
                           negative_inputs_31_39_port, A_neg_shifted(38) => 
                           negative_inputs_31_38_port, A_neg_shifted(37) => 
                           negative_inputs_31_37_port, A_neg_shifted(36) => 
                           negative_inputs_31_36_port, A_neg_shifted(35) => 
                           negative_inputs_31_35_port, A_neg_shifted(34) => 
                           negative_inputs_31_34_port, A_neg_shifted(33) => 
                           negative_inputs_31_33_port, A_neg_shifted(32) => 
                           negative_inputs_31_32_port, A_neg_shifted(31) => 
                           negative_inputs_31_31_port, A_neg_shifted(30) => 
                           negative_inputs_31_30_port, A_neg_shifted(29) => 
                           negative_inputs_31_29_port, A_neg_shifted(28) => 
                           negative_inputs_31_28_port, A_neg_shifted(27) => 
                           negative_inputs_31_27_port, A_neg_shifted(26) => 
                           negative_inputs_31_26_port, A_neg_shifted(25) => 
                           negative_inputs_31_25_port, A_neg_shifted(24) => 
                           negative_inputs_31_24_port, A_neg_shifted(23) => 
                           negative_inputs_31_23_port, A_neg_shifted(22) => 
                           negative_inputs_31_22_port, A_neg_shifted(21) => 
                           negative_inputs_31_21_port, A_neg_shifted(20) => 
                           negative_inputs_31_20_port, A_neg_shifted(19) => 
                           negative_inputs_31_19_port, A_neg_shifted(18) => 
                           negative_inputs_31_18_port, A_neg_shifted(17) => 
                           negative_inputs_31_17_port, A_neg_shifted(16) => 
                           negative_inputs_31_16_port, A_neg_shifted(15) => 
                           negative_inputs_31_15_port, A_neg_shifted(14) => 
                           negative_inputs_31_14_port, A_neg_shifted(13) => 
                           negative_inputs_31_13_port, A_neg_shifted(12) => 
                           negative_inputs_31_12_port, A_neg_shifted(11) => 
                           negative_inputs_31_11_port, A_neg_shifted(10) => 
                           negative_inputs_31_10_port, A_neg_shifted(9) => 
                           negative_inputs_31_9_port, A_neg_shifted(8) => 
                           negative_inputs_31_8_port, A_neg_shifted(7) => 
                           negative_inputs_31_7_port, A_neg_shifted(6) => 
                           negative_inputs_31_6_port, A_neg_shifted(5) => 
                           negative_inputs_31_5_port, A_neg_shifted(4) => 
                           negative_inputs_31_4_port, A_neg_shifted(3) => 
                           negative_inputs_31_3_port, A_neg_shifted(2) => 
                           negative_inputs_31_2_port, A_neg_shifted(1) => 
                           negative_inputs_31_1_port, A_neg_shifted(0) => n8, 
                           Sel(2) => sel_15_2_port, Sel(1) => sel_15_1_port, 
                           Sel(0) => sel_15_0_port, Y(63) => 
                           MuxOutputs_15_63_port, Y(62) => 
                           MuxOutputs_15_62_port, Y(61) => 
                           MuxOutputs_15_61_port, Y(60) => 
                           MuxOutputs_15_60_port, Y(59) => 
                           MuxOutputs_15_59_port, Y(58) => 
                           MuxOutputs_15_58_port, Y(57) => 
                           MuxOutputs_15_57_port, Y(56) => 
                           MuxOutputs_15_56_port, Y(55) => 
                           MuxOutputs_15_55_port, Y(54) => 
                           MuxOutputs_15_54_port, Y(53) => 
                           MuxOutputs_15_53_port, Y(52) => 
                           MuxOutputs_15_52_port, Y(51) => 
                           MuxOutputs_15_51_port, Y(50) => 
                           MuxOutputs_15_50_port, Y(49) => 
                           MuxOutputs_15_49_port, Y(48) => 
                           MuxOutputs_15_48_port, Y(47) => 
                           MuxOutputs_15_47_port, Y(46) => 
                           MuxOutputs_15_46_port, Y(45) => 
                           MuxOutputs_15_45_port, Y(44) => 
                           MuxOutputs_15_44_port, Y(43) => 
                           MuxOutputs_15_43_port, Y(42) => 
                           MuxOutputs_15_42_port, Y(41) => 
                           MuxOutputs_15_41_port, Y(40) => 
                           MuxOutputs_15_40_port, Y(39) => 
                           MuxOutputs_15_39_port, Y(38) => 
                           MuxOutputs_15_38_port, Y(37) => 
                           MuxOutputs_15_37_port, Y(36) => 
                           MuxOutputs_15_36_port, Y(35) => 
                           MuxOutputs_15_35_port, Y(34) => 
                           MuxOutputs_15_34_port, Y(33) => 
                           MuxOutputs_15_33_port, Y(32) => 
                           MuxOutputs_15_32_port, Y(31) => 
                           MuxOutputs_15_31_port, Y(30) => 
                           MuxOutputs_15_30_port, Y(29) => 
                           MuxOutputs_15_29_port, Y(28) => 
                           MuxOutputs_15_28_port, Y(27) => 
                           MuxOutputs_15_27_port, Y(26) => 
                           MuxOutputs_15_26_port, Y(25) => 
                           MuxOutputs_15_25_port, Y(24) => 
                           MuxOutputs_15_24_port, Y(23) => 
                           MuxOutputs_15_23_port, Y(22) => 
                           MuxOutputs_15_22_port, Y(21) => 
                           MuxOutputs_15_21_port, Y(20) => 
                           MuxOutputs_15_20_port, Y(19) => 
                           MuxOutputs_15_19_port, Y(18) => 
                           MuxOutputs_15_18_port, Y(17) => 
                           MuxOutputs_15_17_port, Y(16) => 
                           MuxOutputs_15_16_port, Y(15) => 
                           MuxOutputs_15_15_port, Y(14) => 
                           MuxOutputs_15_14_port, Y(13) => 
                           MuxOutputs_15_13_port, Y(12) => 
                           MuxOutputs_15_12_port, Y(11) => 
                           MuxOutputs_15_11_port, Y(10) => 
                           MuxOutputs_15_10_port, Y(9) => MuxOutputs_15_9_port,
                           Y(8) => MuxOutputs_15_8_port, Y(7) => 
                           MuxOutputs_15_7_port, Y(6) => MuxOutputs_15_6_port, 
                           Y(5) => MuxOutputs_15_5_port, Y(4) => 
                           MuxOutputs_15_4_port, Y(3) => MuxOutputs_15_3_port, 
                           Y(2) => MuxOutputs_15_2_port, Y(1) => 
                           MuxOutputs_15_1_port, Y(0) => MuxOutputs_15_0_port);
   SUM0 : RCA_NbitRca64_31 port map( A(63) => MuxOutputs_0_63_port, A(62) => 
                           MuxOutputs_0_62_port, A(61) => MuxOutputs_0_61_port,
                           A(60) => MuxOutputs_0_60_port, A(59) => 
                           MuxOutputs_0_59_port, A(58) => MuxOutputs_0_58_port,
                           A(57) => MuxOutputs_0_57_port, A(56) => 
                           MuxOutputs_0_56_port, A(55) => MuxOutputs_0_55_port,
                           A(54) => MuxOutputs_0_54_port, A(53) => 
                           MuxOutputs_0_53_port, A(52) => MuxOutputs_0_52_port,
                           A(51) => MuxOutputs_0_51_port, A(50) => 
                           MuxOutputs_0_50_port, A(49) => MuxOutputs_0_49_port,
                           A(48) => MuxOutputs_0_48_port, A(47) => 
                           MuxOutputs_0_47_port, A(46) => MuxOutputs_0_46_port,
                           A(45) => MuxOutputs_0_45_port, A(44) => 
                           MuxOutputs_0_44_port, A(43) => MuxOutputs_0_43_port,
                           A(42) => MuxOutputs_0_42_port, A(41) => 
                           MuxOutputs_0_41_port, A(40) => MuxOutputs_0_40_port,
                           A(39) => MuxOutputs_0_39_port, A(38) => 
                           MuxOutputs_0_38_port, A(37) => MuxOutputs_0_37_port,
                           A(36) => MuxOutputs_0_36_port, A(35) => 
                           MuxOutputs_0_35_port, A(34) => MuxOutputs_0_34_port,
                           A(33) => MuxOutputs_0_33_port, A(32) => 
                           MuxOutputs_0_32_port, A(31) => MuxOutputs_0_31_port,
                           A(30) => MuxOutputs_0_30_port, A(29) => 
                           MuxOutputs_0_29_port, A(28) => MuxOutputs_0_28_port,
                           A(27) => MuxOutputs_0_27_port, A(26) => 
                           MuxOutputs_0_26_port, A(25) => MuxOutputs_0_25_port,
                           A(24) => MuxOutputs_0_24_port, A(23) => 
                           MuxOutputs_0_23_port, A(22) => MuxOutputs_0_22_port,
                           A(21) => MuxOutputs_0_21_port, A(20) => 
                           MuxOutputs_0_20_port, A(19) => MuxOutputs_0_19_port,
                           A(18) => MuxOutputs_0_18_port, A(17) => 
                           MuxOutputs_0_17_port, A(16) => MuxOutputs_0_16_port,
                           A(15) => MuxOutputs_0_15_port, A(14) => 
                           MuxOutputs_0_14_port, A(13) => MuxOutputs_0_13_port,
                           A(12) => MuxOutputs_0_12_port, A(11) => 
                           MuxOutputs_0_11_port, A(10) => MuxOutputs_0_10_port,
                           A(9) => MuxOutputs_0_9_port, A(8) => 
                           MuxOutputs_0_8_port, A(7) => MuxOutputs_0_7_port, 
                           A(6) => MuxOutputs_0_6_port, A(5) => 
                           MuxOutputs_0_5_port, A(4) => MuxOutputs_0_4_port, 
                           A(3) => MuxOutputs_0_3_port, A(2) => 
                           MuxOutputs_0_2_port, A(1) => MuxOutputs_0_1_port, 
                           A(0) => MuxOutputs_0_0_port, B(63) => 
                           MuxOutputs_1_63_port, B(62) => MuxOutputs_1_62_port,
                           B(61) => MuxOutputs_1_61_port, B(60) => 
                           MuxOutputs_1_60_port, B(59) => MuxOutputs_1_59_port,
                           B(58) => MuxOutputs_1_58_port, B(57) => 
                           MuxOutputs_1_57_port, B(56) => MuxOutputs_1_56_port,
                           B(55) => MuxOutputs_1_55_port, B(54) => 
                           MuxOutputs_1_54_port, B(53) => MuxOutputs_1_53_port,
                           B(52) => MuxOutputs_1_52_port, B(51) => 
                           MuxOutputs_1_51_port, B(50) => MuxOutputs_1_50_port,
                           B(49) => MuxOutputs_1_49_port, B(48) => 
                           MuxOutputs_1_48_port, B(47) => MuxOutputs_1_47_port,
                           B(46) => MuxOutputs_1_46_port, B(45) => 
                           MuxOutputs_1_45_port, B(44) => MuxOutputs_1_44_port,
                           B(43) => MuxOutputs_1_43_port, B(42) => 
                           MuxOutputs_1_42_port, B(41) => MuxOutputs_1_41_port,
                           B(40) => MuxOutputs_1_40_port, B(39) => 
                           MuxOutputs_1_39_port, B(38) => MuxOutputs_1_38_port,
                           B(37) => MuxOutputs_1_37_port, B(36) => 
                           MuxOutputs_1_36_port, B(35) => MuxOutputs_1_35_port,
                           B(34) => MuxOutputs_1_34_port, B(33) => 
                           MuxOutputs_1_33_port, B(32) => MuxOutputs_1_32_port,
                           B(31) => MuxOutputs_1_31_port, B(30) => 
                           MuxOutputs_1_30_port, B(29) => MuxOutputs_1_29_port,
                           B(28) => MuxOutputs_1_28_port, B(27) => 
                           MuxOutputs_1_27_port, B(26) => MuxOutputs_1_26_port,
                           B(25) => MuxOutputs_1_25_port, B(24) => 
                           MuxOutputs_1_24_port, B(23) => MuxOutputs_1_23_port,
                           B(22) => MuxOutputs_1_22_port, B(21) => 
                           MuxOutputs_1_21_port, B(20) => MuxOutputs_1_20_port,
                           B(19) => MuxOutputs_1_19_port, B(18) => 
                           MuxOutputs_1_18_port, B(17) => MuxOutputs_1_17_port,
                           B(16) => MuxOutputs_1_16_port, B(15) => 
                           MuxOutputs_1_15_port, B(14) => MuxOutputs_1_14_port,
                           B(13) => MuxOutputs_1_13_port, B(12) => 
                           MuxOutputs_1_12_port, B(11) => MuxOutputs_1_11_port,
                           B(10) => MuxOutputs_1_10_port, B(9) => 
                           MuxOutputs_1_9_port, B(8) => MuxOutputs_1_8_port, 
                           B(7) => MuxOutputs_1_7_port, B(6) => 
                           MuxOutputs_1_6_port, B(5) => MuxOutputs_1_5_port, 
                           B(4) => MuxOutputs_1_4_port, B(3) => 
                           MuxOutputs_1_3_port, B(2) => MuxOutputs_1_2_port, 
                           B(1) => MuxOutputs_1_1_port, B(0) => 
                           MuxOutputs_1_0_port, Ci => X_Logic0_port, S(63) => 
                           SumOutputs_0_63_port, S(62) => SumOutputs_0_62_port,
                           S(61) => SumOutputs_0_61_port, S(60) => 
                           SumOutputs_0_60_port, S(59) => SumOutputs_0_59_port,
                           S(58) => SumOutputs_0_58_port, S(57) => 
                           SumOutputs_0_57_port, S(56) => SumOutputs_0_56_port,
                           S(55) => SumOutputs_0_55_port, S(54) => 
                           SumOutputs_0_54_port, S(53) => SumOutputs_0_53_port,
                           S(52) => SumOutputs_0_52_port, S(51) => 
                           SumOutputs_0_51_port, S(50) => SumOutputs_0_50_port,
                           S(49) => SumOutputs_0_49_port, S(48) => 
                           SumOutputs_0_48_port, S(47) => SumOutputs_0_47_port,
                           S(46) => SumOutputs_0_46_port, S(45) => 
                           SumOutputs_0_45_port, S(44) => SumOutputs_0_44_port,
                           S(43) => SumOutputs_0_43_port, S(42) => 
                           SumOutputs_0_42_port, S(41) => SumOutputs_0_41_port,
                           S(40) => SumOutputs_0_40_port, S(39) => 
                           SumOutputs_0_39_port, S(38) => SumOutputs_0_38_port,
                           S(37) => SumOutputs_0_37_port, S(36) => 
                           SumOutputs_0_36_port, S(35) => SumOutputs_0_35_port,
                           S(34) => SumOutputs_0_34_port, S(33) => 
                           SumOutputs_0_33_port, S(32) => SumOutputs_0_32_port,
                           S(31) => SumOutputs_0_31_port, S(30) => 
                           SumOutputs_0_30_port, S(29) => SumOutputs_0_29_port,
                           S(28) => SumOutputs_0_28_port, S(27) => 
                           SumOutputs_0_27_port, S(26) => SumOutputs_0_26_port,
                           S(25) => SumOutputs_0_25_port, S(24) => 
                           SumOutputs_0_24_port, S(23) => SumOutputs_0_23_port,
                           S(22) => SumOutputs_0_22_port, S(21) => 
                           SumOutputs_0_21_port, S(20) => SumOutputs_0_20_port,
                           S(19) => SumOutputs_0_19_port, S(18) => 
                           SumOutputs_0_18_port, S(17) => SumOutputs_0_17_port,
                           S(16) => SumOutputs_0_16_port, S(15) => 
                           SumOutputs_0_15_port, S(14) => SumOutputs_0_14_port,
                           S(13) => SumOutputs_0_13_port, S(12) => 
                           SumOutputs_0_12_port, S(11) => SumOutputs_0_11_port,
                           S(10) => SumOutputs_0_10_port, S(9) => 
                           SumOutputs_0_9_port, S(8) => SumOutputs_0_8_port, 
                           S(7) => SumOutputs_0_7_port, S(6) => 
                           SumOutputs_0_6_port, S(5) => SumOutputs_0_5_port, 
                           S(4) => SumOutputs_0_4_port, S(3) => 
                           SumOutputs_0_3_port, S(2) => SumOutputs_0_2_port, 
                           S(1) => SumOutputs_0_1_port, S(0) => 
                           SumOutputs_0_0_port, Co => n_1127);
   SUMI_1 : RCA_NbitRca64_30 port map( A(63) => MuxOutputs_2_63_port, A(62) => 
                           MuxOutputs_2_62_port, A(61) => MuxOutputs_2_61_port,
                           A(60) => MuxOutputs_2_60_port, A(59) => 
                           MuxOutputs_2_59_port, A(58) => MuxOutputs_2_58_port,
                           A(57) => MuxOutputs_2_57_port, A(56) => 
                           MuxOutputs_2_56_port, A(55) => MuxOutputs_2_55_port,
                           A(54) => MuxOutputs_2_54_port, A(53) => 
                           MuxOutputs_2_53_port, A(52) => MuxOutputs_2_52_port,
                           A(51) => MuxOutputs_2_51_port, A(50) => 
                           MuxOutputs_2_50_port, A(49) => MuxOutputs_2_49_port,
                           A(48) => MuxOutputs_2_48_port, A(47) => 
                           MuxOutputs_2_47_port, A(46) => MuxOutputs_2_46_port,
                           A(45) => MuxOutputs_2_45_port, A(44) => 
                           MuxOutputs_2_44_port, A(43) => MuxOutputs_2_43_port,
                           A(42) => MuxOutputs_2_42_port, A(41) => 
                           MuxOutputs_2_41_port, A(40) => MuxOutputs_2_40_port,
                           A(39) => MuxOutputs_2_39_port, A(38) => 
                           MuxOutputs_2_38_port, A(37) => MuxOutputs_2_37_port,
                           A(36) => MuxOutputs_2_36_port, A(35) => 
                           MuxOutputs_2_35_port, A(34) => MuxOutputs_2_34_port,
                           A(33) => MuxOutputs_2_33_port, A(32) => 
                           MuxOutputs_2_32_port, A(31) => MuxOutputs_2_31_port,
                           A(30) => MuxOutputs_2_30_port, A(29) => 
                           MuxOutputs_2_29_port, A(28) => MuxOutputs_2_28_port,
                           A(27) => MuxOutputs_2_27_port, A(26) => 
                           MuxOutputs_2_26_port, A(25) => MuxOutputs_2_25_port,
                           A(24) => MuxOutputs_2_24_port, A(23) => 
                           MuxOutputs_2_23_port, A(22) => MuxOutputs_2_22_port,
                           A(21) => MuxOutputs_2_21_port, A(20) => 
                           MuxOutputs_2_20_port, A(19) => MuxOutputs_2_19_port,
                           A(18) => MuxOutputs_2_18_port, A(17) => 
                           MuxOutputs_2_17_port, A(16) => MuxOutputs_2_16_port,
                           A(15) => MuxOutputs_2_15_port, A(14) => 
                           MuxOutputs_2_14_port, A(13) => MuxOutputs_2_13_port,
                           A(12) => MuxOutputs_2_12_port, A(11) => 
                           MuxOutputs_2_11_port, A(10) => MuxOutputs_2_10_port,
                           A(9) => MuxOutputs_2_9_port, A(8) => 
                           MuxOutputs_2_8_port, A(7) => MuxOutputs_2_7_port, 
                           A(6) => MuxOutputs_2_6_port, A(5) => 
                           MuxOutputs_2_5_port, A(4) => MuxOutputs_2_4_port, 
                           A(3) => MuxOutputs_2_3_port, A(2) => 
                           MuxOutputs_2_2_port, A(1) => MuxOutputs_2_1_port, 
                           A(0) => MuxOutputs_2_0_port, B(63) => 
                           SumOutputs_0_63_port, B(62) => SumOutputs_0_62_port,
                           B(61) => SumOutputs_0_61_port, B(60) => 
                           SumOutputs_0_60_port, B(59) => SumOutputs_0_59_port,
                           B(58) => SumOutputs_0_58_port, B(57) => 
                           SumOutputs_0_57_port, B(56) => SumOutputs_0_56_port,
                           B(55) => SumOutputs_0_55_port, B(54) => 
                           SumOutputs_0_54_port, B(53) => SumOutputs_0_53_port,
                           B(52) => SumOutputs_0_52_port, B(51) => 
                           SumOutputs_0_51_port, B(50) => SumOutputs_0_50_port,
                           B(49) => SumOutputs_0_49_port, B(48) => 
                           SumOutputs_0_48_port, B(47) => SumOutputs_0_47_port,
                           B(46) => SumOutputs_0_46_port, B(45) => 
                           SumOutputs_0_45_port, B(44) => SumOutputs_0_44_port,
                           B(43) => SumOutputs_0_43_port, B(42) => 
                           SumOutputs_0_42_port, B(41) => SumOutputs_0_41_port,
                           B(40) => SumOutputs_0_40_port, B(39) => 
                           SumOutputs_0_39_port, B(38) => SumOutputs_0_38_port,
                           B(37) => SumOutputs_0_37_port, B(36) => 
                           SumOutputs_0_36_port, B(35) => SumOutputs_0_35_port,
                           B(34) => SumOutputs_0_34_port, B(33) => 
                           SumOutputs_0_33_port, B(32) => SumOutputs_0_32_port,
                           B(31) => SumOutputs_0_31_port, B(30) => 
                           SumOutputs_0_30_port, B(29) => SumOutputs_0_29_port,
                           B(28) => SumOutputs_0_28_port, B(27) => 
                           SumOutputs_0_27_port, B(26) => SumOutputs_0_26_port,
                           B(25) => SumOutputs_0_25_port, B(24) => 
                           SumOutputs_0_24_port, B(23) => SumOutputs_0_23_port,
                           B(22) => SumOutputs_0_22_port, B(21) => 
                           SumOutputs_0_21_port, B(20) => SumOutputs_0_20_port,
                           B(19) => SumOutputs_0_19_port, B(18) => 
                           SumOutputs_0_18_port, B(17) => SumOutputs_0_17_port,
                           B(16) => SumOutputs_0_16_port, B(15) => 
                           SumOutputs_0_15_port, B(14) => SumOutputs_0_14_port,
                           B(13) => SumOutputs_0_13_port, B(12) => 
                           SumOutputs_0_12_port, B(11) => SumOutputs_0_11_port,
                           B(10) => SumOutputs_0_10_port, B(9) => 
                           SumOutputs_0_9_port, B(8) => SumOutputs_0_8_port, 
                           B(7) => SumOutputs_0_7_port, B(6) => 
                           SumOutputs_0_6_port, B(5) => SumOutputs_0_5_port, 
                           B(4) => SumOutputs_0_4_port, B(3) => 
                           SumOutputs_0_3_port, B(2) => SumOutputs_0_2_port, 
                           B(1) => SumOutputs_0_1_port, B(0) => 
                           SumOutputs_0_0_port, Ci => X_Logic0_port, S(63) => 
                           SumOutputs_1_63_port, S(62) => SumOutputs_1_62_port,
                           S(61) => SumOutputs_1_61_port, S(60) => 
                           SumOutputs_1_60_port, S(59) => SumOutputs_1_59_port,
                           S(58) => SumOutputs_1_58_port, S(57) => 
                           SumOutputs_1_57_port, S(56) => SumOutputs_1_56_port,
                           S(55) => SumOutputs_1_55_port, S(54) => 
                           SumOutputs_1_54_port, S(53) => SumOutputs_1_53_port,
                           S(52) => SumOutputs_1_52_port, S(51) => 
                           SumOutputs_1_51_port, S(50) => SumOutputs_1_50_port,
                           S(49) => SumOutputs_1_49_port, S(48) => 
                           SumOutputs_1_48_port, S(47) => SumOutputs_1_47_port,
                           S(46) => SumOutputs_1_46_port, S(45) => 
                           SumOutputs_1_45_port, S(44) => SumOutputs_1_44_port,
                           S(43) => SumOutputs_1_43_port, S(42) => 
                           SumOutputs_1_42_port, S(41) => SumOutputs_1_41_port,
                           S(40) => SumOutputs_1_40_port, S(39) => 
                           SumOutputs_1_39_port, S(38) => SumOutputs_1_38_port,
                           S(37) => SumOutputs_1_37_port, S(36) => 
                           SumOutputs_1_36_port, S(35) => SumOutputs_1_35_port,
                           S(34) => SumOutputs_1_34_port, S(33) => 
                           SumOutputs_1_33_port, S(32) => SumOutputs_1_32_port,
                           S(31) => SumOutputs_1_31_port, S(30) => 
                           SumOutputs_1_30_port, S(29) => SumOutputs_1_29_port,
                           S(28) => SumOutputs_1_28_port, S(27) => 
                           SumOutputs_1_27_port, S(26) => SumOutputs_1_26_port,
                           S(25) => SumOutputs_1_25_port, S(24) => 
                           SumOutputs_1_24_port, S(23) => SumOutputs_1_23_port,
                           S(22) => SumOutputs_1_22_port, S(21) => 
                           SumOutputs_1_21_port, S(20) => SumOutputs_1_20_port,
                           S(19) => SumOutputs_1_19_port, S(18) => 
                           SumOutputs_1_18_port, S(17) => SumOutputs_1_17_port,
                           S(16) => SumOutputs_1_16_port, S(15) => 
                           SumOutputs_1_15_port, S(14) => SumOutputs_1_14_port,
                           S(13) => SumOutputs_1_13_port, S(12) => 
                           SumOutputs_1_12_port, S(11) => SumOutputs_1_11_port,
                           S(10) => SumOutputs_1_10_port, S(9) => 
                           SumOutputs_1_9_port, S(8) => SumOutputs_1_8_port, 
                           S(7) => SumOutputs_1_7_port, S(6) => 
                           SumOutputs_1_6_port, S(5) => SumOutputs_1_5_port, 
                           S(4) => SumOutputs_1_4_port, S(3) => 
                           SumOutputs_1_3_port, S(2) => SumOutputs_1_2_port, 
                           S(1) => SumOutputs_1_1_port, S(0) => 
                           SumOutputs_1_0_port, Co => n_1128);
   SUMI_2 : RCA_NbitRca64_29 port map( A(63) => MuxOutputs_3_63_port, A(62) => 
                           MuxOutputs_3_62_port, A(61) => MuxOutputs_3_61_port,
                           A(60) => MuxOutputs_3_60_port, A(59) => 
                           MuxOutputs_3_59_port, A(58) => MuxOutputs_3_58_port,
                           A(57) => MuxOutputs_3_57_port, A(56) => 
                           MuxOutputs_3_56_port, A(55) => MuxOutputs_3_55_port,
                           A(54) => MuxOutputs_3_54_port, A(53) => 
                           MuxOutputs_3_53_port, A(52) => MuxOutputs_3_52_port,
                           A(51) => MuxOutputs_3_51_port, A(50) => 
                           MuxOutputs_3_50_port, A(49) => MuxOutputs_3_49_port,
                           A(48) => MuxOutputs_3_48_port, A(47) => 
                           MuxOutputs_3_47_port, A(46) => MuxOutputs_3_46_port,
                           A(45) => MuxOutputs_3_45_port, A(44) => 
                           MuxOutputs_3_44_port, A(43) => MuxOutputs_3_43_port,
                           A(42) => MuxOutputs_3_42_port, A(41) => 
                           MuxOutputs_3_41_port, A(40) => MuxOutputs_3_40_port,
                           A(39) => MuxOutputs_3_39_port, A(38) => 
                           MuxOutputs_3_38_port, A(37) => MuxOutputs_3_37_port,
                           A(36) => MuxOutputs_3_36_port, A(35) => 
                           MuxOutputs_3_35_port, A(34) => MuxOutputs_3_34_port,
                           A(33) => MuxOutputs_3_33_port, A(32) => 
                           MuxOutputs_3_32_port, A(31) => MuxOutputs_3_31_port,
                           A(30) => MuxOutputs_3_30_port, A(29) => 
                           MuxOutputs_3_29_port, A(28) => MuxOutputs_3_28_port,
                           A(27) => MuxOutputs_3_27_port, A(26) => 
                           MuxOutputs_3_26_port, A(25) => MuxOutputs_3_25_port,
                           A(24) => MuxOutputs_3_24_port, A(23) => 
                           MuxOutputs_3_23_port, A(22) => MuxOutputs_3_22_port,
                           A(21) => MuxOutputs_3_21_port, A(20) => 
                           MuxOutputs_3_20_port, A(19) => MuxOutputs_3_19_port,
                           A(18) => MuxOutputs_3_18_port, A(17) => 
                           MuxOutputs_3_17_port, A(16) => MuxOutputs_3_16_port,
                           A(15) => MuxOutputs_3_15_port, A(14) => 
                           MuxOutputs_3_14_port, A(13) => MuxOutputs_3_13_port,
                           A(12) => MuxOutputs_3_12_port, A(11) => 
                           MuxOutputs_3_11_port, A(10) => MuxOutputs_3_10_port,
                           A(9) => MuxOutputs_3_9_port, A(8) => 
                           MuxOutputs_3_8_port, A(7) => MuxOutputs_3_7_port, 
                           A(6) => MuxOutputs_3_6_port, A(5) => 
                           MuxOutputs_3_5_port, A(4) => MuxOutputs_3_4_port, 
                           A(3) => MuxOutputs_3_3_port, A(2) => 
                           MuxOutputs_3_2_port, A(1) => MuxOutputs_3_1_port, 
                           A(0) => MuxOutputs_3_0_port, B(63) => 
                           SumOutputs_1_63_port, B(62) => SumOutputs_1_62_port,
                           B(61) => SumOutputs_1_61_port, B(60) => 
                           SumOutputs_1_60_port, B(59) => SumOutputs_1_59_port,
                           B(58) => SumOutputs_1_58_port, B(57) => 
                           SumOutputs_1_57_port, B(56) => SumOutputs_1_56_port,
                           B(55) => SumOutputs_1_55_port, B(54) => 
                           SumOutputs_1_54_port, B(53) => SumOutputs_1_53_port,
                           B(52) => SumOutputs_1_52_port, B(51) => 
                           SumOutputs_1_51_port, B(50) => SumOutputs_1_50_port,
                           B(49) => SumOutputs_1_49_port, B(48) => 
                           SumOutputs_1_48_port, B(47) => SumOutputs_1_47_port,
                           B(46) => SumOutputs_1_46_port, B(45) => 
                           SumOutputs_1_45_port, B(44) => SumOutputs_1_44_port,
                           B(43) => SumOutputs_1_43_port, B(42) => 
                           SumOutputs_1_42_port, B(41) => SumOutputs_1_41_port,
                           B(40) => SumOutputs_1_40_port, B(39) => 
                           SumOutputs_1_39_port, B(38) => SumOutputs_1_38_port,
                           B(37) => SumOutputs_1_37_port, B(36) => 
                           SumOutputs_1_36_port, B(35) => SumOutputs_1_35_port,
                           B(34) => SumOutputs_1_34_port, B(33) => 
                           SumOutputs_1_33_port, B(32) => SumOutputs_1_32_port,
                           B(31) => SumOutputs_1_31_port, B(30) => 
                           SumOutputs_1_30_port, B(29) => SumOutputs_1_29_port,
                           B(28) => SumOutputs_1_28_port, B(27) => 
                           SumOutputs_1_27_port, B(26) => SumOutputs_1_26_port,
                           B(25) => SumOutputs_1_25_port, B(24) => 
                           SumOutputs_1_24_port, B(23) => SumOutputs_1_23_port,
                           B(22) => SumOutputs_1_22_port, B(21) => 
                           SumOutputs_1_21_port, B(20) => SumOutputs_1_20_port,
                           B(19) => SumOutputs_1_19_port, B(18) => 
                           SumOutputs_1_18_port, B(17) => SumOutputs_1_17_port,
                           B(16) => SumOutputs_1_16_port, B(15) => 
                           SumOutputs_1_15_port, B(14) => SumOutputs_1_14_port,
                           B(13) => SumOutputs_1_13_port, B(12) => 
                           SumOutputs_1_12_port, B(11) => SumOutputs_1_11_port,
                           B(10) => SumOutputs_1_10_port, B(9) => 
                           SumOutputs_1_9_port, B(8) => SumOutputs_1_8_port, 
                           B(7) => SumOutputs_1_7_port, B(6) => 
                           SumOutputs_1_6_port, B(5) => SumOutputs_1_5_port, 
                           B(4) => SumOutputs_1_4_port, B(3) => 
                           SumOutputs_1_3_port, B(2) => SumOutputs_1_2_port, 
                           B(1) => SumOutputs_1_1_port, B(0) => 
                           SumOutputs_1_0_port, Ci => X_Logic0_port, S(63) => 
                           SumOutputs_2_63_port, S(62) => SumOutputs_2_62_port,
                           S(61) => SumOutputs_2_61_port, S(60) => 
                           SumOutputs_2_60_port, S(59) => SumOutputs_2_59_port,
                           S(58) => SumOutputs_2_58_port, S(57) => 
                           SumOutputs_2_57_port, S(56) => SumOutputs_2_56_port,
                           S(55) => SumOutputs_2_55_port, S(54) => 
                           SumOutputs_2_54_port, S(53) => SumOutputs_2_53_port,
                           S(52) => SumOutputs_2_52_port, S(51) => 
                           SumOutputs_2_51_port, S(50) => SumOutputs_2_50_port,
                           S(49) => SumOutputs_2_49_port, S(48) => 
                           SumOutputs_2_48_port, S(47) => SumOutputs_2_47_port,
                           S(46) => SumOutputs_2_46_port, S(45) => 
                           SumOutputs_2_45_port, S(44) => SumOutputs_2_44_port,
                           S(43) => SumOutputs_2_43_port, S(42) => 
                           SumOutputs_2_42_port, S(41) => SumOutputs_2_41_port,
                           S(40) => SumOutputs_2_40_port, S(39) => 
                           SumOutputs_2_39_port, S(38) => SumOutputs_2_38_port,
                           S(37) => SumOutputs_2_37_port, S(36) => 
                           SumOutputs_2_36_port, S(35) => SumOutputs_2_35_port,
                           S(34) => SumOutputs_2_34_port, S(33) => 
                           SumOutputs_2_33_port, S(32) => SumOutputs_2_32_port,
                           S(31) => SumOutputs_2_31_port, S(30) => 
                           SumOutputs_2_30_port, S(29) => SumOutputs_2_29_port,
                           S(28) => SumOutputs_2_28_port, S(27) => 
                           SumOutputs_2_27_port, S(26) => SumOutputs_2_26_port,
                           S(25) => SumOutputs_2_25_port, S(24) => 
                           SumOutputs_2_24_port, S(23) => SumOutputs_2_23_port,
                           S(22) => SumOutputs_2_22_port, S(21) => 
                           SumOutputs_2_21_port, S(20) => SumOutputs_2_20_port,
                           S(19) => SumOutputs_2_19_port, S(18) => 
                           SumOutputs_2_18_port, S(17) => SumOutputs_2_17_port,
                           S(16) => SumOutputs_2_16_port, S(15) => 
                           SumOutputs_2_15_port, S(14) => SumOutputs_2_14_port,
                           S(13) => SumOutputs_2_13_port, S(12) => 
                           SumOutputs_2_12_port, S(11) => SumOutputs_2_11_port,
                           S(10) => SumOutputs_2_10_port, S(9) => 
                           SumOutputs_2_9_port, S(8) => SumOutputs_2_8_port, 
                           S(7) => SumOutputs_2_7_port, S(6) => 
                           SumOutputs_2_6_port, S(5) => SumOutputs_2_5_port, 
                           S(4) => SumOutputs_2_4_port, S(3) => 
                           SumOutputs_2_3_port, S(2) => SumOutputs_2_2_port, 
                           S(1) => SumOutputs_2_1_port, S(0) => 
                           SumOutputs_2_0_port, Co => n_1129);
   SUMI_3 : RCA_NbitRca64_28 port map( A(63) => MuxOutputs_4_63_port, A(62) => 
                           MuxOutputs_4_62_port, A(61) => MuxOutputs_4_61_port,
                           A(60) => MuxOutputs_4_60_port, A(59) => 
                           MuxOutputs_4_59_port, A(58) => MuxOutputs_4_58_port,
                           A(57) => MuxOutputs_4_57_port, A(56) => 
                           MuxOutputs_4_56_port, A(55) => MuxOutputs_4_55_port,
                           A(54) => MuxOutputs_4_54_port, A(53) => 
                           MuxOutputs_4_53_port, A(52) => MuxOutputs_4_52_port,
                           A(51) => MuxOutputs_4_51_port, A(50) => 
                           MuxOutputs_4_50_port, A(49) => MuxOutputs_4_49_port,
                           A(48) => MuxOutputs_4_48_port, A(47) => 
                           MuxOutputs_4_47_port, A(46) => MuxOutputs_4_46_port,
                           A(45) => MuxOutputs_4_45_port, A(44) => 
                           MuxOutputs_4_44_port, A(43) => MuxOutputs_4_43_port,
                           A(42) => MuxOutputs_4_42_port, A(41) => 
                           MuxOutputs_4_41_port, A(40) => MuxOutputs_4_40_port,
                           A(39) => MuxOutputs_4_39_port, A(38) => 
                           MuxOutputs_4_38_port, A(37) => MuxOutputs_4_37_port,
                           A(36) => MuxOutputs_4_36_port, A(35) => 
                           MuxOutputs_4_35_port, A(34) => MuxOutputs_4_34_port,
                           A(33) => MuxOutputs_4_33_port, A(32) => 
                           MuxOutputs_4_32_port, A(31) => MuxOutputs_4_31_port,
                           A(30) => MuxOutputs_4_30_port, A(29) => 
                           MuxOutputs_4_29_port, A(28) => MuxOutputs_4_28_port,
                           A(27) => MuxOutputs_4_27_port, A(26) => 
                           MuxOutputs_4_26_port, A(25) => MuxOutputs_4_25_port,
                           A(24) => MuxOutputs_4_24_port, A(23) => 
                           MuxOutputs_4_23_port, A(22) => MuxOutputs_4_22_port,
                           A(21) => MuxOutputs_4_21_port, A(20) => 
                           MuxOutputs_4_20_port, A(19) => MuxOutputs_4_19_port,
                           A(18) => MuxOutputs_4_18_port, A(17) => 
                           MuxOutputs_4_17_port, A(16) => MuxOutputs_4_16_port,
                           A(15) => MuxOutputs_4_15_port, A(14) => 
                           MuxOutputs_4_14_port, A(13) => MuxOutputs_4_13_port,
                           A(12) => MuxOutputs_4_12_port, A(11) => 
                           MuxOutputs_4_11_port, A(10) => MuxOutputs_4_10_port,
                           A(9) => MuxOutputs_4_9_port, A(8) => 
                           MuxOutputs_4_8_port, A(7) => MuxOutputs_4_7_port, 
                           A(6) => MuxOutputs_4_6_port, A(5) => 
                           MuxOutputs_4_5_port, A(4) => MuxOutputs_4_4_port, 
                           A(3) => MuxOutputs_4_3_port, A(2) => 
                           MuxOutputs_4_2_port, A(1) => MuxOutputs_4_1_port, 
                           A(0) => MuxOutputs_4_0_port, B(63) => 
                           SumOutputs_2_63_port, B(62) => SumOutputs_2_62_port,
                           B(61) => SumOutputs_2_61_port, B(60) => 
                           SumOutputs_2_60_port, B(59) => SumOutputs_2_59_port,
                           B(58) => SumOutputs_2_58_port, B(57) => 
                           SumOutputs_2_57_port, B(56) => SumOutputs_2_56_port,
                           B(55) => SumOutputs_2_55_port, B(54) => 
                           SumOutputs_2_54_port, B(53) => SumOutputs_2_53_port,
                           B(52) => SumOutputs_2_52_port, B(51) => 
                           SumOutputs_2_51_port, B(50) => SumOutputs_2_50_port,
                           B(49) => SumOutputs_2_49_port, B(48) => 
                           SumOutputs_2_48_port, B(47) => SumOutputs_2_47_port,
                           B(46) => SumOutputs_2_46_port, B(45) => 
                           SumOutputs_2_45_port, B(44) => SumOutputs_2_44_port,
                           B(43) => SumOutputs_2_43_port, B(42) => 
                           SumOutputs_2_42_port, B(41) => SumOutputs_2_41_port,
                           B(40) => SumOutputs_2_40_port, B(39) => 
                           SumOutputs_2_39_port, B(38) => SumOutputs_2_38_port,
                           B(37) => SumOutputs_2_37_port, B(36) => 
                           SumOutputs_2_36_port, B(35) => SumOutputs_2_35_port,
                           B(34) => SumOutputs_2_34_port, B(33) => 
                           SumOutputs_2_33_port, B(32) => SumOutputs_2_32_port,
                           B(31) => SumOutputs_2_31_port, B(30) => 
                           SumOutputs_2_30_port, B(29) => SumOutputs_2_29_port,
                           B(28) => SumOutputs_2_28_port, B(27) => 
                           SumOutputs_2_27_port, B(26) => SumOutputs_2_26_port,
                           B(25) => SumOutputs_2_25_port, B(24) => 
                           SumOutputs_2_24_port, B(23) => SumOutputs_2_23_port,
                           B(22) => SumOutputs_2_22_port, B(21) => 
                           SumOutputs_2_21_port, B(20) => SumOutputs_2_20_port,
                           B(19) => SumOutputs_2_19_port, B(18) => 
                           SumOutputs_2_18_port, B(17) => SumOutputs_2_17_port,
                           B(16) => SumOutputs_2_16_port, B(15) => 
                           SumOutputs_2_15_port, B(14) => SumOutputs_2_14_port,
                           B(13) => SumOutputs_2_13_port, B(12) => 
                           SumOutputs_2_12_port, B(11) => SumOutputs_2_11_port,
                           B(10) => SumOutputs_2_10_port, B(9) => 
                           SumOutputs_2_9_port, B(8) => SumOutputs_2_8_port, 
                           B(7) => SumOutputs_2_7_port, B(6) => 
                           SumOutputs_2_6_port, B(5) => SumOutputs_2_5_port, 
                           B(4) => SumOutputs_2_4_port, B(3) => 
                           SumOutputs_2_3_port, B(2) => SumOutputs_2_2_port, 
                           B(1) => SumOutputs_2_1_port, B(0) => 
                           SumOutputs_2_0_port, Ci => X_Logic0_port, S(63) => 
                           SumOutputs_3_63_port, S(62) => SumOutputs_3_62_port,
                           S(61) => SumOutputs_3_61_port, S(60) => 
                           SumOutputs_3_60_port, S(59) => SumOutputs_3_59_port,
                           S(58) => SumOutputs_3_58_port, S(57) => 
                           SumOutputs_3_57_port, S(56) => SumOutputs_3_56_port,
                           S(55) => SumOutputs_3_55_port, S(54) => 
                           SumOutputs_3_54_port, S(53) => SumOutputs_3_53_port,
                           S(52) => SumOutputs_3_52_port, S(51) => 
                           SumOutputs_3_51_port, S(50) => SumOutputs_3_50_port,
                           S(49) => SumOutputs_3_49_port, S(48) => 
                           SumOutputs_3_48_port, S(47) => SumOutputs_3_47_port,
                           S(46) => SumOutputs_3_46_port, S(45) => 
                           SumOutputs_3_45_port, S(44) => SumOutputs_3_44_port,
                           S(43) => SumOutputs_3_43_port, S(42) => 
                           SumOutputs_3_42_port, S(41) => SumOutputs_3_41_port,
                           S(40) => SumOutputs_3_40_port, S(39) => 
                           SumOutputs_3_39_port, S(38) => SumOutputs_3_38_port,
                           S(37) => SumOutputs_3_37_port, S(36) => 
                           SumOutputs_3_36_port, S(35) => SumOutputs_3_35_port,
                           S(34) => SumOutputs_3_34_port, S(33) => 
                           SumOutputs_3_33_port, S(32) => SumOutputs_3_32_port,
                           S(31) => SumOutputs_3_31_port, S(30) => 
                           SumOutputs_3_30_port, S(29) => SumOutputs_3_29_port,
                           S(28) => SumOutputs_3_28_port, S(27) => 
                           SumOutputs_3_27_port, S(26) => SumOutputs_3_26_port,
                           S(25) => SumOutputs_3_25_port, S(24) => 
                           SumOutputs_3_24_port, S(23) => SumOutputs_3_23_port,
                           S(22) => SumOutputs_3_22_port, S(21) => 
                           SumOutputs_3_21_port, S(20) => SumOutputs_3_20_port,
                           S(19) => SumOutputs_3_19_port, S(18) => 
                           SumOutputs_3_18_port, S(17) => SumOutputs_3_17_port,
                           S(16) => SumOutputs_3_16_port, S(15) => 
                           SumOutputs_3_15_port, S(14) => SumOutputs_3_14_port,
                           S(13) => SumOutputs_3_13_port, S(12) => 
                           SumOutputs_3_12_port, S(11) => SumOutputs_3_11_port,
                           S(10) => SumOutputs_3_10_port, S(9) => 
                           SumOutputs_3_9_port, S(8) => SumOutputs_3_8_port, 
                           S(7) => SumOutputs_3_7_port, S(6) => 
                           SumOutputs_3_6_port, S(5) => SumOutputs_3_5_port, 
                           S(4) => SumOutputs_3_4_port, S(3) => 
                           SumOutputs_3_3_port, S(2) => SumOutputs_3_2_port, 
                           S(1) => SumOutputs_3_1_port, S(0) => 
                           SumOutputs_3_0_port, Co => n_1130);
   SUMI_4 : RCA_NbitRca64_27 port map( A(63) => MuxOutputs_5_63_port, A(62) => 
                           MuxOutputs_5_62_port, A(61) => MuxOutputs_5_61_port,
                           A(60) => MuxOutputs_5_60_port, A(59) => 
                           MuxOutputs_5_59_port, A(58) => MuxOutputs_5_58_port,
                           A(57) => MuxOutputs_5_57_port, A(56) => 
                           MuxOutputs_5_56_port, A(55) => MuxOutputs_5_55_port,
                           A(54) => MuxOutputs_5_54_port, A(53) => 
                           MuxOutputs_5_53_port, A(52) => MuxOutputs_5_52_port,
                           A(51) => MuxOutputs_5_51_port, A(50) => 
                           MuxOutputs_5_50_port, A(49) => MuxOutputs_5_49_port,
                           A(48) => MuxOutputs_5_48_port, A(47) => 
                           MuxOutputs_5_47_port, A(46) => MuxOutputs_5_46_port,
                           A(45) => MuxOutputs_5_45_port, A(44) => 
                           MuxOutputs_5_44_port, A(43) => MuxOutputs_5_43_port,
                           A(42) => MuxOutputs_5_42_port, A(41) => 
                           MuxOutputs_5_41_port, A(40) => MuxOutputs_5_40_port,
                           A(39) => MuxOutputs_5_39_port, A(38) => 
                           MuxOutputs_5_38_port, A(37) => MuxOutputs_5_37_port,
                           A(36) => MuxOutputs_5_36_port, A(35) => 
                           MuxOutputs_5_35_port, A(34) => MuxOutputs_5_34_port,
                           A(33) => MuxOutputs_5_33_port, A(32) => 
                           MuxOutputs_5_32_port, A(31) => MuxOutputs_5_31_port,
                           A(30) => MuxOutputs_5_30_port, A(29) => 
                           MuxOutputs_5_29_port, A(28) => MuxOutputs_5_28_port,
                           A(27) => MuxOutputs_5_27_port, A(26) => 
                           MuxOutputs_5_26_port, A(25) => MuxOutputs_5_25_port,
                           A(24) => MuxOutputs_5_24_port, A(23) => 
                           MuxOutputs_5_23_port, A(22) => MuxOutputs_5_22_port,
                           A(21) => MuxOutputs_5_21_port, A(20) => 
                           MuxOutputs_5_20_port, A(19) => MuxOutputs_5_19_port,
                           A(18) => MuxOutputs_5_18_port, A(17) => 
                           MuxOutputs_5_17_port, A(16) => MuxOutputs_5_16_port,
                           A(15) => MuxOutputs_5_15_port, A(14) => 
                           MuxOutputs_5_14_port, A(13) => MuxOutputs_5_13_port,
                           A(12) => MuxOutputs_5_12_port, A(11) => 
                           MuxOutputs_5_11_port, A(10) => MuxOutputs_5_10_port,
                           A(9) => MuxOutputs_5_9_port, A(8) => 
                           MuxOutputs_5_8_port, A(7) => MuxOutputs_5_7_port, 
                           A(6) => MuxOutputs_5_6_port, A(5) => 
                           MuxOutputs_5_5_port, A(4) => MuxOutputs_5_4_port, 
                           A(3) => MuxOutputs_5_3_port, A(2) => 
                           MuxOutputs_5_2_port, A(1) => MuxOutputs_5_1_port, 
                           A(0) => MuxOutputs_5_0_port, B(63) => 
                           SumOutputs_3_63_port, B(62) => SumOutputs_3_62_port,
                           B(61) => SumOutputs_3_61_port, B(60) => 
                           SumOutputs_3_60_port, B(59) => SumOutputs_3_59_port,
                           B(58) => SumOutputs_3_58_port, B(57) => 
                           SumOutputs_3_57_port, B(56) => SumOutputs_3_56_port,
                           B(55) => SumOutputs_3_55_port, B(54) => 
                           SumOutputs_3_54_port, B(53) => SumOutputs_3_53_port,
                           B(52) => SumOutputs_3_52_port, B(51) => 
                           SumOutputs_3_51_port, B(50) => SumOutputs_3_50_port,
                           B(49) => SumOutputs_3_49_port, B(48) => 
                           SumOutputs_3_48_port, B(47) => SumOutputs_3_47_port,
                           B(46) => SumOutputs_3_46_port, B(45) => 
                           SumOutputs_3_45_port, B(44) => SumOutputs_3_44_port,
                           B(43) => SumOutputs_3_43_port, B(42) => 
                           SumOutputs_3_42_port, B(41) => SumOutputs_3_41_port,
                           B(40) => SumOutputs_3_40_port, B(39) => 
                           SumOutputs_3_39_port, B(38) => SumOutputs_3_38_port,
                           B(37) => SumOutputs_3_37_port, B(36) => 
                           SumOutputs_3_36_port, B(35) => SumOutputs_3_35_port,
                           B(34) => SumOutputs_3_34_port, B(33) => 
                           SumOutputs_3_33_port, B(32) => SumOutputs_3_32_port,
                           B(31) => SumOutputs_3_31_port, B(30) => 
                           SumOutputs_3_30_port, B(29) => SumOutputs_3_29_port,
                           B(28) => SumOutputs_3_28_port, B(27) => 
                           SumOutputs_3_27_port, B(26) => SumOutputs_3_26_port,
                           B(25) => SumOutputs_3_25_port, B(24) => 
                           SumOutputs_3_24_port, B(23) => SumOutputs_3_23_port,
                           B(22) => SumOutputs_3_22_port, B(21) => 
                           SumOutputs_3_21_port, B(20) => SumOutputs_3_20_port,
                           B(19) => SumOutputs_3_19_port, B(18) => 
                           SumOutputs_3_18_port, B(17) => SumOutputs_3_17_port,
                           B(16) => SumOutputs_3_16_port, B(15) => 
                           SumOutputs_3_15_port, B(14) => SumOutputs_3_14_port,
                           B(13) => SumOutputs_3_13_port, B(12) => 
                           SumOutputs_3_12_port, B(11) => SumOutputs_3_11_port,
                           B(10) => SumOutputs_3_10_port, B(9) => 
                           SumOutputs_3_9_port, B(8) => SumOutputs_3_8_port, 
                           B(7) => SumOutputs_3_7_port, B(6) => 
                           SumOutputs_3_6_port, B(5) => SumOutputs_3_5_port, 
                           B(4) => SumOutputs_3_4_port, B(3) => 
                           SumOutputs_3_3_port, B(2) => SumOutputs_3_2_port, 
                           B(1) => SumOutputs_3_1_port, B(0) => 
                           SumOutputs_3_0_port, Ci => X_Logic0_port, S(63) => 
                           SumOutputs_4_63_port, S(62) => SumOutputs_4_62_port,
                           S(61) => SumOutputs_4_61_port, S(60) => 
                           SumOutputs_4_60_port, S(59) => SumOutputs_4_59_port,
                           S(58) => SumOutputs_4_58_port, S(57) => 
                           SumOutputs_4_57_port, S(56) => SumOutputs_4_56_port,
                           S(55) => SumOutputs_4_55_port, S(54) => 
                           SumOutputs_4_54_port, S(53) => SumOutputs_4_53_port,
                           S(52) => SumOutputs_4_52_port, S(51) => 
                           SumOutputs_4_51_port, S(50) => SumOutputs_4_50_port,
                           S(49) => SumOutputs_4_49_port, S(48) => 
                           SumOutputs_4_48_port, S(47) => SumOutputs_4_47_port,
                           S(46) => SumOutputs_4_46_port, S(45) => 
                           SumOutputs_4_45_port, S(44) => SumOutputs_4_44_port,
                           S(43) => SumOutputs_4_43_port, S(42) => 
                           SumOutputs_4_42_port, S(41) => SumOutputs_4_41_port,
                           S(40) => SumOutputs_4_40_port, S(39) => 
                           SumOutputs_4_39_port, S(38) => SumOutputs_4_38_port,
                           S(37) => SumOutputs_4_37_port, S(36) => 
                           SumOutputs_4_36_port, S(35) => SumOutputs_4_35_port,
                           S(34) => SumOutputs_4_34_port, S(33) => 
                           SumOutputs_4_33_port, S(32) => SumOutputs_4_32_port,
                           S(31) => SumOutputs_4_31_port, S(30) => 
                           SumOutputs_4_30_port, S(29) => SumOutputs_4_29_port,
                           S(28) => SumOutputs_4_28_port, S(27) => 
                           SumOutputs_4_27_port, S(26) => SumOutputs_4_26_port,
                           S(25) => SumOutputs_4_25_port, S(24) => 
                           SumOutputs_4_24_port, S(23) => SumOutputs_4_23_port,
                           S(22) => SumOutputs_4_22_port, S(21) => 
                           SumOutputs_4_21_port, S(20) => SumOutputs_4_20_port,
                           S(19) => SumOutputs_4_19_port, S(18) => 
                           SumOutputs_4_18_port, S(17) => SumOutputs_4_17_port,
                           S(16) => SumOutputs_4_16_port, S(15) => 
                           SumOutputs_4_15_port, S(14) => SumOutputs_4_14_port,
                           S(13) => SumOutputs_4_13_port, S(12) => 
                           SumOutputs_4_12_port, S(11) => SumOutputs_4_11_port,
                           S(10) => SumOutputs_4_10_port, S(9) => 
                           SumOutputs_4_9_port, S(8) => SumOutputs_4_8_port, 
                           S(7) => SumOutputs_4_7_port, S(6) => 
                           SumOutputs_4_6_port, S(5) => SumOutputs_4_5_port, 
                           S(4) => SumOutputs_4_4_port, S(3) => 
                           SumOutputs_4_3_port, S(2) => SumOutputs_4_2_port, 
                           S(1) => SumOutputs_4_1_port, S(0) => 
                           SumOutputs_4_0_port, Co => n_1131);
   SUMI_5 : RCA_NbitRca64_26 port map( A(63) => MuxOutputs_6_63_port, A(62) => 
                           MuxOutputs_6_62_port, A(61) => MuxOutputs_6_61_port,
                           A(60) => MuxOutputs_6_60_port, A(59) => 
                           MuxOutputs_6_59_port, A(58) => MuxOutputs_6_58_port,
                           A(57) => MuxOutputs_6_57_port, A(56) => 
                           MuxOutputs_6_56_port, A(55) => MuxOutputs_6_55_port,
                           A(54) => MuxOutputs_6_54_port, A(53) => 
                           MuxOutputs_6_53_port, A(52) => MuxOutputs_6_52_port,
                           A(51) => MuxOutputs_6_51_port, A(50) => 
                           MuxOutputs_6_50_port, A(49) => MuxOutputs_6_49_port,
                           A(48) => MuxOutputs_6_48_port, A(47) => 
                           MuxOutputs_6_47_port, A(46) => MuxOutputs_6_46_port,
                           A(45) => MuxOutputs_6_45_port, A(44) => 
                           MuxOutputs_6_44_port, A(43) => MuxOutputs_6_43_port,
                           A(42) => MuxOutputs_6_42_port, A(41) => 
                           MuxOutputs_6_41_port, A(40) => MuxOutputs_6_40_port,
                           A(39) => MuxOutputs_6_39_port, A(38) => 
                           MuxOutputs_6_38_port, A(37) => MuxOutputs_6_37_port,
                           A(36) => MuxOutputs_6_36_port, A(35) => 
                           MuxOutputs_6_35_port, A(34) => MuxOutputs_6_34_port,
                           A(33) => MuxOutputs_6_33_port, A(32) => 
                           MuxOutputs_6_32_port, A(31) => MuxOutputs_6_31_port,
                           A(30) => MuxOutputs_6_30_port, A(29) => 
                           MuxOutputs_6_29_port, A(28) => MuxOutputs_6_28_port,
                           A(27) => MuxOutputs_6_27_port, A(26) => 
                           MuxOutputs_6_26_port, A(25) => MuxOutputs_6_25_port,
                           A(24) => MuxOutputs_6_24_port, A(23) => 
                           MuxOutputs_6_23_port, A(22) => MuxOutputs_6_22_port,
                           A(21) => MuxOutputs_6_21_port, A(20) => 
                           MuxOutputs_6_20_port, A(19) => MuxOutputs_6_19_port,
                           A(18) => MuxOutputs_6_18_port, A(17) => 
                           MuxOutputs_6_17_port, A(16) => MuxOutputs_6_16_port,
                           A(15) => MuxOutputs_6_15_port, A(14) => 
                           MuxOutputs_6_14_port, A(13) => MuxOutputs_6_13_port,
                           A(12) => MuxOutputs_6_12_port, A(11) => 
                           MuxOutputs_6_11_port, A(10) => MuxOutputs_6_10_port,
                           A(9) => MuxOutputs_6_9_port, A(8) => 
                           MuxOutputs_6_8_port, A(7) => MuxOutputs_6_7_port, 
                           A(6) => MuxOutputs_6_6_port, A(5) => 
                           MuxOutputs_6_5_port, A(4) => MuxOutputs_6_4_port, 
                           A(3) => MuxOutputs_6_3_port, A(2) => 
                           MuxOutputs_6_2_port, A(1) => MuxOutputs_6_1_port, 
                           A(0) => MuxOutputs_6_0_port, B(63) => 
                           SumOutputs_4_63_port, B(62) => SumOutputs_4_62_port,
                           B(61) => SumOutputs_4_61_port, B(60) => 
                           SumOutputs_4_60_port, B(59) => SumOutputs_4_59_port,
                           B(58) => SumOutputs_4_58_port, B(57) => 
                           SumOutputs_4_57_port, B(56) => SumOutputs_4_56_port,
                           B(55) => SumOutputs_4_55_port, B(54) => 
                           SumOutputs_4_54_port, B(53) => SumOutputs_4_53_port,
                           B(52) => SumOutputs_4_52_port, B(51) => 
                           SumOutputs_4_51_port, B(50) => SumOutputs_4_50_port,
                           B(49) => SumOutputs_4_49_port, B(48) => 
                           SumOutputs_4_48_port, B(47) => SumOutputs_4_47_port,
                           B(46) => SumOutputs_4_46_port, B(45) => 
                           SumOutputs_4_45_port, B(44) => SumOutputs_4_44_port,
                           B(43) => SumOutputs_4_43_port, B(42) => 
                           SumOutputs_4_42_port, B(41) => SumOutputs_4_41_port,
                           B(40) => SumOutputs_4_40_port, B(39) => 
                           SumOutputs_4_39_port, B(38) => SumOutputs_4_38_port,
                           B(37) => SumOutputs_4_37_port, B(36) => 
                           SumOutputs_4_36_port, B(35) => SumOutputs_4_35_port,
                           B(34) => SumOutputs_4_34_port, B(33) => 
                           SumOutputs_4_33_port, B(32) => SumOutputs_4_32_port,
                           B(31) => SumOutputs_4_31_port, B(30) => 
                           SumOutputs_4_30_port, B(29) => SumOutputs_4_29_port,
                           B(28) => SumOutputs_4_28_port, B(27) => 
                           SumOutputs_4_27_port, B(26) => SumOutputs_4_26_port,
                           B(25) => SumOutputs_4_25_port, B(24) => 
                           SumOutputs_4_24_port, B(23) => SumOutputs_4_23_port,
                           B(22) => SumOutputs_4_22_port, B(21) => 
                           SumOutputs_4_21_port, B(20) => SumOutputs_4_20_port,
                           B(19) => SumOutputs_4_19_port, B(18) => 
                           SumOutputs_4_18_port, B(17) => SumOutputs_4_17_port,
                           B(16) => SumOutputs_4_16_port, B(15) => 
                           SumOutputs_4_15_port, B(14) => SumOutputs_4_14_port,
                           B(13) => SumOutputs_4_13_port, B(12) => 
                           SumOutputs_4_12_port, B(11) => SumOutputs_4_11_port,
                           B(10) => SumOutputs_4_10_port, B(9) => 
                           SumOutputs_4_9_port, B(8) => SumOutputs_4_8_port, 
                           B(7) => SumOutputs_4_7_port, B(6) => 
                           SumOutputs_4_6_port, B(5) => SumOutputs_4_5_port, 
                           B(4) => SumOutputs_4_4_port, B(3) => 
                           SumOutputs_4_3_port, B(2) => SumOutputs_4_2_port, 
                           B(1) => SumOutputs_4_1_port, B(0) => 
                           SumOutputs_4_0_port, Ci => X_Logic0_port, S(63) => 
                           SumOutputs_5_63_port, S(62) => SumOutputs_5_62_port,
                           S(61) => SumOutputs_5_61_port, S(60) => 
                           SumOutputs_5_60_port, S(59) => SumOutputs_5_59_port,
                           S(58) => SumOutputs_5_58_port, S(57) => 
                           SumOutputs_5_57_port, S(56) => SumOutputs_5_56_port,
                           S(55) => SumOutputs_5_55_port, S(54) => 
                           SumOutputs_5_54_port, S(53) => SumOutputs_5_53_port,
                           S(52) => SumOutputs_5_52_port, S(51) => 
                           SumOutputs_5_51_port, S(50) => SumOutputs_5_50_port,
                           S(49) => SumOutputs_5_49_port, S(48) => 
                           SumOutputs_5_48_port, S(47) => SumOutputs_5_47_port,
                           S(46) => SumOutputs_5_46_port, S(45) => 
                           SumOutputs_5_45_port, S(44) => SumOutputs_5_44_port,
                           S(43) => SumOutputs_5_43_port, S(42) => 
                           SumOutputs_5_42_port, S(41) => SumOutputs_5_41_port,
                           S(40) => SumOutputs_5_40_port, S(39) => 
                           SumOutputs_5_39_port, S(38) => SumOutputs_5_38_port,
                           S(37) => SumOutputs_5_37_port, S(36) => 
                           SumOutputs_5_36_port, S(35) => SumOutputs_5_35_port,
                           S(34) => SumOutputs_5_34_port, S(33) => 
                           SumOutputs_5_33_port, S(32) => SumOutputs_5_32_port,
                           S(31) => SumOutputs_5_31_port, S(30) => 
                           SumOutputs_5_30_port, S(29) => SumOutputs_5_29_port,
                           S(28) => SumOutputs_5_28_port, S(27) => 
                           SumOutputs_5_27_port, S(26) => SumOutputs_5_26_port,
                           S(25) => SumOutputs_5_25_port, S(24) => 
                           SumOutputs_5_24_port, S(23) => SumOutputs_5_23_port,
                           S(22) => SumOutputs_5_22_port, S(21) => 
                           SumOutputs_5_21_port, S(20) => SumOutputs_5_20_port,
                           S(19) => SumOutputs_5_19_port, S(18) => 
                           SumOutputs_5_18_port, S(17) => SumOutputs_5_17_port,
                           S(16) => SumOutputs_5_16_port, S(15) => 
                           SumOutputs_5_15_port, S(14) => SumOutputs_5_14_port,
                           S(13) => SumOutputs_5_13_port, S(12) => 
                           SumOutputs_5_12_port, S(11) => SumOutputs_5_11_port,
                           S(10) => SumOutputs_5_10_port, S(9) => 
                           SumOutputs_5_9_port, S(8) => SumOutputs_5_8_port, 
                           S(7) => SumOutputs_5_7_port, S(6) => 
                           SumOutputs_5_6_port, S(5) => SumOutputs_5_5_port, 
                           S(4) => SumOutputs_5_4_port, S(3) => 
                           SumOutputs_5_3_port, S(2) => SumOutputs_5_2_port, 
                           S(1) => SumOutputs_5_1_port, S(0) => 
                           SumOutputs_5_0_port, Co => n_1132);
   SUMI_6 : RCA_NbitRca64_25 port map( A(63) => MuxOutputs_7_63_port, A(62) => 
                           MuxOutputs_7_62_port, A(61) => MuxOutputs_7_61_port,
                           A(60) => MuxOutputs_7_60_port, A(59) => 
                           MuxOutputs_7_59_port, A(58) => MuxOutputs_7_58_port,
                           A(57) => MuxOutputs_7_57_port, A(56) => 
                           MuxOutputs_7_56_port, A(55) => MuxOutputs_7_55_port,
                           A(54) => MuxOutputs_7_54_port, A(53) => 
                           MuxOutputs_7_53_port, A(52) => MuxOutputs_7_52_port,
                           A(51) => MuxOutputs_7_51_port, A(50) => 
                           MuxOutputs_7_50_port, A(49) => MuxOutputs_7_49_port,
                           A(48) => MuxOutputs_7_48_port, A(47) => 
                           MuxOutputs_7_47_port, A(46) => MuxOutputs_7_46_port,
                           A(45) => MuxOutputs_7_45_port, A(44) => 
                           MuxOutputs_7_44_port, A(43) => MuxOutputs_7_43_port,
                           A(42) => MuxOutputs_7_42_port, A(41) => 
                           MuxOutputs_7_41_port, A(40) => MuxOutputs_7_40_port,
                           A(39) => MuxOutputs_7_39_port, A(38) => 
                           MuxOutputs_7_38_port, A(37) => MuxOutputs_7_37_port,
                           A(36) => MuxOutputs_7_36_port, A(35) => 
                           MuxOutputs_7_35_port, A(34) => MuxOutputs_7_34_port,
                           A(33) => MuxOutputs_7_33_port, A(32) => 
                           MuxOutputs_7_32_port, A(31) => MuxOutputs_7_31_port,
                           A(30) => MuxOutputs_7_30_port, A(29) => 
                           MuxOutputs_7_29_port, A(28) => MuxOutputs_7_28_port,
                           A(27) => MuxOutputs_7_27_port, A(26) => 
                           MuxOutputs_7_26_port, A(25) => MuxOutputs_7_25_port,
                           A(24) => MuxOutputs_7_24_port, A(23) => 
                           MuxOutputs_7_23_port, A(22) => MuxOutputs_7_22_port,
                           A(21) => MuxOutputs_7_21_port, A(20) => 
                           MuxOutputs_7_20_port, A(19) => MuxOutputs_7_19_port,
                           A(18) => MuxOutputs_7_18_port, A(17) => 
                           MuxOutputs_7_17_port, A(16) => MuxOutputs_7_16_port,
                           A(15) => MuxOutputs_7_15_port, A(14) => 
                           MuxOutputs_7_14_port, A(13) => MuxOutputs_7_13_port,
                           A(12) => MuxOutputs_7_12_port, A(11) => 
                           MuxOutputs_7_11_port, A(10) => MuxOutputs_7_10_port,
                           A(9) => MuxOutputs_7_9_port, A(8) => 
                           MuxOutputs_7_8_port, A(7) => MuxOutputs_7_7_port, 
                           A(6) => MuxOutputs_7_6_port, A(5) => 
                           MuxOutputs_7_5_port, A(4) => MuxOutputs_7_4_port, 
                           A(3) => MuxOutputs_7_3_port, A(2) => 
                           MuxOutputs_7_2_port, A(1) => MuxOutputs_7_1_port, 
                           A(0) => MuxOutputs_7_0_port, B(63) => 
                           SumOutputs_5_63_port, B(62) => SumOutputs_5_62_port,
                           B(61) => SumOutputs_5_61_port, B(60) => 
                           SumOutputs_5_60_port, B(59) => SumOutputs_5_59_port,
                           B(58) => SumOutputs_5_58_port, B(57) => 
                           SumOutputs_5_57_port, B(56) => SumOutputs_5_56_port,
                           B(55) => SumOutputs_5_55_port, B(54) => 
                           SumOutputs_5_54_port, B(53) => SumOutputs_5_53_port,
                           B(52) => SumOutputs_5_52_port, B(51) => 
                           SumOutputs_5_51_port, B(50) => SumOutputs_5_50_port,
                           B(49) => SumOutputs_5_49_port, B(48) => 
                           SumOutputs_5_48_port, B(47) => SumOutputs_5_47_port,
                           B(46) => SumOutputs_5_46_port, B(45) => 
                           SumOutputs_5_45_port, B(44) => SumOutputs_5_44_port,
                           B(43) => SumOutputs_5_43_port, B(42) => 
                           SumOutputs_5_42_port, B(41) => SumOutputs_5_41_port,
                           B(40) => SumOutputs_5_40_port, B(39) => 
                           SumOutputs_5_39_port, B(38) => SumOutputs_5_38_port,
                           B(37) => SumOutputs_5_37_port, B(36) => 
                           SumOutputs_5_36_port, B(35) => SumOutputs_5_35_port,
                           B(34) => SumOutputs_5_34_port, B(33) => 
                           SumOutputs_5_33_port, B(32) => SumOutputs_5_32_port,
                           B(31) => SumOutputs_5_31_port, B(30) => 
                           SumOutputs_5_30_port, B(29) => SumOutputs_5_29_port,
                           B(28) => SumOutputs_5_28_port, B(27) => 
                           SumOutputs_5_27_port, B(26) => SumOutputs_5_26_port,
                           B(25) => SumOutputs_5_25_port, B(24) => 
                           SumOutputs_5_24_port, B(23) => SumOutputs_5_23_port,
                           B(22) => SumOutputs_5_22_port, B(21) => 
                           SumOutputs_5_21_port, B(20) => SumOutputs_5_20_port,
                           B(19) => SumOutputs_5_19_port, B(18) => 
                           SumOutputs_5_18_port, B(17) => SumOutputs_5_17_port,
                           B(16) => SumOutputs_5_16_port, B(15) => 
                           SumOutputs_5_15_port, B(14) => SumOutputs_5_14_port,
                           B(13) => SumOutputs_5_13_port, B(12) => 
                           SumOutputs_5_12_port, B(11) => SumOutputs_5_11_port,
                           B(10) => SumOutputs_5_10_port, B(9) => 
                           SumOutputs_5_9_port, B(8) => SumOutputs_5_8_port, 
                           B(7) => SumOutputs_5_7_port, B(6) => 
                           SumOutputs_5_6_port, B(5) => SumOutputs_5_5_port, 
                           B(4) => SumOutputs_5_4_port, B(3) => 
                           SumOutputs_5_3_port, B(2) => SumOutputs_5_2_port, 
                           B(1) => SumOutputs_5_1_port, B(0) => 
                           SumOutputs_5_0_port, Ci => X_Logic0_port, S(63) => 
                           SumOutputs_6_63_port, S(62) => SumOutputs_6_62_port,
                           S(61) => SumOutputs_6_61_port, S(60) => 
                           SumOutputs_6_60_port, S(59) => SumOutputs_6_59_port,
                           S(58) => SumOutputs_6_58_port, S(57) => 
                           SumOutputs_6_57_port, S(56) => SumOutputs_6_56_port,
                           S(55) => SumOutputs_6_55_port, S(54) => 
                           SumOutputs_6_54_port, S(53) => SumOutputs_6_53_port,
                           S(52) => SumOutputs_6_52_port, S(51) => 
                           SumOutputs_6_51_port, S(50) => SumOutputs_6_50_port,
                           S(49) => SumOutputs_6_49_port, S(48) => 
                           SumOutputs_6_48_port, S(47) => SumOutputs_6_47_port,
                           S(46) => SumOutputs_6_46_port, S(45) => 
                           SumOutputs_6_45_port, S(44) => SumOutputs_6_44_port,
                           S(43) => SumOutputs_6_43_port, S(42) => 
                           SumOutputs_6_42_port, S(41) => SumOutputs_6_41_port,
                           S(40) => SumOutputs_6_40_port, S(39) => 
                           SumOutputs_6_39_port, S(38) => SumOutputs_6_38_port,
                           S(37) => SumOutputs_6_37_port, S(36) => 
                           SumOutputs_6_36_port, S(35) => SumOutputs_6_35_port,
                           S(34) => SumOutputs_6_34_port, S(33) => 
                           SumOutputs_6_33_port, S(32) => SumOutputs_6_32_port,
                           S(31) => SumOutputs_6_31_port, S(30) => 
                           SumOutputs_6_30_port, S(29) => SumOutputs_6_29_port,
                           S(28) => SumOutputs_6_28_port, S(27) => 
                           SumOutputs_6_27_port, S(26) => SumOutputs_6_26_port,
                           S(25) => SumOutputs_6_25_port, S(24) => 
                           SumOutputs_6_24_port, S(23) => SumOutputs_6_23_port,
                           S(22) => SumOutputs_6_22_port, S(21) => 
                           SumOutputs_6_21_port, S(20) => SumOutputs_6_20_port,
                           S(19) => SumOutputs_6_19_port, S(18) => 
                           SumOutputs_6_18_port, S(17) => SumOutputs_6_17_port,
                           S(16) => SumOutputs_6_16_port, S(15) => 
                           SumOutputs_6_15_port, S(14) => SumOutputs_6_14_port,
                           S(13) => SumOutputs_6_13_port, S(12) => 
                           SumOutputs_6_12_port, S(11) => SumOutputs_6_11_port,
                           S(10) => SumOutputs_6_10_port, S(9) => 
                           SumOutputs_6_9_port, S(8) => SumOutputs_6_8_port, 
                           S(7) => SumOutputs_6_7_port, S(6) => 
                           SumOutputs_6_6_port, S(5) => SumOutputs_6_5_port, 
                           S(4) => SumOutputs_6_4_port, S(3) => 
                           SumOutputs_6_3_port, S(2) => SumOutputs_6_2_port, 
                           S(1) => SumOutputs_6_1_port, S(0) => 
                           SumOutputs_6_0_port, Co => n_1133);
   SUMI_7 : RCA_NbitRca64_24 port map( A(63) => MuxOutputs_8_63_port, A(62) => 
                           MuxOutputs_8_62_port, A(61) => MuxOutputs_8_61_port,
                           A(60) => MuxOutputs_8_60_port, A(59) => 
                           MuxOutputs_8_59_port, A(58) => MuxOutputs_8_58_port,
                           A(57) => MuxOutputs_8_57_port, A(56) => 
                           MuxOutputs_8_56_port, A(55) => MuxOutputs_8_55_port,
                           A(54) => MuxOutputs_8_54_port, A(53) => 
                           MuxOutputs_8_53_port, A(52) => MuxOutputs_8_52_port,
                           A(51) => MuxOutputs_8_51_port, A(50) => 
                           MuxOutputs_8_50_port, A(49) => MuxOutputs_8_49_port,
                           A(48) => MuxOutputs_8_48_port, A(47) => 
                           MuxOutputs_8_47_port, A(46) => MuxOutputs_8_46_port,
                           A(45) => MuxOutputs_8_45_port, A(44) => 
                           MuxOutputs_8_44_port, A(43) => MuxOutputs_8_43_port,
                           A(42) => MuxOutputs_8_42_port, A(41) => 
                           MuxOutputs_8_41_port, A(40) => MuxOutputs_8_40_port,
                           A(39) => MuxOutputs_8_39_port, A(38) => 
                           MuxOutputs_8_38_port, A(37) => MuxOutputs_8_37_port,
                           A(36) => MuxOutputs_8_36_port, A(35) => 
                           MuxOutputs_8_35_port, A(34) => MuxOutputs_8_34_port,
                           A(33) => MuxOutputs_8_33_port, A(32) => 
                           MuxOutputs_8_32_port, A(31) => MuxOutputs_8_31_port,
                           A(30) => MuxOutputs_8_30_port, A(29) => 
                           MuxOutputs_8_29_port, A(28) => MuxOutputs_8_28_port,
                           A(27) => MuxOutputs_8_27_port, A(26) => 
                           MuxOutputs_8_26_port, A(25) => MuxOutputs_8_25_port,
                           A(24) => MuxOutputs_8_24_port, A(23) => 
                           MuxOutputs_8_23_port, A(22) => MuxOutputs_8_22_port,
                           A(21) => MuxOutputs_8_21_port, A(20) => 
                           MuxOutputs_8_20_port, A(19) => MuxOutputs_8_19_port,
                           A(18) => MuxOutputs_8_18_port, A(17) => 
                           MuxOutputs_8_17_port, A(16) => MuxOutputs_8_16_port,
                           A(15) => MuxOutputs_8_15_port, A(14) => 
                           MuxOutputs_8_14_port, A(13) => MuxOutputs_8_13_port,
                           A(12) => MuxOutputs_8_12_port, A(11) => 
                           MuxOutputs_8_11_port, A(10) => MuxOutputs_8_10_port,
                           A(9) => MuxOutputs_8_9_port, A(8) => 
                           MuxOutputs_8_8_port, A(7) => MuxOutputs_8_7_port, 
                           A(6) => MuxOutputs_8_6_port, A(5) => 
                           MuxOutputs_8_5_port, A(4) => MuxOutputs_8_4_port, 
                           A(3) => MuxOutputs_8_3_port, A(2) => 
                           MuxOutputs_8_2_port, A(1) => MuxOutputs_8_1_port, 
                           A(0) => MuxOutputs_8_0_port, B(63) => 
                           SumOutputs_6_63_port, B(62) => SumOutputs_6_62_port,
                           B(61) => SumOutputs_6_61_port, B(60) => 
                           SumOutputs_6_60_port, B(59) => SumOutputs_6_59_port,
                           B(58) => SumOutputs_6_58_port, B(57) => 
                           SumOutputs_6_57_port, B(56) => SumOutputs_6_56_port,
                           B(55) => SumOutputs_6_55_port, B(54) => 
                           SumOutputs_6_54_port, B(53) => SumOutputs_6_53_port,
                           B(52) => SumOutputs_6_52_port, B(51) => 
                           SumOutputs_6_51_port, B(50) => SumOutputs_6_50_port,
                           B(49) => SumOutputs_6_49_port, B(48) => 
                           SumOutputs_6_48_port, B(47) => SumOutputs_6_47_port,
                           B(46) => SumOutputs_6_46_port, B(45) => 
                           SumOutputs_6_45_port, B(44) => SumOutputs_6_44_port,
                           B(43) => SumOutputs_6_43_port, B(42) => 
                           SumOutputs_6_42_port, B(41) => SumOutputs_6_41_port,
                           B(40) => SumOutputs_6_40_port, B(39) => 
                           SumOutputs_6_39_port, B(38) => SumOutputs_6_38_port,
                           B(37) => SumOutputs_6_37_port, B(36) => 
                           SumOutputs_6_36_port, B(35) => SumOutputs_6_35_port,
                           B(34) => SumOutputs_6_34_port, B(33) => 
                           SumOutputs_6_33_port, B(32) => SumOutputs_6_32_port,
                           B(31) => SumOutputs_6_31_port, B(30) => 
                           SumOutputs_6_30_port, B(29) => SumOutputs_6_29_port,
                           B(28) => SumOutputs_6_28_port, B(27) => 
                           SumOutputs_6_27_port, B(26) => SumOutputs_6_26_port,
                           B(25) => SumOutputs_6_25_port, B(24) => 
                           SumOutputs_6_24_port, B(23) => SumOutputs_6_23_port,
                           B(22) => SumOutputs_6_22_port, B(21) => 
                           SumOutputs_6_21_port, B(20) => SumOutputs_6_20_port,
                           B(19) => SumOutputs_6_19_port, B(18) => 
                           SumOutputs_6_18_port, B(17) => SumOutputs_6_17_port,
                           B(16) => SumOutputs_6_16_port, B(15) => 
                           SumOutputs_6_15_port, B(14) => SumOutputs_6_14_port,
                           B(13) => SumOutputs_6_13_port, B(12) => 
                           SumOutputs_6_12_port, B(11) => SumOutputs_6_11_port,
                           B(10) => SumOutputs_6_10_port, B(9) => 
                           SumOutputs_6_9_port, B(8) => SumOutputs_6_8_port, 
                           B(7) => SumOutputs_6_7_port, B(6) => 
                           SumOutputs_6_6_port, B(5) => SumOutputs_6_5_port, 
                           B(4) => SumOutputs_6_4_port, B(3) => 
                           SumOutputs_6_3_port, B(2) => SumOutputs_6_2_port, 
                           B(1) => SumOutputs_6_1_port, B(0) => 
                           SumOutputs_6_0_port, Ci => X_Logic0_port, S(63) => 
                           SumOutputs_7_63_port, S(62) => SumOutputs_7_62_port,
                           S(61) => SumOutputs_7_61_port, S(60) => 
                           SumOutputs_7_60_port, S(59) => SumOutputs_7_59_port,
                           S(58) => SumOutputs_7_58_port, S(57) => 
                           SumOutputs_7_57_port, S(56) => SumOutputs_7_56_port,
                           S(55) => SumOutputs_7_55_port, S(54) => 
                           SumOutputs_7_54_port, S(53) => SumOutputs_7_53_port,
                           S(52) => SumOutputs_7_52_port, S(51) => 
                           SumOutputs_7_51_port, S(50) => SumOutputs_7_50_port,
                           S(49) => SumOutputs_7_49_port, S(48) => 
                           SumOutputs_7_48_port, S(47) => SumOutputs_7_47_port,
                           S(46) => SumOutputs_7_46_port, S(45) => 
                           SumOutputs_7_45_port, S(44) => SumOutputs_7_44_port,
                           S(43) => SumOutputs_7_43_port, S(42) => 
                           SumOutputs_7_42_port, S(41) => SumOutputs_7_41_port,
                           S(40) => SumOutputs_7_40_port, S(39) => 
                           SumOutputs_7_39_port, S(38) => SumOutputs_7_38_port,
                           S(37) => SumOutputs_7_37_port, S(36) => 
                           SumOutputs_7_36_port, S(35) => SumOutputs_7_35_port,
                           S(34) => SumOutputs_7_34_port, S(33) => 
                           SumOutputs_7_33_port, S(32) => SumOutputs_7_32_port,
                           S(31) => SumOutputs_7_31_port, S(30) => 
                           SumOutputs_7_30_port, S(29) => SumOutputs_7_29_port,
                           S(28) => SumOutputs_7_28_port, S(27) => 
                           SumOutputs_7_27_port, S(26) => SumOutputs_7_26_port,
                           S(25) => SumOutputs_7_25_port, S(24) => 
                           SumOutputs_7_24_port, S(23) => SumOutputs_7_23_port,
                           S(22) => SumOutputs_7_22_port, S(21) => 
                           SumOutputs_7_21_port, S(20) => SumOutputs_7_20_port,
                           S(19) => SumOutputs_7_19_port, S(18) => 
                           SumOutputs_7_18_port, S(17) => SumOutputs_7_17_port,
                           S(16) => SumOutputs_7_16_port, S(15) => 
                           SumOutputs_7_15_port, S(14) => SumOutputs_7_14_port,
                           S(13) => SumOutputs_7_13_port, S(12) => 
                           SumOutputs_7_12_port, S(11) => SumOutputs_7_11_port,
                           S(10) => SumOutputs_7_10_port, S(9) => 
                           SumOutputs_7_9_port, S(8) => SumOutputs_7_8_port, 
                           S(7) => SumOutputs_7_7_port, S(6) => 
                           SumOutputs_7_6_port, S(5) => SumOutputs_7_5_port, 
                           S(4) => SumOutputs_7_4_port, S(3) => 
                           SumOutputs_7_3_port, S(2) => SumOutputs_7_2_port, 
                           S(1) => SumOutputs_7_1_port, S(0) => 
                           SumOutputs_7_0_port, Co => n_1134);
   SUMI_8 : RCA_NbitRca64_23 port map( A(63) => MuxOutputs_9_63_port, A(62) => 
                           MuxOutputs_9_62_port, A(61) => MuxOutputs_9_61_port,
                           A(60) => MuxOutputs_9_60_port, A(59) => 
                           MuxOutputs_9_59_port, A(58) => MuxOutputs_9_58_port,
                           A(57) => MuxOutputs_9_57_port, A(56) => 
                           MuxOutputs_9_56_port, A(55) => MuxOutputs_9_55_port,
                           A(54) => MuxOutputs_9_54_port, A(53) => 
                           MuxOutputs_9_53_port, A(52) => MuxOutputs_9_52_port,
                           A(51) => MuxOutputs_9_51_port, A(50) => 
                           MuxOutputs_9_50_port, A(49) => MuxOutputs_9_49_port,
                           A(48) => MuxOutputs_9_48_port, A(47) => 
                           MuxOutputs_9_47_port, A(46) => MuxOutputs_9_46_port,
                           A(45) => MuxOutputs_9_45_port, A(44) => 
                           MuxOutputs_9_44_port, A(43) => MuxOutputs_9_43_port,
                           A(42) => MuxOutputs_9_42_port, A(41) => 
                           MuxOutputs_9_41_port, A(40) => MuxOutputs_9_40_port,
                           A(39) => MuxOutputs_9_39_port, A(38) => 
                           MuxOutputs_9_38_port, A(37) => MuxOutputs_9_37_port,
                           A(36) => MuxOutputs_9_36_port, A(35) => 
                           MuxOutputs_9_35_port, A(34) => MuxOutputs_9_34_port,
                           A(33) => MuxOutputs_9_33_port, A(32) => 
                           MuxOutputs_9_32_port, A(31) => MuxOutputs_9_31_port,
                           A(30) => MuxOutputs_9_30_port, A(29) => 
                           MuxOutputs_9_29_port, A(28) => MuxOutputs_9_28_port,
                           A(27) => MuxOutputs_9_27_port, A(26) => 
                           MuxOutputs_9_26_port, A(25) => MuxOutputs_9_25_port,
                           A(24) => MuxOutputs_9_24_port, A(23) => 
                           MuxOutputs_9_23_port, A(22) => MuxOutputs_9_22_port,
                           A(21) => MuxOutputs_9_21_port, A(20) => 
                           MuxOutputs_9_20_port, A(19) => MuxOutputs_9_19_port,
                           A(18) => MuxOutputs_9_18_port, A(17) => 
                           MuxOutputs_9_17_port, A(16) => MuxOutputs_9_16_port,
                           A(15) => MuxOutputs_9_15_port, A(14) => 
                           MuxOutputs_9_14_port, A(13) => MuxOutputs_9_13_port,
                           A(12) => MuxOutputs_9_12_port, A(11) => 
                           MuxOutputs_9_11_port, A(10) => MuxOutputs_9_10_port,
                           A(9) => MuxOutputs_9_9_port, A(8) => 
                           MuxOutputs_9_8_port, A(7) => MuxOutputs_9_7_port, 
                           A(6) => MuxOutputs_9_6_port, A(5) => 
                           MuxOutputs_9_5_port, A(4) => MuxOutputs_9_4_port, 
                           A(3) => MuxOutputs_9_3_port, A(2) => 
                           MuxOutputs_9_2_port, A(1) => MuxOutputs_9_1_port, 
                           A(0) => MuxOutputs_9_0_port, B(63) => 
                           SumOutputs_7_63_port, B(62) => SumOutputs_7_62_port,
                           B(61) => SumOutputs_7_61_port, B(60) => 
                           SumOutputs_7_60_port, B(59) => SumOutputs_7_59_port,
                           B(58) => SumOutputs_7_58_port, B(57) => 
                           SumOutputs_7_57_port, B(56) => SumOutputs_7_56_port,
                           B(55) => SumOutputs_7_55_port, B(54) => 
                           SumOutputs_7_54_port, B(53) => SumOutputs_7_53_port,
                           B(52) => SumOutputs_7_52_port, B(51) => 
                           SumOutputs_7_51_port, B(50) => SumOutputs_7_50_port,
                           B(49) => SumOutputs_7_49_port, B(48) => 
                           SumOutputs_7_48_port, B(47) => SumOutputs_7_47_port,
                           B(46) => SumOutputs_7_46_port, B(45) => 
                           SumOutputs_7_45_port, B(44) => SumOutputs_7_44_port,
                           B(43) => SumOutputs_7_43_port, B(42) => 
                           SumOutputs_7_42_port, B(41) => SumOutputs_7_41_port,
                           B(40) => SumOutputs_7_40_port, B(39) => 
                           SumOutputs_7_39_port, B(38) => SumOutputs_7_38_port,
                           B(37) => SumOutputs_7_37_port, B(36) => 
                           SumOutputs_7_36_port, B(35) => SumOutputs_7_35_port,
                           B(34) => SumOutputs_7_34_port, B(33) => 
                           SumOutputs_7_33_port, B(32) => SumOutputs_7_32_port,
                           B(31) => SumOutputs_7_31_port, B(30) => 
                           SumOutputs_7_30_port, B(29) => SumOutputs_7_29_port,
                           B(28) => SumOutputs_7_28_port, B(27) => 
                           SumOutputs_7_27_port, B(26) => SumOutputs_7_26_port,
                           B(25) => SumOutputs_7_25_port, B(24) => 
                           SumOutputs_7_24_port, B(23) => SumOutputs_7_23_port,
                           B(22) => SumOutputs_7_22_port, B(21) => 
                           SumOutputs_7_21_port, B(20) => SumOutputs_7_20_port,
                           B(19) => SumOutputs_7_19_port, B(18) => 
                           SumOutputs_7_18_port, B(17) => SumOutputs_7_17_port,
                           B(16) => SumOutputs_7_16_port, B(15) => 
                           SumOutputs_7_15_port, B(14) => SumOutputs_7_14_port,
                           B(13) => SumOutputs_7_13_port, B(12) => 
                           SumOutputs_7_12_port, B(11) => SumOutputs_7_11_port,
                           B(10) => SumOutputs_7_10_port, B(9) => 
                           SumOutputs_7_9_port, B(8) => SumOutputs_7_8_port, 
                           B(7) => SumOutputs_7_7_port, B(6) => 
                           SumOutputs_7_6_port, B(5) => SumOutputs_7_5_port, 
                           B(4) => SumOutputs_7_4_port, B(3) => 
                           SumOutputs_7_3_port, B(2) => SumOutputs_7_2_port, 
                           B(1) => SumOutputs_7_1_port, B(0) => 
                           SumOutputs_7_0_port, Ci => X_Logic0_port, S(63) => 
                           SumOutputs_8_63_port, S(62) => SumOutputs_8_62_port,
                           S(61) => SumOutputs_8_61_port, S(60) => 
                           SumOutputs_8_60_port, S(59) => SumOutputs_8_59_port,
                           S(58) => SumOutputs_8_58_port, S(57) => 
                           SumOutputs_8_57_port, S(56) => SumOutputs_8_56_port,
                           S(55) => SumOutputs_8_55_port, S(54) => 
                           SumOutputs_8_54_port, S(53) => SumOutputs_8_53_port,
                           S(52) => SumOutputs_8_52_port, S(51) => 
                           SumOutputs_8_51_port, S(50) => SumOutputs_8_50_port,
                           S(49) => SumOutputs_8_49_port, S(48) => 
                           SumOutputs_8_48_port, S(47) => SumOutputs_8_47_port,
                           S(46) => SumOutputs_8_46_port, S(45) => 
                           SumOutputs_8_45_port, S(44) => SumOutputs_8_44_port,
                           S(43) => SumOutputs_8_43_port, S(42) => 
                           SumOutputs_8_42_port, S(41) => SumOutputs_8_41_port,
                           S(40) => SumOutputs_8_40_port, S(39) => 
                           SumOutputs_8_39_port, S(38) => SumOutputs_8_38_port,
                           S(37) => SumOutputs_8_37_port, S(36) => 
                           SumOutputs_8_36_port, S(35) => SumOutputs_8_35_port,
                           S(34) => SumOutputs_8_34_port, S(33) => 
                           SumOutputs_8_33_port, S(32) => SumOutputs_8_32_port,
                           S(31) => SumOutputs_8_31_port, S(30) => 
                           SumOutputs_8_30_port, S(29) => SumOutputs_8_29_port,
                           S(28) => SumOutputs_8_28_port, S(27) => 
                           SumOutputs_8_27_port, S(26) => SumOutputs_8_26_port,
                           S(25) => SumOutputs_8_25_port, S(24) => 
                           SumOutputs_8_24_port, S(23) => SumOutputs_8_23_port,
                           S(22) => SumOutputs_8_22_port, S(21) => 
                           SumOutputs_8_21_port, S(20) => SumOutputs_8_20_port,
                           S(19) => SumOutputs_8_19_port, S(18) => 
                           SumOutputs_8_18_port, S(17) => SumOutputs_8_17_port,
                           S(16) => SumOutputs_8_16_port, S(15) => 
                           SumOutputs_8_15_port, S(14) => SumOutputs_8_14_port,
                           S(13) => SumOutputs_8_13_port, S(12) => 
                           SumOutputs_8_12_port, S(11) => SumOutputs_8_11_port,
                           S(10) => SumOutputs_8_10_port, S(9) => 
                           SumOutputs_8_9_port, S(8) => SumOutputs_8_8_port, 
                           S(7) => SumOutputs_8_7_port, S(6) => 
                           SumOutputs_8_6_port, S(5) => SumOutputs_8_5_port, 
                           S(4) => SumOutputs_8_4_port, S(3) => 
                           SumOutputs_8_3_port, S(2) => SumOutputs_8_2_port, 
                           S(1) => SumOutputs_8_1_port, S(0) => 
                           SumOutputs_8_0_port, Co => n_1135);
   SUMI_9 : RCA_NbitRca64_22 port map( A(63) => MuxOutputs_10_63_port, A(62) =>
                           MuxOutputs_10_62_port, A(61) => 
                           MuxOutputs_10_61_port, A(60) => 
                           MuxOutputs_10_60_port, A(59) => 
                           MuxOutputs_10_59_port, A(58) => 
                           MuxOutputs_10_58_port, A(57) => 
                           MuxOutputs_10_57_port, A(56) => 
                           MuxOutputs_10_56_port, A(55) => 
                           MuxOutputs_10_55_port, A(54) => 
                           MuxOutputs_10_54_port, A(53) => 
                           MuxOutputs_10_53_port, A(52) => 
                           MuxOutputs_10_52_port, A(51) => 
                           MuxOutputs_10_51_port, A(50) => 
                           MuxOutputs_10_50_port, A(49) => 
                           MuxOutputs_10_49_port, A(48) => 
                           MuxOutputs_10_48_port, A(47) => 
                           MuxOutputs_10_47_port, A(46) => 
                           MuxOutputs_10_46_port, A(45) => 
                           MuxOutputs_10_45_port, A(44) => 
                           MuxOutputs_10_44_port, A(43) => 
                           MuxOutputs_10_43_port, A(42) => 
                           MuxOutputs_10_42_port, A(41) => 
                           MuxOutputs_10_41_port, A(40) => 
                           MuxOutputs_10_40_port, A(39) => 
                           MuxOutputs_10_39_port, A(38) => 
                           MuxOutputs_10_38_port, A(37) => 
                           MuxOutputs_10_37_port, A(36) => 
                           MuxOutputs_10_36_port, A(35) => 
                           MuxOutputs_10_35_port, A(34) => 
                           MuxOutputs_10_34_port, A(33) => 
                           MuxOutputs_10_33_port, A(32) => 
                           MuxOutputs_10_32_port, A(31) => 
                           MuxOutputs_10_31_port, A(30) => 
                           MuxOutputs_10_30_port, A(29) => 
                           MuxOutputs_10_29_port, A(28) => 
                           MuxOutputs_10_28_port, A(27) => 
                           MuxOutputs_10_27_port, A(26) => 
                           MuxOutputs_10_26_port, A(25) => 
                           MuxOutputs_10_25_port, A(24) => 
                           MuxOutputs_10_24_port, A(23) => 
                           MuxOutputs_10_23_port, A(22) => 
                           MuxOutputs_10_22_port, A(21) => 
                           MuxOutputs_10_21_port, A(20) => 
                           MuxOutputs_10_20_port, A(19) => 
                           MuxOutputs_10_19_port, A(18) => 
                           MuxOutputs_10_18_port, A(17) => 
                           MuxOutputs_10_17_port, A(16) => 
                           MuxOutputs_10_16_port, A(15) => 
                           MuxOutputs_10_15_port, A(14) => 
                           MuxOutputs_10_14_port, A(13) => 
                           MuxOutputs_10_13_port, A(12) => 
                           MuxOutputs_10_12_port, A(11) => 
                           MuxOutputs_10_11_port, A(10) => 
                           MuxOutputs_10_10_port, A(9) => MuxOutputs_10_9_port,
                           A(8) => MuxOutputs_10_8_port, A(7) => 
                           MuxOutputs_10_7_port, A(6) => MuxOutputs_10_6_port, 
                           A(5) => MuxOutputs_10_5_port, A(4) => 
                           MuxOutputs_10_4_port, A(3) => MuxOutputs_10_3_port, 
                           A(2) => MuxOutputs_10_2_port, A(1) => 
                           MuxOutputs_10_1_port, A(0) => MuxOutputs_10_0_port, 
                           B(63) => SumOutputs_8_63_port, B(62) => 
                           SumOutputs_8_62_port, B(61) => SumOutputs_8_61_port,
                           B(60) => SumOutputs_8_60_port, B(59) => 
                           SumOutputs_8_59_port, B(58) => SumOutputs_8_58_port,
                           B(57) => SumOutputs_8_57_port, B(56) => 
                           SumOutputs_8_56_port, B(55) => SumOutputs_8_55_port,
                           B(54) => SumOutputs_8_54_port, B(53) => 
                           SumOutputs_8_53_port, B(52) => SumOutputs_8_52_port,
                           B(51) => SumOutputs_8_51_port, B(50) => 
                           SumOutputs_8_50_port, B(49) => SumOutputs_8_49_port,
                           B(48) => SumOutputs_8_48_port, B(47) => 
                           SumOutputs_8_47_port, B(46) => SumOutputs_8_46_port,
                           B(45) => SumOutputs_8_45_port, B(44) => 
                           SumOutputs_8_44_port, B(43) => SumOutputs_8_43_port,
                           B(42) => SumOutputs_8_42_port, B(41) => 
                           SumOutputs_8_41_port, B(40) => SumOutputs_8_40_port,
                           B(39) => SumOutputs_8_39_port, B(38) => 
                           SumOutputs_8_38_port, B(37) => SumOutputs_8_37_port,
                           B(36) => SumOutputs_8_36_port, B(35) => 
                           SumOutputs_8_35_port, B(34) => SumOutputs_8_34_port,
                           B(33) => SumOutputs_8_33_port, B(32) => 
                           SumOutputs_8_32_port, B(31) => SumOutputs_8_31_port,
                           B(30) => SumOutputs_8_30_port, B(29) => 
                           SumOutputs_8_29_port, B(28) => SumOutputs_8_28_port,
                           B(27) => SumOutputs_8_27_port, B(26) => 
                           SumOutputs_8_26_port, B(25) => SumOutputs_8_25_port,
                           B(24) => SumOutputs_8_24_port, B(23) => 
                           SumOutputs_8_23_port, B(22) => SumOutputs_8_22_port,
                           B(21) => SumOutputs_8_21_port, B(20) => 
                           SumOutputs_8_20_port, B(19) => SumOutputs_8_19_port,
                           B(18) => SumOutputs_8_18_port, B(17) => 
                           SumOutputs_8_17_port, B(16) => SumOutputs_8_16_port,
                           B(15) => SumOutputs_8_15_port, B(14) => 
                           SumOutputs_8_14_port, B(13) => SumOutputs_8_13_port,
                           B(12) => SumOutputs_8_12_port, B(11) => 
                           SumOutputs_8_11_port, B(10) => SumOutputs_8_10_port,
                           B(9) => SumOutputs_8_9_port, B(8) => 
                           SumOutputs_8_8_port, B(7) => SumOutputs_8_7_port, 
                           B(6) => SumOutputs_8_6_port, B(5) => 
                           SumOutputs_8_5_port, B(4) => SumOutputs_8_4_port, 
                           B(3) => SumOutputs_8_3_port, B(2) => 
                           SumOutputs_8_2_port, B(1) => SumOutputs_8_1_port, 
                           B(0) => SumOutputs_8_0_port, Ci => X_Logic0_port, 
                           S(63) => SumOutputs_9_63_port, S(62) => 
                           SumOutputs_9_62_port, S(61) => SumOutputs_9_61_port,
                           S(60) => SumOutputs_9_60_port, S(59) => 
                           SumOutputs_9_59_port, S(58) => SumOutputs_9_58_port,
                           S(57) => SumOutputs_9_57_port, S(56) => 
                           SumOutputs_9_56_port, S(55) => SumOutputs_9_55_port,
                           S(54) => SumOutputs_9_54_port, S(53) => 
                           SumOutputs_9_53_port, S(52) => SumOutputs_9_52_port,
                           S(51) => SumOutputs_9_51_port, S(50) => 
                           SumOutputs_9_50_port, S(49) => SumOutputs_9_49_port,
                           S(48) => SumOutputs_9_48_port, S(47) => 
                           SumOutputs_9_47_port, S(46) => SumOutputs_9_46_port,
                           S(45) => SumOutputs_9_45_port, S(44) => 
                           SumOutputs_9_44_port, S(43) => SumOutputs_9_43_port,
                           S(42) => SumOutputs_9_42_port, S(41) => 
                           SumOutputs_9_41_port, S(40) => SumOutputs_9_40_port,
                           S(39) => SumOutputs_9_39_port, S(38) => 
                           SumOutputs_9_38_port, S(37) => SumOutputs_9_37_port,
                           S(36) => SumOutputs_9_36_port, S(35) => 
                           SumOutputs_9_35_port, S(34) => SumOutputs_9_34_port,
                           S(33) => SumOutputs_9_33_port, S(32) => 
                           SumOutputs_9_32_port, S(31) => SumOutputs_9_31_port,
                           S(30) => SumOutputs_9_30_port, S(29) => 
                           SumOutputs_9_29_port, S(28) => SumOutputs_9_28_port,
                           S(27) => SumOutputs_9_27_port, S(26) => 
                           SumOutputs_9_26_port, S(25) => SumOutputs_9_25_port,
                           S(24) => SumOutputs_9_24_port, S(23) => 
                           SumOutputs_9_23_port, S(22) => SumOutputs_9_22_port,
                           S(21) => SumOutputs_9_21_port, S(20) => 
                           SumOutputs_9_20_port, S(19) => SumOutputs_9_19_port,
                           S(18) => SumOutputs_9_18_port, S(17) => 
                           SumOutputs_9_17_port, S(16) => SumOutputs_9_16_port,
                           S(15) => SumOutputs_9_15_port, S(14) => 
                           SumOutputs_9_14_port, S(13) => SumOutputs_9_13_port,
                           S(12) => SumOutputs_9_12_port, S(11) => 
                           SumOutputs_9_11_port, S(10) => SumOutputs_9_10_port,
                           S(9) => SumOutputs_9_9_port, S(8) => 
                           SumOutputs_9_8_port, S(7) => SumOutputs_9_7_port, 
                           S(6) => SumOutputs_9_6_port, S(5) => 
                           SumOutputs_9_5_port, S(4) => SumOutputs_9_4_port, 
                           S(3) => SumOutputs_9_3_port, S(2) => 
                           SumOutputs_9_2_port, S(1) => SumOutputs_9_1_port, 
                           S(0) => SumOutputs_9_0_port, Co => n_1136);
   SUMI_10 : RCA_NbitRca64_21 port map( A(63) => MuxOutputs_11_63_port, A(62) 
                           => MuxOutputs_11_62_port, A(61) => 
                           MuxOutputs_11_61_port, A(60) => 
                           MuxOutputs_11_60_port, A(59) => 
                           MuxOutputs_11_59_port, A(58) => 
                           MuxOutputs_11_58_port, A(57) => 
                           MuxOutputs_11_57_port, A(56) => 
                           MuxOutputs_11_56_port, A(55) => 
                           MuxOutputs_11_55_port, A(54) => 
                           MuxOutputs_11_54_port, A(53) => 
                           MuxOutputs_11_53_port, A(52) => 
                           MuxOutputs_11_52_port, A(51) => 
                           MuxOutputs_11_51_port, A(50) => 
                           MuxOutputs_11_50_port, A(49) => 
                           MuxOutputs_11_49_port, A(48) => 
                           MuxOutputs_11_48_port, A(47) => 
                           MuxOutputs_11_47_port, A(46) => 
                           MuxOutputs_11_46_port, A(45) => 
                           MuxOutputs_11_45_port, A(44) => 
                           MuxOutputs_11_44_port, A(43) => 
                           MuxOutputs_11_43_port, A(42) => 
                           MuxOutputs_11_42_port, A(41) => 
                           MuxOutputs_11_41_port, A(40) => 
                           MuxOutputs_11_40_port, A(39) => 
                           MuxOutputs_11_39_port, A(38) => 
                           MuxOutputs_11_38_port, A(37) => 
                           MuxOutputs_11_37_port, A(36) => 
                           MuxOutputs_11_36_port, A(35) => 
                           MuxOutputs_11_35_port, A(34) => 
                           MuxOutputs_11_34_port, A(33) => 
                           MuxOutputs_11_33_port, A(32) => 
                           MuxOutputs_11_32_port, A(31) => 
                           MuxOutputs_11_31_port, A(30) => 
                           MuxOutputs_11_30_port, A(29) => 
                           MuxOutputs_11_29_port, A(28) => 
                           MuxOutputs_11_28_port, A(27) => 
                           MuxOutputs_11_27_port, A(26) => 
                           MuxOutputs_11_26_port, A(25) => 
                           MuxOutputs_11_25_port, A(24) => 
                           MuxOutputs_11_24_port, A(23) => 
                           MuxOutputs_11_23_port, A(22) => 
                           MuxOutputs_11_22_port, A(21) => 
                           MuxOutputs_11_21_port, A(20) => 
                           MuxOutputs_11_20_port, A(19) => 
                           MuxOutputs_11_19_port, A(18) => 
                           MuxOutputs_11_18_port, A(17) => 
                           MuxOutputs_11_17_port, A(16) => 
                           MuxOutputs_11_16_port, A(15) => 
                           MuxOutputs_11_15_port, A(14) => 
                           MuxOutputs_11_14_port, A(13) => 
                           MuxOutputs_11_13_port, A(12) => 
                           MuxOutputs_11_12_port, A(11) => 
                           MuxOutputs_11_11_port, A(10) => 
                           MuxOutputs_11_10_port, A(9) => MuxOutputs_11_9_port,
                           A(8) => MuxOutputs_11_8_port, A(7) => 
                           MuxOutputs_11_7_port, A(6) => MuxOutputs_11_6_port, 
                           A(5) => MuxOutputs_11_5_port, A(4) => 
                           MuxOutputs_11_4_port, A(3) => MuxOutputs_11_3_port, 
                           A(2) => MuxOutputs_11_2_port, A(1) => 
                           MuxOutputs_11_1_port, A(0) => MuxOutputs_11_0_port, 
                           B(63) => SumOutputs_9_63_port, B(62) => 
                           SumOutputs_9_62_port, B(61) => SumOutputs_9_61_port,
                           B(60) => SumOutputs_9_60_port, B(59) => 
                           SumOutputs_9_59_port, B(58) => SumOutputs_9_58_port,
                           B(57) => SumOutputs_9_57_port, B(56) => 
                           SumOutputs_9_56_port, B(55) => SumOutputs_9_55_port,
                           B(54) => SumOutputs_9_54_port, B(53) => 
                           SumOutputs_9_53_port, B(52) => SumOutputs_9_52_port,
                           B(51) => SumOutputs_9_51_port, B(50) => 
                           SumOutputs_9_50_port, B(49) => SumOutputs_9_49_port,
                           B(48) => SumOutputs_9_48_port, B(47) => 
                           SumOutputs_9_47_port, B(46) => SumOutputs_9_46_port,
                           B(45) => SumOutputs_9_45_port, B(44) => 
                           SumOutputs_9_44_port, B(43) => SumOutputs_9_43_port,
                           B(42) => SumOutputs_9_42_port, B(41) => 
                           SumOutputs_9_41_port, B(40) => SumOutputs_9_40_port,
                           B(39) => SumOutputs_9_39_port, B(38) => 
                           SumOutputs_9_38_port, B(37) => SumOutputs_9_37_port,
                           B(36) => SumOutputs_9_36_port, B(35) => 
                           SumOutputs_9_35_port, B(34) => SumOutputs_9_34_port,
                           B(33) => SumOutputs_9_33_port, B(32) => 
                           SumOutputs_9_32_port, B(31) => SumOutputs_9_31_port,
                           B(30) => SumOutputs_9_30_port, B(29) => 
                           SumOutputs_9_29_port, B(28) => SumOutputs_9_28_port,
                           B(27) => SumOutputs_9_27_port, B(26) => 
                           SumOutputs_9_26_port, B(25) => SumOutputs_9_25_port,
                           B(24) => SumOutputs_9_24_port, B(23) => 
                           SumOutputs_9_23_port, B(22) => SumOutputs_9_22_port,
                           B(21) => SumOutputs_9_21_port, B(20) => 
                           SumOutputs_9_20_port, B(19) => SumOutputs_9_19_port,
                           B(18) => SumOutputs_9_18_port, B(17) => 
                           SumOutputs_9_17_port, B(16) => SumOutputs_9_16_port,
                           B(15) => SumOutputs_9_15_port, B(14) => 
                           SumOutputs_9_14_port, B(13) => SumOutputs_9_13_port,
                           B(12) => SumOutputs_9_12_port, B(11) => 
                           SumOutputs_9_11_port, B(10) => SumOutputs_9_10_port,
                           B(9) => SumOutputs_9_9_port, B(8) => 
                           SumOutputs_9_8_port, B(7) => SumOutputs_9_7_port, 
                           B(6) => SumOutputs_9_6_port, B(5) => 
                           SumOutputs_9_5_port, B(4) => SumOutputs_9_4_port, 
                           B(3) => SumOutputs_9_3_port, B(2) => 
                           SumOutputs_9_2_port, B(1) => SumOutputs_9_1_port, 
                           B(0) => SumOutputs_9_0_port, Ci => X_Logic0_port, 
                           S(63) => SumOutputs_10_63_port, S(62) => 
                           SumOutputs_10_62_port, S(61) => 
                           SumOutputs_10_61_port, S(60) => 
                           SumOutputs_10_60_port, S(59) => 
                           SumOutputs_10_59_port, S(58) => 
                           SumOutputs_10_58_port, S(57) => 
                           SumOutputs_10_57_port, S(56) => 
                           SumOutputs_10_56_port, S(55) => 
                           SumOutputs_10_55_port, S(54) => 
                           SumOutputs_10_54_port, S(53) => 
                           SumOutputs_10_53_port, S(52) => 
                           SumOutputs_10_52_port, S(51) => 
                           SumOutputs_10_51_port, S(50) => 
                           SumOutputs_10_50_port, S(49) => 
                           SumOutputs_10_49_port, S(48) => 
                           SumOutputs_10_48_port, S(47) => 
                           SumOutputs_10_47_port, S(46) => 
                           SumOutputs_10_46_port, S(45) => 
                           SumOutputs_10_45_port, S(44) => 
                           SumOutputs_10_44_port, S(43) => 
                           SumOutputs_10_43_port, S(42) => 
                           SumOutputs_10_42_port, S(41) => 
                           SumOutputs_10_41_port, S(40) => 
                           SumOutputs_10_40_port, S(39) => 
                           SumOutputs_10_39_port, S(38) => 
                           SumOutputs_10_38_port, S(37) => 
                           SumOutputs_10_37_port, S(36) => 
                           SumOutputs_10_36_port, S(35) => 
                           SumOutputs_10_35_port, S(34) => 
                           SumOutputs_10_34_port, S(33) => 
                           SumOutputs_10_33_port, S(32) => 
                           SumOutputs_10_32_port, S(31) => 
                           SumOutputs_10_31_port, S(30) => 
                           SumOutputs_10_30_port, S(29) => 
                           SumOutputs_10_29_port, S(28) => 
                           SumOutputs_10_28_port, S(27) => 
                           SumOutputs_10_27_port, S(26) => 
                           SumOutputs_10_26_port, S(25) => 
                           SumOutputs_10_25_port, S(24) => 
                           SumOutputs_10_24_port, S(23) => 
                           SumOutputs_10_23_port, S(22) => 
                           SumOutputs_10_22_port, S(21) => 
                           SumOutputs_10_21_port, S(20) => 
                           SumOutputs_10_20_port, S(19) => 
                           SumOutputs_10_19_port, S(18) => 
                           SumOutputs_10_18_port, S(17) => 
                           SumOutputs_10_17_port, S(16) => 
                           SumOutputs_10_16_port, S(15) => 
                           SumOutputs_10_15_port, S(14) => 
                           SumOutputs_10_14_port, S(13) => 
                           SumOutputs_10_13_port, S(12) => 
                           SumOutputs_10_12_port, S(11) => 
                           SumOutputs_10_11_port, S(10) => 
                           SumOutputs_10_10_port, S(9) => SumOutputs_10_9_port,
                           S(8) => SumOutputs_10_8_port, S(7) => 
                           SumOutputs_10_7_port, S(6) => SumOutputs_10_6_port, 
                           S(5) => SumOutputs_10_5_port, S(4) => 
                           SumOutputs_10_4_port, S(3) => SumOutputs_10_3_port, 
                           S(2) => SumOutputs_10_2_port, S(1) => 
                           SumOutputs_10_1_port, S(0) => SumOutputs_10_0_port, 
                           Co => n_1137);
   SUMI_11 : RCA_NbitRca64_20 port map( A(63) => MuxOutputs_12_63_port, A(62) 
                           => MuxOutputs_12_62_port, A(61) => 
                           MuxOutputs_12_61_port, A(60) => 
                           MuxOutputs_12_60_port, A(59) => 
                           MuxOutputs_12_59_port, A(58) => 
                           MuxOutputs_12_58_port, A(57) => 
                           MuxOutputs_12_57_port, A(56) => 
                           MuxOutputs_12_56_port, A(55) => 
                           MuxOutputs_12_55_port, A(54) => 
                           MuxOutputs_12_54_port, A(53) => 
                           MuxOutputs_12_53_port, A(52) => 
                           MuxOutputs_12_52_port, A(51) => 
                           MuxOutputs_12_51_port, A(50) => 
                           MuxOutputs_12_50_port, A(49) => 
                           MuxOutputs_12_49_port, A(48) => 
                           MuxOutputs_12_48_port, A(47) => 
                           MuxOutputs_12_47_port, A(46) => 
                           MuxOutputs_12_46_port, A(45) => 
                           MuxOutputs_12_45_port, A(44) => 
                           MuxOutputs_12_44_port, A(43) => 
                           MuxOutputs_12_43_port, A(42) => 
                           MuxOutputs_12_42_port, A(41) => 
                           MuxOutputs_12_41_port, A(40) => 
                           MuxOutputs_12_40_port, A(39) => 
                           MuxOutputs_12_39_port, A(38) => 
                           MuxOutputs_12_38_port, A(37) => 
                           MuxOutputs_12_37_port, A(36) => 
                           MuxOutputs_12_36_port, A(35) => 
                           MuxOutputs_12_35_port, A(34) => 
                           MuxOutputs_12_34_port, A(33) => 
                           MuxOutputs_12_33_port, A(32) => 
                           MuxOutputs_12_32_port, A(31) => 
                           MuxOutputs_12_31_port, A(30) => 
                           MuxOutputs_12_30_port, A(29) => 
                           MuxOutputs_12_29_port, A(28) => 
                           MuxOutputs_12_28_port, A(27) => 
                           MuxOutputs_12_27_port, A(26) => 
                           MuxOutputs_12_26_port, A(25) => 
                           MuxOutputs_12_25_port, A(24) => 
                           MuxOutputs_12_24_port, A(23) => 
                           MuxOutputs_12_23_port, A(22) => 
                           MuxOutputs_12_22_port, A(21) => 
                           MuxOutputs_12_21_port, A(20) => 
                           MuxOutputs_12_20_port, A(19) => 
                           MuxOutputs_12_19_port, A(18) => 
                           MuxOutputs_12_18_port, A(17) => 
                           MuxOutputs_12_17_port, A(16) => 
                           MuxOutputs_12_16_port, A(15) => 
                           MuxOutputs_12_15_port, A(14) => 
                           MuxOutputs_12_14_port, A(13) => 
                           MuxOutputs_12_13_port, A(12) => 
                           MuxOutputs_12_12_port, A(11) => 
                           MuxOutputs_12_11_port, A(10) => 
                           MuxOutputs_12_10_port, A(9) => MuxOutputs_12_9_port,
                           A(8) => MuxOutputs_12_8_port, A(7) => 
                           MuxOutputs_12_7_port, A(6) => MuxOutputs_12_6_port, 
                           A(5) => MuxOutputs_12_5_port, A(4) => 
                           MuxOutputs_12_4_port, A(3) => MuxOutputs_12_3_port, 
                           A(2) => MuxOutputs_12_2_port, A(1) => 
                           MuxOutputs_12_1_port, A(0) => MuxOutputs_12_0_port, 
                           B(63) => SumOutputs_10_63_port, B(62) => 
                           SumOutputs_10_62_port, B(61) => 
                           SumOutputs_10_61_port, B(60) => 
                           SumOutputs_10_60_port, B(59) => 
                           SumOutputs_10_59_port, B(58) => 
                           SumOutputs_10_58_port, B(57) => 
                           SumOutputs_10_57_port, B(56) => 
                           SumOutputs_10_56_port, B(55) => 
                           SumOutputs_10_55_port, B(54) => 
                           SumOutputs_10_54_port, B(53) => 
                           SumOutputs_10_53_port, B(52) => 
                           SumOutputs_10_52_port, B(51) => 
                           SumOutputs_10_51_port, B(50) => 
                           SumOutputs_10_50_port, B(49) => 
                           SumOutputs_10_49_port, B(48) => 
                           SumOutputs_10_48_port, B(47) => 
                           SumOutputs_10_47_port, B(46) => 
                           SumOutputs_10_46_port, B(45) => 
                           SumOutputs_10_45_port, B(44) => 
                           SumOutputs_10_44_port, B(43) => 
                           SumOutputs_10_43_port, B(42) => 
                           SumOutputs_10_42_port, B(41) => 
                           SumOutputs_10_41_port, B(40) => 
                           SumOutputs_10_40_port, B(39) => 
                           SumOutputs_10_39_port, B(38) => 
                           SumOutputs_10_38_port, B(37) => 
                           SumOutputs_10_37_port, B(36) => 
                           SumOutputs_10_36_port, B(35) => 
                           SumOutputs_10_35_port, B(34) => 
                           SumOutputs_10_34_port, B(33) => 
                           SumOutputs_10_33_port, B(32) => 
                           SumOutputs_10_32_port, B(31) => 
                           SumOutputs_10_31_port, B(30) => 
                           SumOutputs_10_30_port, B(29) => 
                           SumOutputs_10_29_port, B(28) => 
                           SumOutputs_10_28_port, B(27) => 
                           SumOutputs_10_27_port, B(26) => 
                           SumOutputs_10_26_port, B(25) => 
                           SumOutputs_10_25_port, B(24) => 
                           SumOutputs_10_24_port, B(23) => 
                           SumOutputs_10_23_port, B(22) => 
                           SumOutputs_10_22_port, B(21) => 
                           SumOutputs_10_21_port, B(20) => 
                           SumOutputs_10_20_port, B(19) => 
                           SumOutputs_10_19_port, B(18) => 
                           SumOutputs_10_18_port, B(17) => 
                           SumOutputs_10_17_port, B(16) => 
                           SumOutputs_10_16_port, B(15) => 
                           SumOutputs_10_15_port, B(14) => 
                           SumOutputs_10_14_port, B(13) => 
                           SumOutputs_10_13_port, B(12) => 
                           SumOutputs_10_12_port, B(11) => 
                           SumOutputs_10_11_port, B(10) => 
                           SumOutputs_10_10_port, B(9) => SumOutputs_10_9_port,
                           B(8) => SumOutputs_10_8_port, B(7) => 
                           SumOutputs_10_7_port, B(6) => SumOutputs_10_6_port, 
                           B(5) => SumOutputs_10_5_port, B(4) => 
                           SumOutputs_10_4_port, B(3) => SumOutputs_10_3_port, 
                           B(2) => SumOutputs_10_2_port, B(1) => 
                           SumOutputs_10_1_port, B(0) => SumOutputs_10_0_port, 
                           Ci => X_Logic0_port, S(63) => SumOutputs_11_63_port,
                           S(62) => SumOutputs_11_62_port, S(61) => 
                           SumOutputs_11_61_port, S(60) => 
                           SumOutputs_11_60_port, S(59) => 
                           SumOutputs_11_59_port, S(58) => 
                           SumOutputs_11_58_port, S(57) => 
                           SumOutputs_11_57_port, S(56) => 
                           SumOutputs_11_56_port, S(55) => 
                           SumOutputs_11_55_port, S(54) => 
                           SumOutputs_11_54_port, S(53) => 
                           SumOutputs_11_53_port, S(52) => 
                           SumOutputs_11_52_port, S(51) => 
                           SumOutputs_11_51_port, S(50) => 
                           SumOutputs_11_50_port, S(49) => 
                           SumOutputs_11_49_port, S(48) => 
                           SumOutputs_11_48_port, S(47) => 
                           SumOutputs_11_47_port, S(46) => 
                           SumOutputs_11_46_port, S(45) => 
                           SumOutputs_11_45_port, S(44) => 
                           SumOutputs_11_44_port, S(43) => 
                           SumOutputs_11_43_port, S(42) => 
                           SumOutputs_11_42_port, S(41) => 
                           SumOutputs_11_41_port, S(40) => 
                           SumOutputs_11_40_port, S(39) => 
                           SumOutputs_11_39_port, S(38) => 
                           SumOutputs_11_38_port, S(37) => 
                           SumOutputs_11_37_port, S(36) => 
                           SumOutputs_11_36_port, S(35) => 
                           SumOutputs_11_35_port, S(34) => 
                           SumOutputs_11_34_port, S(33) => 
                           SumOutputs_11_33_port, S(32) => 
                           SumOutputs_11_32_port, S(31) => 
                           SumOutputs_11_31_port, S(30) => 
                           SumOutputs_11_30_port, S(29) => 
                           SumOutputs_11_29_port, S(28) => 
                           SumOutputs_11_28_port, S(27) => 
                           SumOutputs_11_27_port, S(26) => 
                           SumOutputs_11_26_port, S(25) => 
                           SumOutputs_11_25_port, S(24) => 
                           SumOutputs_11_24_port, S(23) => 
                           SumOutputs_11_23_port, S(22) => 
                           SumOutputs_11_22_port, S(21) => 
                           SumOutputs_11_21_port, S(20) => 
                           SumOutputs_11_20_port, S(19) => 
                           SumOutputs_11_19_port, S(18) => 
                           SumOutputs_11_18_port, S(17) => 
                           SumOutputs_11_17_port, S(16) => 
                           SumOutputs_11_16_port, S(15) => 
                           SumOutputs_11_15_port, S(14) => 
                           SumOutputs_11_14_port, S(13) => 
                           SumOutputs_11_13_port, S(12) => 
                           SumOutputs_11_12_port, S(11) => 
                           SumOutputs_11_11_port, S(10) => 
                           SumOutputs_11_10_port, S(9) => SumOutputs_11_9_port,
                           S(8) => SumOutputs_11_8_port, S(7) => 
                           SumOutputs_11_7_port, S(6) => SumOutputs_11_6_port, 
                           S(5) => SumOutputs_11_5_port, S(4) => 
                           SumOutputs_11_4_port, S(3) => SumOutputs_11_3_port, 
                           S(2) => SumOutputs_11_2_port, S(1) => 
                           SumOutputs_11_1_port, S(0) => SumOutputs_11_0_port, 
                           Co => n_1138);
   SUMI_12 : RCA_NbitRca64_19 port map( A(63) => MuxOutputs_13_63_port, A(62) 
                           => MuxOutputs_13_62_port, A(61) => 
                           MuxOutputs_13_61_port, A(60) => 
                           MuxOutputs_13_60_port, A(59) => 
                           MuxOutputs_13_59_port, A(58) => 
                           MuxOutputs_13_58_port, A(57) => 
                           MuxOutputs_13_57_port, A(56) => 
                           MuxOutputs_13_56_port, A(55) => 
                           MuxOutputs_13_55_port, A(54) => 
                           MuxOutputs_13_54_port, A(53) => 
                           MuxOutputs_13_53_port, A(52) => 
                           MuxOutputs_13_52_port, A(51) => 
                           MuxOutputs_13_51_port, A(50) => 
                           MuxOutputs_13_50_port, A(49) => 
                           MuxOutputs_13_49_port, A(48) => 
                           MuxOutputs_13_48_port, A(47) => 
                           MuxOutputs_13_47_port, A(46) => 
                           MuxOutputs_13_46_port, A(45) => 
                           MuxOutputs_13_45_port, A(44) => 
                           MuxOutputs_13_44_port, A(43) => 
                           MuxOutputs_13_43_port, A(42) => 
                           MuxOutputs_13_42_port, A(41) => 
                           MuxOutputs_13_41_port, A(40) => 
                           MuxOutputs_13_40_port, A(39) => 
                           MuxOutputs_13_39_port, A(38) => 
                           MuxOutputs_13_38_port, A(37) => 
                           MuxOutputs_13_37_port, A(36) => 
                           MuxOutputs_13_36_port, A(35) => 
                           MuxOutputs_13_35_port, A(34) => 
                           MuxOutputs_13_34_port, A(33) => 
                           MuxOutputs_13_33_port, A(32) => 
                           MuxOutputs_13_32_port, A(31) => 
                           MuxOutputs_13_31_port, A(30) => 
                           MuxOutputs_13_30_port, A(29) => 
                           MuxOutputs_13_29_port, A(28) => 
                           MuxOutputs_13_28_port, A(27) => 
                           MuxOutputs_13_27_port, A(26) => 
                           MuxOutputs_13_26_port, A(25) => 
                           MuxOutputs_13_25_port, A(24) => 
                           MuxOutputs_13_24_port, A(23) => 
                           MuxOutputs_13_23_port, A(22) => 
                           MuxOutputs_13_22_port, A(21) => 
                           MuxOutputs_13_21_port, A(20) => 
                           MuxOutputs_13_20_port, A(19) => 
                           MuxOutputs_13_19_port, A(18) => 
                           MuxOutputs_13_18_port, A(17) => 
                           MuxOutputs_13_17_port, A(16) => 
                           MuxOutputs_13_16_port, A(15) => 
                           MuxOutputs_13_15_port, A(14) => 
                           MuxOutputs_13_14_port, A(13) => 
                           MuxOutputs_13_13_port, A(12) => 
                           MuxOutputs_13_12_port, A(11) => 
                           MuxOutputs_13_11_port, A(10) => 
                           MuxOutputs_13_10_port, A(9) => MuxOutputs_13_9_port,
                           A(8) => MuxOutputs_13_8_port, A(7) => 
                           MuxOutputs_13_7_port, A(6) => MuxOutputs_13_6_port, 
                           A(5) => MuxOutputs_13_5_port, A(4) => 
                           MuxOutputs_13_4_port, A(3) => MuxOutputs_13_3_port, 
                           A(2) => MuxOutputs_13_2_port, A(1) => 
                           MuxOutputs_13_1_port, A(0) => MuxOutputs_13_0_port, 
                           B(63) => SumOutputs_11_63_port, B(62) => 
                           SumOutputs_11_62_port, B(61) => 
                           SumOutputs_11_61_port, B(60) => 
                           SumOutputs_11_60_port, B(59) => 
                           SumOutputs_11_59_port, B(58) => 
                           SumOutputs_11_58_port, B(57) => 
                           SumOutputs_11_57_port, B(56) => 
                           SumOutputs_11_56_port, B(55) => 
                           SumOutputs_11_55_port, B(54) => 
                           SumOutputs_11_54_port, B(53) => 
                           SumOutputs_11_53_port, B(52) => 
                           SumOutputs_11_52_port, B(51) => 
                           SumOutputs_11_51_port, B(50) => 
                           SumOutputs_11_50_port, B(49) => 
                           SumOutputs_11_49_port, B(48) => 
                           SumOutputs_11_48_port, B(47) => 
                           SumOutputs_11_47_port, B(46) => 
                           SumOutputs_11_46_port, B(45) => 
                           SumOutputs_11_45_port, B(44) => 
                           SumOutputs_11_44_port, B(43) => 
                           SumOutputs_11_43_port, B(42) => 
                           SumOutputs_11_42_port, B(41) => 
                           SumOutputs_11_41_port, B(40) => 
                           SumOutputs_11_40_port, B(39) => 
                           SumOutputs_11_39_port, B(38) => 
                           SumOutputs_11_38_port, B(37) => 
                           SumOutputs_11_37_port, B(36) => 
                           SumOutputs_11_36_port, B(35) => 
                           SumOutputs_11_35_port, B(34) => 
                           SumOutputs_11_34_port, B(33) => 
                           SumOutputs_11_33_port, B(32) => 
                           SumOutputs_11_32_port, B(31) => 
                           SumOutputs_11_31_port, B(30) => 
                           SumOutputs_11_30_port, B(29) => 
                           SumOutputs_11_29_port, B(28) => 
                           SumOutputs_11_28_port, B(27) => 
                           SumOutputs_11_27_port, B(26) => 
                           SumOutputs_11_26_port, B(25) => 
                           SumOutputs_11_25_port, B(24) => 
                           SumOutputs_11_24_port, B(23) => 
                           SumOutputs_11_23_port, B(22) => 
                           SumOutputs_11_22_port, B(21) => 
                           SumOutputs_11_21_port, B(20) => 
                           SumOutputs_11_20_port, B(19) => 
                           SumOutputs_11_19_port, B(18) => 
                           SumOutputs_11_18_port, B(17) => 
                           SumOutputs_11_17_port, B(16) => 
                           SumOutputs_11_16_port, B(15) => 
                           SumOutputs_11_15_port, B(14) => 
                           SumOutputs_11_14_port, B(13) => 
                           SumOutputs_11_13_port, B(12) => 
                           SumOutputs_11_12_port, B(11) => 
                           SumOutputs_11_11_port, B(10) => 
                           SumOutputs_11_10_port, B(9) => SumOutputs_11_9_port,
                           B(8) => SumOutputs_11_8_port, B(7) => 
                           SumOutputs_11_7_port, B(6) => SumOutputs_11_6_port, 
                           B(5) => SumOutputs_11_5_port, B(4) => 
                           SumOutputs_11_4_port, B(3) => SumOutputs_11_3_port, 
                           B(2) => SumOutputs_11_2_port, B(1) => 
                           SumOutputs_11_1_port, B(0) => SumOutputs_11_0_port, 
                           Ci => X_Logic0_port, S(63) => SumOutputs_12_63_port,
                           S(62) => SumOutputs_12_62_port, S(61) => 
                           SumOutputs_12_61_port, S(60) => 
                           SumOutputs_12_60_port, S(59) => 
                           SumOutputs_12_59_port, S(58) => 
                           SumOutputs_12_58_port, S(57) => 
                           SumOutputs_12_57_port, S(56) => 
                           SumOutputs_12_56_port, S(55) => 
                           SumOutputs_12_55_port, S(54) => 
                           SumOutputs_12_54_port, S(53) => 
                           SumOutputs_12_53_port, S(52) => 
                           SumOutputs_12_52_port, S(51) => 
                           SumOutputs_12_51_port, S(50) => 
                           SumOutputs_12_50_port, S(49) => 
                           SumOutputs_12_49_port, S(48) => 
                           SumOutputs_12_48_port, S(47) => 
                           SumOutputs_12_47_port, S(46) => 
                           SumOutputs_12_46_port, S(45) => 
                           SumOutputs_12_45_port, S(44) => 
                           SumOutputs_12_44_port, S(43) => 
                           SumOutputs_12_43_port, S(42) => 
                           SumOutputs_12_42_port, S(41) => 
                           SumOutputs_12_41_port, S(40) => 
                           SumOutputs_12_40_port, S(39) => 
                           SumOutputs_12_39_port, S(38) => 
                           SumOutputs_12_38_port, S(37) => 
                           SumOutputs_12_37_port, S(36) => 
                           SumOutputs_12_36_port, S(35) => 
                           SumOutputs_12_35_port, S(34) => 
                           SumOutputs_12_34_port, S(33) => 
                           SumOutputs_12_33_port, S(32) => 
                           SumOutputs_12_32_port, S(31) => 
                           SumOutputs_12_31_port, S(30) => 
                           SumOutputs_12_30_port, S(29) => 
                           SumOutputs_12_29_port, S(28) => 
                           SumOutputs_12_28_port, S(27) => 
                           SumOutputs_12_27_port, S(26) => 
                           SumOutputs_12_26_port, S(25) => 
                           SumOutputs_12_25_port, S(24) => 
                           SumOutputs_12_24_port, S(23) => 
                           SumOutputs_12_23_port, S(22) => 
                           SumOutputs_12_22_port, S(21) => 
                           SumOutputs_12_21_port, S(20) => 
                           SumOutputs_12_20_port, S(19) => 
                           SumOutputs_12_19_port, S(18) => 
                           SumOutputs_12_18_port, S(17) => 
                           SumOutputs_12_17_port, S(16) => 
                           SumOutputs_12_16_port, S(15) => 
                           SumOutputs_12_15_port, S(14) => 
                           SumOutputs_12_14_port, S(13) => 
                           SumOutputs_12_13_port, S(12) => 
                           SumOutputs_12_12_port, S(11) => 
                           SumOutputs_12_11_port, S(10) => 
                           SumOutputs_12_10_port, S(9) => SumOutputs_12_9_port,
                           S(8) => SumOutputs_12_8_port, S(7) => 
                           SumOutputs_12_7_port, S(6) => SumOutputs_12_6_port, 
                           S(5) => SumOutputs_12_5_port, S(4) => 
                           SumOutputs_12_4_port, S(3) => SumOutputs_12_3_port, 
                           S(2) => SumOutputs_12_2_port, S(1) => 
                           SumOutputs_12_1_port, S(0) => SumOutputs_12_0_port, 
                           Co => n_1139);
   SUMI_13 : RCA_NbitRca64_18 port map( A(63) => MuxOutputs_14_63_port, A(62) 
                           => MuxOutputs_14_62_port, A(61) => 
                           MuxOutputs_14_61_port, A(60) => 
                           MuxOutputs_14_60_port, A(59) => 
                           MuxOutputs_14_59_port, A(58) => 
                           MuxOutputs_14_58_port, A(57) => 
                           MuxOutputs_14_57_port, A(56) => 
                           MuxOutputs_14_56_port, A(55) => 
                           MuxOutputs_14_55_port, A(54) => 
                           MuxOutputs_14_54_port, A(53) => 
                           MuxOutputs_14_53_port, A(52) => 
                           MuxOutputs_14_52_port, A(51) => 
                           MuxOutputs_14_51_port, A(50) => 
                           MuxOutputs_14_50_port, A(49) => 
                           MuxOutputs_14_49_port, A(48) => 
                           MuxOutputs_14_48_port, A(47) => 
                           MuxOutputs_14_47_port, A(46) => 
                           MuxOutputs_14_46_port, A(45) => 
                           MuxOutputs_14_45_port, A(44) => 
                           MuxOutputs_14_44_port, A(43) => 
                           MuxOutputs_14_43_port, A(42) => 
                           MuxOutputs_14_42_port, A(41) => 
                           MuxOutputs_14_41_port, A(40) => 
                           MuxOutputs_14_40_port, A(39) => 
                           MuxOutputs_14_39_port, A(38) => 
                           MuxOutputs_14_38_port, A(37) => 
                           MuxOutputs_14_37_port, A(36) => 
                           MuxOutputs_14_36_port, A(35) => 
                           MuxOutputs_14_35_port, A(34) => 
                           MuxOutputs_14_34_port, A(33) => 
                           MuxOutputs_14_33_port, A(32) => 
                           MuxOutputs_14_32_port, A(31) => 
                           MuxOutputs_14_31_port, A(30) => 
                           MuxOutputs_14_30_port, A(29) => 
                           MuxOutputs_14_29_port, A(28) => 
                           MuxOutputs_14_28_port, A(27) => 
                           MuxOutputs_14_27_port, A(26) => 
                           MuxOutputs_14_26_port, A(25) => 
                           MuxOutputs_14_25_port, A(24) => 
                           MuxOutputs_14_24_port, A(23) => 
                           MuxOutputs_14_23_port, A(22) => 
                           MuxOutputs_14_22_port, A(21) => 
                           MuxOutputs_14_21_port, A(20) => 
                           MuxOutputs_14_20_port, A(19) => 
                           MuxOutputs_14_19_port, A(18) => 
                           MuxOutputs_14_18_port, A(17) => 
                           MuxOutputs_14_17_port, A(16) => 
                           MuxOutputs_14_16_port, A(15) => 
                           MuxOutputs_14_15_port, A(14) => 
                           MuxOutputs_14_14_port, A(13) => 
                           MuxOutputs_14_13_port, A(12) => 
                           MuxOutputs_14_12_port, A(11) => 
                           MuxOutputs_14_11_port, A(10) => 
                           MuxOutputs_14_10_port, A(9) => MuxOutputs_14_9_port,
                           A(8) => MuxOutputs_14_8_port, A(7) => 
                           MuxOutputs_14_7_port, A(6) => MuxOutputs_14_6_port, 
                           A(5) => MuxOutputs_14_5_port, A(4) => 
                           MuxOutputs_14_4_port, A(3) => MuxOutputs_14_3_port, 
                           A(2) => MuxOutputs_14_2_port, A(1) => 
                           MuxOutputs_14_1_port, A(0) => MuxOutputs_14_0_port, 
                           B(63) => SumOutputs_12_63_port, B(62) => 
                           SumOutputs_12_62_port, B(61) => 
                           SumOutputs_12_61_port, B(60) => 
                           SumOutputs_12_60_port, B(59) => 
                           SumOutputs_12_59_port, B(58) => 
                           SumOutputs_12_58_port, B(57) => 
                           SumOutputs_12_57_port, B(56) => 
                           SumOutputs_12_56_port, B(55) => 
                           SumOutputs_12_55_port, B(54) => 
                           SumOutputs_12_54_port, B(53) => 
                           SumOutputs_12_53_port, B(52) => 
                           SumOutputs_12_52_port, B(51) => 
                           SumOutputs_12_51_port, B(50) => 
                           SumOutputs_12_50_port, B(49) => 
                           SumOutputs_12_49_port, B(48) => 
                           SumOutputs_12_48_port, B(47) => 
                           SumOutputs_12_47_port, B(46) => 
                           SumOutputs_12_46_port, B(45) => 
                           SumOutputs_12_45_port, B(44) => 
                           SumOutputs_12_44_port, B(43) => 
                           SumOutputs_12_43_port, B(42) => 
                           SumOutputs_12_42_port, B(41) => 
                           SumOutputs_12_41_port, B(40) => 
                           SumOutputs_12_40_port, B(39) => 
                           SumOutputs_12_39_port, B(38) => 
                           SumOutputs_12_38_port, B(37) => 
                           SumOutputs_12_37_port, B(36) => 
                           SumOutputs_12_36_port, B(35) => 
                           SumOutputs_12_35_port, B(34) => 
                           SumOutputs_12_34_port, B(33) => 
                           SumOutputs_12_33_port, B(32) => 
                           SumOutputs_12_32_port, B(31) => 
                           SumOutputs_12_31_port, B(30) => 
                           SumOutputs_12_30_port, B(29) => 
                           SumOutputs_12_29_port, B(28) => 
                           SumOutputs_12_28_port, B(27) => 
                           SumOutputs_12_27_port, B(26) => 
                           SumOutputs_12_26_port, B(25) => 
                           SumOutputs_12_25_port, B(24) => 
                           SumOutputs_12_24_port, B(23) => 
                           SumOutputs_12_23_port, B(22) => 
                           SumOutputs_12_22_port, B(21) => 
                           SumOutputs_12_21_port, B(20) => 
                           SumOutputs_12_20_port, B(19) => 
                           SumOutputs_12_19_port, B(18) => 
                           SumOutputs_12_18_port, B(17) => 
                           SumOutputs_12_17_port, B(16) => 
                           SumOutputs_12_16_port, B(15) => 
                           SumOutputs_12_15_port, B(14) => 
                           SumOutputs_12_14_port, B(13) => 
                           SumOutputs_12_13_port, B(12) => 
                           SumOutputs_12_12_port, B(11) => 
                           SumOutputs_12_11_port, B(10) => 
                           SumOutputs_12_10_port, B(9) => SumOutputs_12_9_port,
                           B(8) => SumOutputs_12_8_port, B(7) => 
                           SumOutputs_12_7_port, B(6) => SumOutputs_12_6_port, 
                           B(5) => SumOutputs_12_5_port, B(4) => 
                           SumOutputs_12_4_port, B(3) => SumOutputs_12_3_port, 
                           B(2) => SumOutputs_12_2_port, B(1) => 
                           SumOutputs_12_1_port, B(0) => SumOutputs_12_0_port, 
                           Ci => X_Logic0_port, S(63) => SumOutputs_13_63_port,
                           S(62) => SumOutputs_13_62_port, S(61) => 
                           SumOutputs_13_61_port, S(60) => 
                           SumOutputs_13_60_port, S(59) => 
                           SumOutputs_13_59_port, S(58) => 
                           SumOutputs_13_58_port, S(57) => 
                           SumOutputs_13_57_port, S(56) => 
                           SumOutputs_13_56_port, S(55) => 
                           SumOutputs_13_55_port, S(54) => 
                           SumOutputs_13_54_port, S(53) => 
                           SumOutputs_13_53_port, S(52) => 
                           SumOutputs_13_52_port, S(51) => 
                           SumOutputs_13_51_port, S(50) => 
                           SumOutputs_13_50_port, S(49) => 
                           SumOutputs_13_49_port, S(48) => 
                           SumOutputs_13_48_port, S(47) => 
                           SumOutputs_13_47_port, S(46) => 
                           SumOutputs_13_46_port, S(45) => 
                           SumOutputs_13_45_port, S(44) => 
                           SumOutputs_13_44_port, S(43) => 
                           SumOutputs_13_43_port, S(42) => 
                           SumOutputs_13_42_port, S(41) => 
                           SumOutputs_13_41_port, S(40) => 
                           SumOutputs_13_40_port, S(39) => 
                           SumOutputs_13_39_port, S(38) => 
                           SumOutputs_13_38_port, S(37) => 
                           SumOutputs_13_37_port, S(36) => 
                           SumOutputs_13_36_port, S(35) => 
                           SumOutputs_13_35_port, S(34) => 
                           SumOutputs_13_34_port, S(33) => 
                           SumOutputs_13_33_port, S(32) => 
                           SumOutputs_13_32_port, S(31) => 
                           SumOutputs_13_31_port, S(30) => 
                           SumOutputs_13_30_port, S(29) => 
                           SumOutputs_13_29_port, S(28) => 
                           SumOutputs_13_28_port, S(27) => 
                           SumOutputs_13_27_port, S(26) => 
                           SumOutputs_13_26_port, S(25) => 
                           SumOutputs_13_25_port, S(24) => 
                           SumOutputs_13_24_port, S(23) => 
                           SumOutputs_13_23_port, S(22) => 
                           SumOutputs_13_22_port, S(21) => 
                           SumOutputs_13_21_port, S(20) => 
                           SumOutputs_13_20_port, S(19) => 
                           SumOutputs_13_19_port, S(18) => 
                           SumOutputs_13_18_port, S(17) => 
                           SumOutputs_13_17_port, S(16) => 
                           SumOutputs_13_16_port, S(15) => 
                           SumOutputs_13_15_port, S(14) => 
                           SumOutputs_13_14_port, S(13) => 
                           SumOutputs_13_13_port, S(12) => 
                           SumOutputs_13_12_port, S(11) => 
                           SumOutputs_13_11_port, S(10) => 
                           SumOutputs_13_10_port, S(9) => SumOutputs_13_9_port,
                           S(8) => SumOutputs_13_8_port, S(7) => 
                           SumOutputs_13_7_port, S(6) => SumOutputs_13_6_port, 
                           S(5) => SumOutputs_13_5_port, S(4) => 
                           SumOutputs_13_4_port, S(3) => SumOutputs_13_3_port, 
                           S(2) => SumOutputs_13_2_port, S(1) => 
                           SumOutputs_13_1_port, S(0) => SumOutputs_13_0_port, 
                           Co => n_1140);
   SUMI_14 : RCA_NbitRca64_17 port map( A(63) => MuxOutputs_15_63_port, A(62) 
                           => MuxOutputs_15_62_port, A(61) => 
                           MuxOutputs_15_61_port, A(60) => 
                           MuxOutputs_15_60_port, A(59) => 
                           MuxOutputs_15_59_port, A(58) => 
                           MuxOutputs_15_58_port, A(57) => 
                           MuxOutputs_15_57_port, A(56) => 
                           MuxOutputs_15_56_port, A(55) => 
                           MuxOutputs_15_55_port, A(54) => 
                           MuxOutputs_15_54_port, A(53) => 
                           MuxOutputs_15_53_port, A(52) => 
                           MuxOutputs_15_52_port, A(51) => 
                           MuxOutputs_15_51_port, A(50) => 
                           MuxOutputs_15_50_port, A(49) => 
                           MuxOutputs_15_49_port, A(48) => 
                           MuxOutputs_15_48_port, A(47) => 
                           MuxOutputs_15_47_port, A(46) => 
                           MuxOutputs_15_46_port, A(45) => 
                           MuxOutputs_15_45_port, A(44) => 
                           MuxOutputs_15_44_port, A(43) => 
                           MuxOutputs_15_43_port, A(42) => 
                           MuxOutputs_15_42_port, A(41) => 
                           MuxOutputs_15_41_port, A(40) => 
                           MuxOutputs_15_40_port, A(39) => 
                           MuxOutputs_15_39_port, A(38) => 
                           MuxOutputs_15_38_port, A(37) => 
                           MuxOutputs_15_37_port, A(36) => 
                           MuxOutputs_15_36_port, A(35) => 
                           MuxOutputs_15_35_port, A(34) => 
                           MuxOutputs_15_34_port, A(33) => 
                           MuxOutputs_15_33_port, A(32) => 
                           MuxOutputs_15_32_port, A(31) => 
                           MuxOutputs_15_31_port, A(30) => 
                           MuxOutputs_15_30_port, A(29) => 
                           MuxOutputs_15_29_port, A(28) => 
                           MuxOutputs_15_28_port, A(27) => 
                           MuxOutputs_15_27_port, A(26) => 
                           MuxOutputs_15_26_port, A(25) => 
                           MuxOutputs_15_25_port, A(24) => 
                           MuxOutputs_15_24_port, A(23) => 
                           MuxOutputs_15_23_port, A(22) => 
                           MuxOutputs_15_22_port, A(21) => 
                           MuxOutputs_15_21_port, A(20) => 
                           MuxOutputs_15_20_port, A(19) => 
                           MuxOutputs_15_19_port, A(18) => 
                           MuxOutputs_15_18_port, A(17) => 
                           MuxOutputs_15_17_port, A(16) => 
                           MuxOutputs_15_16_port, A(15) => 
                           MuxOutputs_15_15_port, A(14) => 
                           MuxOutputs_15_14_port, A(13) => 
                           MuxOutputs_15_13_port, A(12) => 
                           MuxOutputs_15_12_port, A(11) => 
                           MuxOutputs_15_11_port, A(10) => 
                           MuxOutputs_15_10_port, A(9) => MuxOutputs_15_9_port,
                           A(8) => MuxOutputs_15_8_port, A(7) => 
                           MuxOutputs_15_7_port, A(6) => MuxOutputs_15_6_port, 
                           A(5) => MuxOutputs_15_5_port, A(4) => 
                           MuxOutputs_15_4_port, A(3) => MuxOutputs_15_3_port, 
                           A(2) => MuxOutputs_15_2_port, A(1) => 
                           MuxOutputs_15_1_port, A(0) => MuxOutputs_15_0_port, 
                           B(63) => SumOutputs_13_63_port, B(62) => 
                           SumOutputs_13_62_port, B(61) => 
                           SumOutputs_13_61_port, B(60) => 
                           SumOutputs_13_60_port, B(59) => 
                           SumOutputs_13_59_port, B(58) => 
                           SumOutputs_13_58_port, B(57) => 
                           SumOutputs_13_57_port, B(56) => 
                           SumOutputs_13_56_port, B(55) => 
                           SumOutputs_13_55_port, B(54) => 
                           SumOutputs_13_54_port, B(53) => 
                           SumOutputs_13_53_port, B(52) => 
                           SumOutputs_13_52_port, B(51) => 
                           SumOutputs_13_51_port, B(50) => 
                           SumOutputs_13_50_port, B(49) => 
                           SumOutputs_13_49_port, B(48) => 
                           SumOutputs_13_48_port, B(47) => 
                           SumOutputs_13_47_port, B(46) => 
                           SumOutputs_13_46_port, B(45) => 
                           SumOutputs_13_45_port, B(44) => 
                           SumOutputs_13_44_port, B(43) => 
                           SumOutputs_13_43_port, B(42) => 
                           SumOutputs_13_42_port, B(41) => 
                           SumOutputs_13_41_port, B(40) => 
                           SumOutputs_13_40_port, B(39) => 
                           SumOutputs_13_39_port, B(38) => 
                           SumOutputs_13_38_port, B(37) => 
                           SumOutputs_13_37_port, B(36) => 
                           SumOutputs_13_36_port, B(35) => 
                           SumOutputs_13_35_port, B(34) => 
                           SumOutputs_13_34_port, B(33) => 
                           SumOutputs_13_33_port, B(32) => 
                           SumOutputs_13_32_port, B(31) => 
                           SumOutputs_13_31_port, B(30) => 
                           SumOutputs_13_30_port, B(29) => 
                           SumOutputs_13_29_port, B(28) => 
                           SumOutputs_13_28_port, B(27) => 
                           SumOutputs_13_27_port, B(26) => 
                           SumOutputs_13_26_port, B(25) => 
                           SumOutputs_13_25_port, B(24) => 
                           SumOutputs_13_24_port, B(23) => 
                           SumOutputs_13_23_port, B(22) => 
                           SumOutputs_13_22_port, B(21) => 
                           SumOutputs_13_21_port, B(20) => 
                           SumOutputs_13_20_port, B(19) => 
                           SumOutputs_13_19_port, B(18) => 
                           SumOutputs_13_18_port, B(17) => 
                           SumOutputs_13_17_port, B(16) => 
                           SumOutputs_13_16_port, B(15) => 
                           SumOutputs_13_15_port, B(14) => 
                           SumOutputs_13_14_port, B(13) => 
                           SumOutputs_13_13_port, B(12) => 
                           SumOutputs_13_12_port, B(11) => 
                           SumOutputs_13_11_port, B(10) => 
                           SumOutputs_13_10_port, B(9) => SumOutputs_13_9_port,
                           B(8) => SumOutputs_13_8_port, B(7) => 
                           SumOutputs_13_7_port, B(6) => SumOutputs_13_6_port, 
                           B(5) => SumOutputs_13_5_port, B(4) => 
                           SumOutputs_13_4_port, B(3) => SumOutputs_13_3_port, 
                           B(2) => SumOutputs_13_2_port, B(1) => 
                           SumOutputs_13_1_port, B(0) => SumOutputs_13_0_port, 
                           Ci => X_Logic0_port, S(63) => P(63), S(62) => P(62),
                           S(61) => P(61), S(60) => P(60), S(59) => P(59), 
                           S(58) => P(58), S(57) => P(57), S(56) => P(56), 
                           S(55) => P(55), S(54) => P(54), S(53) => P(53), 
                           S(52) => P(52), S(51) => P(51), S(50) => P(50), 
                           S(49) => P(49), S(48) => P(48), S(47) => P(47), 
                           S(46) => P(46), S(45) => P(45), S(44) => P(44), 
                           S(43) => P(43), S(42) => P(42), S(41) => P(41), 
                           S(40) => P(40), S(39) => P(39), S(38) => P(38), 
                           S(37) => P(37), S(36) => P(36), S(35) => P(35), 
                           S(34) => P(34), S(33) => P(33), S(32) => P(32), 
                           S(31) => P(31), S(30) => P(30), S(29) => P(29), 
                           S(28) => P(28), S(27) => P(27), S(26) => P(26), 
                           S(25) => P(25), S(24) => P(24), S(23) => P(23), 
                           S(22) => P(22), S(21) => P(21), S(20) => P(20), 
                           S(19) => P(19), S(18) => P(18), S(17) => P(17), 
                           S(16) => P(16), S(15) => P(15), S(14) => P(14), 
                           S(13) => P(13), S(12) => P(12), S(11) => P(11), 
                           S(10) => P(10), S(9) => P(9), S(8) => P(8), S(7) => 
                           P(7), S(6) => P(6), S(5) => P(5), S(4) => P(4), S(3)
                           => P(3), S(2) => P(2), S(1) => P(1), S(0) => P(0), 
                           Co => n_1141);
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   n8 <= '0';
   U3 : BUF_X1 port map( A => negative_inputs_0_4_port, Z => n12);
   U4 : BUF_X1 port map( A => negative_inputs_0_14_port, Z => n9);
   U5 : BUF_X1 port map( A => negative_inputs_0_17_port, Z => n10);
   U6 : CLKBUF_X1 port map( A => negative_inputs_0_3_port, Z => n14);
   U7 : BUF_X1 port map( A => negative_inputs_0_5_port, Z => n11);
   U8 : CLKBUF_X1 port map( A => negative_inputs_1_3_port, Z => n13);
   U9 : CLKBUF_X1 port map( A => negative_inputs_5_11_port, Z => n54);
   U11 : CLKBUF_X1 port map( A => negative_inputs_5_7_port, Z => n46);
   U12 : BUF_X1 port map( A => A(1), Z => n15);
   U13 : CLKBUF_X1 port map( A => negative_inputs_5_10_port, Z => n52);
   U14 : CLKBUF_X1 port map( A => negative_inputs_5_12_port, Z => n56);
   U15 : CLKBUF_X1 port map( A => negative_inputs_5_14_port, Z => n60);
   U16 : CLKBUF_X1 port map( A => negative_inputs_5_19_port, Z => n70);
   U17 : CLKBUF_X1 port map( A => negative_inputs_5_13_port, Z => n58);
   U18 : CLKBUF_X1 port map( A => negative_inputs_5_15_port, Z => n62);
   U19 : BUF_X1 port map( A => negative_inputs_5_8_port, Z => n48);
   U20 : BUF_X1 port map( A => A(0), Z => n18);
   U21 : INV_X1 port map( A => negative_inputs_1_42_port, ZN => n16);
   U22 : INV_X1 port map( A => n16, ZN => n17);
   U23 : CLKBUF_X1 port map( A => negative_inputs_5_9_port, Z => n50);
   U24 : CLKBUF_X1 port map( A => negative_inputs_11_47_port, Z => n115);
   U25 : CLKBUF_X1 port map( A => negative_inputs_12_47_port, Z => n113);
   U26 : CLKBUF_X1 port map( A => negative_inputs_13_47_port, Z => n111);
   U27 : CLKBUF_X1 port map( A => negative_inputs_15_16_port, Z => n45);
   U28 : CLKBUF_X1 port map( A => negative_inputs_15_17_port, Z => n47);
   U29 : CLKBUF_X1 port map( A => negative_inputs_15_19_port, Z => n51);
   U30 : CLKBUF_X1 port map( A => negative_inputs_15_20_port, Z => n53);
   U31 : CLKBUF_X1 port map( A => negative_inputs_15_21_port, Z => n55);
   U32 : CLKBUF_X1 port map( A => negative_inputs_15_22_port, Z => n57);
   U33 : CLKBUF_X1 port map( A => negative_inputs_15_23_port, Z => n59);
   U34 : CLKBUF_X1 port map( A => negative_inputs_15_24_port, Z => n61);
   U35 : CLKBUF_X1 port map( A => negative_inputs_15_27_port, Z => n67);
   U36 : CLKBUF_X1 port map( A => negative_inputs_15_26_port, Z => n65);
   U37 : CLKBUF_X1 port map( A => negative_inputs_15_25_port, Z => n63);
   U38 : CLKBUF_X1 port map( A => negative_inputs_15_29_port, Z => n71);
   U39 : CLKBUF_X1 port map( A => negative_inputs_15_28_port, Z => n69);
   U40 : CLKBUF_X1 port map( A => negative_inputs_15_31_port, Z => n75);
   U41 : CLKBUF_X1 port map( A => negative_inputs_15_30_port, Z => n73);
   U42 : CLKBUF_X1 port map( A => negative_inputs_15_32_port, Z => n77);
   U43 : CLKBUF_X1 port map( A => negative_inputs_15_33_port, Z => n79);
   U44 : CLKBUF_X1 port map( A => negative_inputs_15_34_port, Z => n81);
   U45 : CLKBUF_X1 port map( A => negative_inputs_15_35_port, Z => n83);
   U46 : CLKBUF_X1 port map( A => negative_inputs_15_36_port, Z => n85);
   U47 : CLKBUF_X1 port map( A => negative_inputs_14_47_port, Z => n109);
   U48 : CLKBUF_X1 port map( A => negative_inputs_15_37_port, Z => n87);
   U49 : CLKBUF_X1 port map( A => negative_inputs_15_38_port, Z => n89);
   U50 : CLKBUF_X1 port map( A => negative_inputs_15_39_port, Z => n91);
   U51 : CLKBUF_X1 port map( A => negative_inputs_15_40_port, Z => n93);
   U52 : CLKBUF_X1 port map( A => negative_inputs_15_41_port, Z => n95);
   U53 : CLKBUF_X1 port map( A => negative_inputs_15_42_port, Z => n97);
   U54 : CLKBUF_X1 port map( A => negative_inputs_15_43_port, Z => n99);
   U55 : CLKBUF_X1 port map( A => negative_inputs_15_44_port, Z => n101);
   U56 : CLKBUF_X1 port map( A => negative_inputs_15_45_port, Z => n103);
   U57 : CLKBUF_X1 port map( A => negative_inputs_15_46_port, Z => n105);
   U58 : CLKBUF_X1 port map( A => negative_inputs_15_47_port, Z => n107);
   U59 : CLKBUF_X1 port map( A => negative_inputs_15_15_port, Z => n43);
   U60 : CLKBUF_X1 port map( A => positive_inputs_15_15_port, Z => n121);
   U61 : CLKBUF_X1 port map( A => negative_inputs_15_18_port, Z => n49);
   U62 : CLKBUF_X1 port map( A => negative_inputs_10_47_port, Z => n116);
   U63 : BUF_X2 port map( A => negative_inputs_0_49_port, Z => n41);
   U64 : BUF_X2 port map( A => negative_inputs_0_51_port, Z => n39);
   U65 : BUF_X2 port map( A => negative_inputs_0_52_port, Z => n40);
   U66 : BUF_X1 port map( A => positive_inputs_5_19_port, Z => n148);
   U67 : BUF_X1 port map( A => positive_inputs_5_20_port, Z => n150);
   U68 : BUF_X1 port map( A => positive_inputs_5_21_port, Z => n152);
   U69 : BUF_X1 port map( A => positive_inputs_5_22_port, Z => n154);
   U70 : BUF_X1 port map( A => positive_inputs_5_23_port, Z => n156);
   U71 : BUF_X1 port map( A => positive_inputs_5_24_port, Z => n158);
   U72 : BUF_X1 port map( A => positive_inputs_5_25_port, Z => n160);
   U73 : BUF_X1 port map( A => positive_inputs_5_26_port, Z => n162);
   U74 : BUF_X1 port map( A => positive_inputs_5_27_port, Z => n164);
   U75 : BUF_X1 port map( A => positive_inputs_5_28_port, Z => n166);
   U76 : BUF_X1 port map( A => positive_inputs_5_29_port, Z => n168);
   U77 : BUF_X1 port map( A => positive_inputs_5_30_port, Z => n170);
   U78 : BUF_X1 port map( A => positive_inputs_5_31_port, Z => n172);
   U79 : BUF_X1 port map( A => positive_inputs_5_32_port, Z => n174);
   U80 : BUF_X1 port map( A => positive_inputs_5_33_port, Z => n176);
   U81 : BUF_X1 port map( A => positive_inputs_5_34_port, Z => n178);
   U82 : BUF_X1 port map( A => positive_inputs_3_37_port, Z => n22);
   U83 : BUF_X1 port map( A => positive_inputs_2_37_port, Z => n23);
   U84 : BUF_X1 port map( A => positive_inputs_1_37_port, Z => n24);
   U85 : BUF_X1 port map( A => positive_inputs_5_35_port, Z => n180);
   U86 : BUF_X1 port map( A => positive_inputs_5_36_port, Z => n19);
   U87 : BUF_X1 port map( A => positive_inputs_5_37_port, Z => n20);
   U88 : BUF_X1 port map( A => positive_inputs_4_37_port, Z => n21);
   U89 : BUF_X1 port map( A => positive_inputs_2_47_port, Z => n38);
   U90 : BUF_X1 port map( A => positive_inputs_4_47_port, Z => n37);
   U91 : BUF_X1 port map( A => positive_inputs_5_47_port, Z => n36);
   U92 : BUF_X1 port map( A => positive_inputs_6_47_port, Z => n35);
   U93 : BUF_X1 port map( A => positive_inputs_7_47_port, Z => n34);
   U94 : BUF_X1 port map( A => positive_inputs_8_47_port, Z => n33);
   U95 : BUF_X1 port map( A => positive_inputs_9_47_port, Z => n32);
   U96 : BUF_X1 port map( A => positive_inputs_10_47_port, Z => n31);
   U97 : BUF_X1 port map( A => negative_inputs_1_37_port, Z => n114);
   U98 : BUF_X1 port map( A => negative_inputs_2_37_port, Z => n112);
   U99 : BUF_X1 port map( A => negative_inputs_3_37_port, Z => n110);
   U100 : BUF_X1 port map( A => negative_inputs_5_6_port, Z => n44);
   U101 : BUF_X1 port map( A => negative_inputs_5_16_port, Z => n64);
   U102 : BUF_X1 port map( A => negative_inputs_5_17_port, Z => n66);
   U103 : BUF_X1 port map( A => negative_inputs_5_18_port, Z => n68);
   U104 : BUF_X1 port map( A => negative_inputs_5_20_port, Z => n72);
   U105 : BUF_X1 port map( A => negative_inputs_5_21_port, Z => n74);
   U106 : BUF_X1 port map( A => negative_inputs_5_22_port, Z => n76);
   U107 : BUF_X1 port map( A => negative_inputs_5_24_port, Z => n80);
   U108 : CLKBUF_X1 port map( A => negative_inputs_4_37_port, Z => n108);
   U109 : BUF_X1 port map( A => negative_inputs_5_25_port, Z => n82);
   U110 : BUF_X1 port map( A => negative_inputs_5_26_port, Z => n84);
   U111 : BUF_X1 port map( A => negative_inputs_5_27_port, Z => n86);
   U112 : BUF_X1 port map( A => negative_inputs_5_28_port, Z => n88);
   U113 : BUF_X1 port map( A => negative_inputs_5_30_port, Z => n92);
   U114 : BUF_X1 port map( A => negative_inputs_5_31_port, Z => n94);
   U115 : BUF_X1 port map( A => negative_inputs_5_32_port, Z => n96);
   U116 : BUF_X1 port map( A => negative_inputs_5_33_port, Z => n98);
   U117 : BUF_X1 port map( A => negative_inputs_5_34_port, Z => n100);
   U118 : BUF_X1 port map( A => negative_inputs_5_35_port, Z => n102);
   U119 : BUF_X1 port map( A => negative_inputs_5_36_port, Z => n104);
   U120 : BUF_X1 port map( A => negative_inputs_5_37_port, Z => n106);
   U121 : BUF_X1 port map( A => negative_inputs_5_23_port, Z => n78);
   U122 : BUF_X1 port map( A => negative_inputs_5_29_port, Z => n90);
   U123 : BUF_X1 port map( A => negative_inputs_7_47_port, Z => n119);
   U124 : BUF_X1 port map( A => negative_inputs_8_47_port, Z => n118);
   U125 : BUF_X1 port map( A => negative_inputs_9_47_port, Z => n117);
   U126 : BUF_X1 port map( A => negative_inputs_5_5_port, Z => n42);
   U127 : BUF_X1 port map( A => positive_inputs_15_16_port, Z => n123);
   U128 : BUF_X1 port map( A => positive_inputs_15_18_port, Z => n127);
   U129 : BUF_X1 port map( A => positive_inputs_15_19_port, Z => n129);
   U130 : BUF_X1 port map( A => positive_inputs_15_17_port, Z => n125);
   U131 : BUF_X1 port map( A => positive_inputs_15_20_port, Z => n131);
   U132 : BUF_X1 port map( A => positive_inputs_15_21_port, Z => n133);
   U133 : BUF_X1 port map( A => positive_inputs_15_22_port, Z => n135);
   U134 : BUF_X1 port map( A => positive_inputs_15_23_port, Z => n137);
   U135 : BUF_X1 port map( A => positive_inputs_15_24_port, Z => n139);
   U136 : BUF_X1 port map( A => positive_inputs_15_25_port, Z => n141);
   U137 : BUF_X1 port map( A => positive_inputs_15_26_port, Z => n143);
   U138 : BUF_X1 port map( A => positive_inputs_15_27_port, Z => n145);
   U139 : BUF_X1 port map( A => positive_inputs_15_28_port, Z => n147);
   U140 : BUF_X1 port map( A => positive_inputs_15_29_port, Z => n149);
   U141 : BUF_X1 port map( A => positive_inputs_15_30_port, Z => n151);
   U142 : BUF_X1 port map( A => positive_inputs_15_31_port, Z => n153);
   U143 : BUF_X1 port map( A => positive_inputs_15_32_port, Z => n155);
   U144 : BUF_X1 port map( A => positive_inputs_15_33_port, Z => n157);
   U145 : BUF_X1 port map( A => positive_inputs_15_34_port, Z => n159);
   U146 : BUF_X1 port map( A => positive_inputs_15_35_port, Z => n161);
   U147 : BUF_X1 port map( A => positive_inputs_15_36_port, Z => n163);
   U148 : BUF_X1 port map( A => positive_inputs_15_37_port, Z => n165);
   U149 : BUF_X1 port map( A => positive_inputs_15_38_port, Z => n167);
   U150 : BUF_X1 port map( A => positive_inputs_15_39_port, Z => n169);
   U151 : BUF_X1 port map( A => positive_inputs_15_40_port, Z => n171);
   U152 : BUF_X1 port map( A => positive_inputs_11_47_port, Z => n30);
   U153 : BUF_X1 port map( A => positive_inputs_15_41_port, Z => n173);
   U154 : BUF_X1 port map( A => positive_inputs_15_42_port, Z => n175);
   U155 : BUF_X1 port map( A => positive_inputs_13_47_port, Z => n28);
   U156 : BUF_X1 port map( A => positive_inputs_12_47_port, Z => n29);
   U157 : BUF_X1 port map( A => positive_inputs_15_43_port, Z => n177);
   U158 : BUF_X1 port map( A => positive_inputs_15_46_port, Z => n25);
   U159 : BUF_X1 port map( A => positive_inputs_15_44_port, Z => n179);
   U160 : BUF_X1 port map( A => positive_inputs_15_47_port, Z => n26);
   U161 : BUF_X1 port map( A => positive_inputs_14_47_port, Z => n27);
   U162 : BUF_X1 port map( A => positive_inputs_15_45_port, Z => n181);
   U163 : BUF_X1 port map( A => positive_inputs_5_6_port, Z => n122);
   U164 : BUF_X1 port map( A => positive_inputs_5_5_port, Z => n120);
   U165 : BUF_X1 port map( A => positive_inputs_5_8_port, Z => n126);
   U166 : BUF_X1 port map( A => positive_inputs_5_9_port, Z => n128);
   U167 : BUF_X1 port map( A => positive_inputs_5_7_port, Z => n124);
   U168 : BUF_X1 port map( A => positive_inputs_5_10_port, Z => n130);
   U169 : BUF_X1 port map( A => positive_inputs_5_11_port, Z => n132);
   U170 : BUF_X1 port map( A => positive_inputs_5_12_port, Z => n134);
   U171 : BUF_X1 port map( A => positive_inputs_5_13_port, Z => n136);
   U172 : BUF_X1 port map( A => positive_inputs_5_14_port, Z => n138);
   U173 : BUF_X1 port map( A => positive_inputs_5_15_port, Z => n140);
   U174 : BUF_X1 port map( A => positive_inputs_5_16_port, Z => n142);
   U175 : BUF_X1 port map( A => positive_inputs_5_17_port, Z => n144);
   U176 : BUF_X1 port map( A => positive_inputs_5_18_port, Z => n146);

end SYN_STRUCTURAL;
