
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_register_file is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_register_file;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_register_file.all;

entity register_file is

   port( CLK, RESET, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
         ADD_RD2 : in std_logic_vector (4 downto 0);  DATAIN : in 
         std_logic_vector (31 downto 0);  OUT1, OUT2 : out std_logic_vector (31
         downto 0));

end register_file;

architecture SYN_Behavioral of register_file is

   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component TINV_X1
      port( I, EN : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
      n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, 
      n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, 
      n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, 
      n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, 
      n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, 
      n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, 
      n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, 
      n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, 
      n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, 
      n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, 
      n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, 
      n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, 
      n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, 
      n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, 
      n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, 
      n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, 
      n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, 
      n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, 
      n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, 
      n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, 
      n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, 
      n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, 
      n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, 
      n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, 
      n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, 
      n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, 
      n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, 
      n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, 
      n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, 
      n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, 
      n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, 
      n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, 
      n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, 
      n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, 
      n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, 
      n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, 
      n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, 
      n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, 
      n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, 
      n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, 
      n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, 
      n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, 
      n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, 
      n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, 
      n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, 
      n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, 
      n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, 
      n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, 
      n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, 
      n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, 
      n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, 
      n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, 
      n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, 
      n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, 
      n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, 
      n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, 
      n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, 
      n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, 
      n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, 
      n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, 
      n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, 
      n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, 
      n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, 
      n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, 
      n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, 
      n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, 
      n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, 
      n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, 
      n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, 
      n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, 
      n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, 
      n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, 
      n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, 
      n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, 
      n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, 
      n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, 
      n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, 
      n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, 
      n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, 
      n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, 
      n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, 
      n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, 
      n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, 
      n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, 
      n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, 
      n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, 
      n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, 
      n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, 
      n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, 
      n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, 
      n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, 
      n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, 
      n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, 
      n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, 
      n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, 
      n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, 
      n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, 
      n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, 
      n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, 
      n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, 
      n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, 
      n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, 
      n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, 
      n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, 
      n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, 
      n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, 
      n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, 
      n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, 
      n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, 
      n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, 
      n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, 
      n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, 
      n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, 
      n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, 
      n2633, n2634, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, 
      n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, 
      n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, 
      n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, 
      n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, 
      n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, 
      n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, 
      n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, 
      n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, 
      n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, 
      n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, 
      n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, 
      n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, 
      n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, 
      n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, 
      n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, 
      n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, 
      n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, 
      n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, 
      n4930, n4931, n4932, n4933, n7879, n7880, n7881, n7882, n7883, n7884, 
      n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, 
      n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, 
      n7905, n7906, n7907, n7908, n7909, n7910, n7975, n7976, n7977, n7978, 
      n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, 
      n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, 
      n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, 
      n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, 
      n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, 
      n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, 
      n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, 
      n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, 
      n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, 
      n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, 
      n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, 
      n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, 
      n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, 
      n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, 
      n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, 
      n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, 
      n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, 
      n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, 
      n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, 
      n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, 
      n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, 
      n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, 
      n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, 
      n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, 
      n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, 
      n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, 
      n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, 
      n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, 
      n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, 
      n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, 
      n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, 
      n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, 
      n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, 
      n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, 
      n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, 
      n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, 
      n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, 
      n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, 
      n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, 
      n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, 
      n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, 
      n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, 
      n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, 
      n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, 
      n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, 
      n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, 
      n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, 
      n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, 
      n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, 
      n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, 
      n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, 
      n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, 
      n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, 
      n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, 
      n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, 
      n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, 
      n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, 
      n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, 
      n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, 
      n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, 
      n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, 
      n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, 
      n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, 
      n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, 
      n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, 
      n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, 
      n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, 
      n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, 
      n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, 
      n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, 
      n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, 
      n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, 
      n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, 
      n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, 
      n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, 
      n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, 
      n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, 
      n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, 
      n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, 
      n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, 
      n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, 
      n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, 
      n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, 
      n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, 
      n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, 
      n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, 
      n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, 
      n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, 
      n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, 
      n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, 
      n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, 
      n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, 
      n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, 
      n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, 
      n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, 
      n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, 
      n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, 
      n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, 
      n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, 
      n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, 
      n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, 
      n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, 
      n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, 
      n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, 
      n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, 
      n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, 
      n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, 
      n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, 
      n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, 
      n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, 
      n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, 
      n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, 
      n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, 
      n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, 
      n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, 
      n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, 
      n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, 
      n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, 
      n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, 
      n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, 
      n9921, n9922, n9923, n9925, n9926, n9927, n9928, n9929, n9930, n9931, 
      n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, 
      n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, 
      n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, 
      n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, 
      n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, 
      n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, 
      n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, 
      n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010, 
      n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019, 
      n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028, 
      n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037, 
      n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046, 
      n10047, n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055, 
      n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064, 
      n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073, 
      n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082, 
      n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091, 
      n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099, n10100, 
      n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109, 
      n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118, 
      n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127, 
      n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136, 
      n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145, 
      n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154, 
      n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163, 
      n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171, n10172, 
      n10173, n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181, 
      n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189, n10190, 
      n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199, 
      n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208, 
      n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217, 
      n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226, 
      n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234, n10235, 
      n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243, n10244, 
      n10245, n10246, n10247, n10248, n10249, n10250, n10251, n10252, n10253, 
      n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10261, n10262, 
      n10263, n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271, 
      n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280, 
      n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289, 
      n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298, 
      n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307, 
      n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315, n10316, 
      n10317, n10318, n10319, n10320, n10321, n10322, n10323, n10324, n10325, 
      n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333, n10334, 
      n10335, n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343, 
      n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352, 
      n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361, 
      n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370, 
      n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379, 
      n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387, n10388, 
      n10389, n10390, n10391, n10392, n10393, n10394, n10395, n10396, n10397, 
      n10398, n10399, n10400, n10401, n10402, n10403, n10404, n10405, n10406, 
      n10407, n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415, 
      n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424, 
      n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433, 
      n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442, 
      n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450, n10451, 
      n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459, n10460, 
      n10461, n10462, n10463, n10464, n10465, n10466, n10467, n10468, n10469, 
      n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477, n10478, 
      n10479, n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487, 
      n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496, 
      n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505, 
      n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514, 
      n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522, n10523, 
      n10525, n10526, n10527, n10528, n10529, n10530, n10531, n10532, n10533, 
      n10534, n10535, n10536, n10537, n10538, n10539, n10540, n10541, n10542, 
      n10543, n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551, 
      n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560, 
      n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569, 
      n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577, n10578, 
      n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586, n10587, 
      n10588, n10589, n10590, n10591, n10592, n10593, n10594, n10595, n10596, 
      n10597, n10598, n10599, n10600, n10601, n10602, n10603, n10604, n10605, 
      n10606, n10607, n10608, n10609, n10610, n10611, n10612, n10613, n10614, 
      n10615, n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623, 
      n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632, 
      n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641, 
      n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649, n10650, 
      n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658, n10659, 
      n10660, n10661, n10662, n10663, n10664, n10665, n10666, n10667, n10668, 
      n10669, n10670, n10671, n10672, n10673, n10674, n10675, n10676, n10677, 
      n10678, n10679, n10680, n10681, n10682, n10683, n10684, n10685, n10686, 
      n10687, n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695, 
      n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704, 
      n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713, 
      n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721, n10722, 
      n10723, n10724, n10725, n10726, n10727, n10728, n10729, n10730, n10731, 
      n10732, n10733, n10734, n10735, n10736, n10737, n10738, n10739, n10740, 
      n10741, n10742, n10743, n10744, n10745, n10746, n10747, n10748, n10749, 
      n10750, n10751, n10752, n10753, n10754, n10755, n10756, n10757, n10758, 
      n10759, n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767, 
      n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776, 
      n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785, 
      n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793, n10794, 
      n10795, n10796, n10797, n10798, n10799, n10800, n10801, n10802, n10803, 
      n10804, n10805, n10806, n10807, n10808, n10809, n10810, n10811, n10812, 
      n10813, n10814, n10815, n10816, n10817, n10818, n10819, n10820, n10821, 
      n10822, n10823, n10824, n10825, n10826, n10827, n10828, n10829, n10830, 
      n10831, n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839, 
      n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848, 
      n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857, 
      n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865, n10866, 
      n10867, n10868, n10869, n10870, n10871, n10872, n10873, n10874, n10875, 
      n10876, n10877, n10878, n10879, n10880, n10881, n10882, n10883, n10884, 
      n10885, n10886, n10887, n10888, n10889, n10890, n10891, n10892, n10893, 
      n10894, n10895, n10896, n10897, n10898, n10899, n10900, n10901, n10902, 
      n10903, n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911, 
      n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920, 
      n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929, 
      n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937, n10938, 
      n10939, n10940, n10941, n10942, n10943, n10944, n10945, n10946, n10947, 
      n10948, n10949, n10950, n10951, n10952, n10953, n10954, n10955, n10956, 
      n10957, n10958, n10959, n10960, n10961, n10962, n10963, n10964, n10965, 
      n10966, n10967, n10968, n10969, n10970, n10971, n10972, n10973, n10974, 
      n10975, n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983, 
      n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992, 
      n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001, 
      n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009, n11010, 
      n11011, n11012, n11013, n11014, n11015, n11016, n11017, n11018, n11019, 
      n11020, n11021, n11022, n11023, n11024, n11025, n11026, n11027, n11028, 
      n11029, n11030, n11031, n11032, n11033, n11034, n11035, n11036, n11037, 
      n11038, n11039, n11040, n11041, n11042, n11043, n11044, n11045, n11046, 
      n11047, n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055, 
      n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064, 
      n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073, 
      n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081, n11082, 
      n11083, n11084, n11085, n11086, n11087, n11088, n11089, n11090, n11091, 
      n11092, n11093, n11094, n11095, n11096, n11097, n11098, n11099, n11100, 
      n11101, n11102, n11103, n11104, n11105, n11106, n11107, n11108, n11109, 
      n11110, n11111, n11112, n11113, n11114, n11115, n11116, n11117, n11118, 
      n11119, n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127, 
      n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136, 
      n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145, 
      n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153, n11154, 
      n11155, n11156, n11157, n11158, n11159, n11160, n11161, n11162, n11163, 
      n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11203, n11204, 
      n11205, n11206, n11207, n11208, n11209, n11210, n11211, n11212, n11213, 
      n11214, n11215, n11216, n11217, n11218, n11219, n11220, n11221, n11222, 
      n11223, n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231, 
      n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240, 
      n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249, 
      n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258, 
      n11259, n11260, n11261, n11262, n11263, n11264, n11265, n11266, n11267, 
      n11268, n11269, n11270, n11271, n11272, n11273, n11274, n11275, n11276, 
      n11277, n11278, n11279, n11280, n11281, n11282, n11283, n11284, n11285, 
      n11286, n11287, n11288, n11289, n11290, n11291, n11324, n11325, n11326, 
      n11327, n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335, 
      n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344, 
      n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353, 
      n11354, n11355, n11388, n11389, n11390, n11391, n11392, n11393, n11394, 
      n11395, n11396, n11397, n11398, n11399, n11400, n11401, n11402, n11403, 
      n11404, n11405, n11406, n11407, n11408, n11409, n11410, n11411, n11412, 
      n11413, n11414, n11415, n11416, n11417, n11418, n11419, n11484, n11485, 
      n11486, n11487, n11488, n11489, n11490, n11491, n11492, n11493, n11494, 
      n11495, n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503, 
      n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512, 
      n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521, 
      n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530, 
      n11531, n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539, 
      n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547, n11548, 
      n11549, n11550, n11551, n11552, n11553, n11554, n11555, n11556, n11557, 
      n11558, n11559, n11560, n11561, n11562, n11563, n11564, n11565, n11566, 
      n11567, n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575, 
      n11576, n11577, n11578, n11579, n11580, n11613, n11614, n11615, n11616, 
      n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625, 
      n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633, n11634, 
      n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642, n11643, 
      n11644, n11677, n11678, n11679, n11680, n11681, n11682, n11683, n11684, 
      n11685, n11686, n11687, n11688, n11689, n11690, n11691, n11692, n11693, 
      n11694, n11695, n11696, n11697, n11698, n11699, n11700, n11701, n11702, 
      n11703, n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711, 
      n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720, 
      n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729, 
      n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738, 
      n11739, n11740, n11741, n11742, n11743, n11744, n11745, n11746, n11747, 
      n11748, n11749, n11750, n11751, n11752, n11753, n11754, n11755, n11756, 
      n11757, n11758, n11759, n11760, n11761, n11762, n11763, n11764, n11765, 
      n11766, n11767, n11768, n11769, n11770, n11771, n11772, n11837, n11838, 
      n11839, n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847, 
      n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856, 
      n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865, 
      n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873, n11874, 
      n11875, n11876, n11877, n11878, n11879, n11880, n11881, n11882, n11883, 
      n11884, n11885, n11886, n11887, n11888, n11889, n11890, n11891, n11892, 
      n11893, n11894, n11895, n11896, n11897, n11898, n11899, n11900, n11901, 
      n11902, n11903, n11904, n11905, n11906, n11907, n11908, n11909, n11910, 
      n11911, n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919, 
      n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928, 
      n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937, 
      n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945, n11946, 
      n11947, n11948, n11949, n11950, n11951, n11952, n11953, n11954, n11955, 
      n11956, n11957, n11958, n11959, n11960, n11961, n11962, n11963, n11964, 
      n11965, n11966, n11967, n11968, n11969, n11970, n11971, n11972, n11973, 
      n11974, n11975, n11976, n11977, n11978, n11979, n11980, n11981, n11982, 
      n11983, n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991, 
      n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000, 
      n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009, 
      n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017, n12018, 
      n12019, n12020, n12021, n12022, n12023, n12024, n12025, n12026, n12027, 
      n12028, n12029, n12030, n12031, n12032, n12033, n12034, n12035, n12036, 
      n12037, n12038, n12039, n12040, n12041, n12042, n12043, n12044, n12045, 
      n12046, n12047, n12048, n12049, n12050, n12051, n12052, n12053, n12054, 
      n12055, n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063, 
      n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072, 
      n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081, 
      n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089, n12090, 
      n12091, n12092, n12093, n12094, n12095, n12096, n12097, n12098, n12099, 
      n12100, n12101, n12102, n12103, n12104, n12105, n12106, n12107, n12108, 
      n12109, n12110, n12111, n12112, n12113, n12114, n12115, n12116, n12117, 
      n12118, n12119, n12120, n12121, n12122, n12123, n12124, n12125, n12126, 
      n12127, n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135, 
      n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144, 
      n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153, 
      n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161, n12162, 
      n12163, n12164, n12165, n12166, n12167, n12168, n12169, n12170, n12171, 
      n12172, n12173, n12174, n12175, n12176, n12177, n12178, n12179, n12180, 
      n12181, n12182, n12183, n12184, n12185, n12186, n12187, n12188, n12189, 
      n12190, n12191, n12192, n12193, n12194, n12195, n12196, n12197, n12198, 
      n12199, n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207, 
      n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216, 
      n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225, 
      n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233, n12234, 
      n12235, n12236, n12237, n12238, n12239, n12240, n12241, n12242, n12243, 
      n12244, n12245, n12246, n12247, n12248, n12249, n12250, n12251, n12252, 
      n12253, n12254, n12255, n12256, n12257, n12258, n12259, n12260, n12261, 
      n12262, n12263, n12264, n12265, n12266, n12267, n12268, n12269, n12270, 
      n12271, n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279, 
      n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288, 
      n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297, 
      n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305, n12306, 
      n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314, n12315, 
      n12316, n12317, n12318, n12319, n12320, n12321, n12322, n12323, n12324, 
      n12325, n12326, n12327, n12328, n12329, n12330, n12331, n12332, n12333, 
      n12334, n12335, n12336, n12337, n12338, n12339, n12340, n12341, n12342, 
      n12343, n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351, 
      n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360, 
      n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369, 
      n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377, n12378, 
      n12379, n12380, n12381, n12382, n12383, n12384, n12385, n12386, n12387, 
      n12388, n12389, n12390, n12391, n12392, n12393, n12394, n12395, n12396, 
      n12397, n12398, n12399, n12400, n12401, n12402, n12403, n12404, n12405, 
      n12406, n12407, n12408, n12409, n12410, n12411, n12412, n12413, n12414, 
      n12415, n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423, 
      n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432, 
      n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441, 
      n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449, n12450, 
      n12451, n12452, n12453, n12454, n12455, n12456, n12457, n12458, n12459, 
      n12460, n12461, n12462, n12463, n12464, n12465, n12466, n12467, n12468, 
      n12469, n12470, n12471, n12472, n12473, n12474, n12475, n12476, n12477, 
      n12478, n12479, n12480, n12481, n12482, n12483, n12484, n12485, n12486, 
      n12487, n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495, 
      n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504, 
      n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513, 
      n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521, n12522, 
      n12523, n12524, n_1000, n_1001, n_1002, n_1003, n_1004, n_1005, n_1006, 
      n_1007, n_1008, n_1009, n_1010, n_1011, n_1012, n_1013, n_1014, n_1015, 
      n_1016, n_1017, n_1018, n_1019, n_1020, n_1021, n_1022, n_1023, n_1024, 
      n_1025, n_1026, n_1027, n_1028, n_1029, n_1030, n_1031, n_1032, n_1033, 
      n_1034, n_1035, n_1036, n_1037, n_1038, n_1039, n_1040, n_1041, n_1042, 
      n_1043, n_1044, n_1045, n_1046, n_1047, n_1048, n_1049, n_1050, n_1051, 
      n_1052, n_1053, n_1054, n_1055, n_1056, n_1057, n_1058, n_1059, n_1060, 
      n_1061, n_1062, n_1063, n_1064, n_1065, n_1066, n_1067, n_1068, n_1069, 
      n_1070, n_1071, n_1072, n_1073, n_1074, n_1075, n_1076, n_1077, n_1078, 
      n_1079, n_1080, n_1081, n_1082, n_1083, n_1084, n_1085, n_1086, n_1087, 
      n_1088, n_1089, n_1090, n_1091, n_1092, n_1093, n_1094, n_1095, n_1096, 
      n_1097, n_1098, n_1099, n_1100, n_1101, n_1102, n_1103, n_1104, n_1105, 
      n_1106, n_1107, n_1108, n_1109, n_1110, n_1111, n_1112, n_1113, n_1114, 
      n_1115, n_1116, n_1117, n_1118, n_1119, n_1120, n_1121, n_1122, n_1123, 
      n_1124, n_1125, n_1126, n_1127, n_1128, n_1129, n_1130, n_1131, n_1132, 
      n_1133, n_1134, n_1135, n_1136, n_1137, n_1138, n_1139, n_1140, n_1141, 
      n_1142, n_1143, n_1144, n_1145, n_1146, n_1147, n_1148, n_1149, n_1150, 
      n_1151, n_1152, n_1153, n_1154, n_1155, n_1156, n_1157, n_1158, n_1159, 
      n_1160, n_1161, n_1162, n_1163, n_1164, n_1165, n_1166, n_1167, n_1168, 
      n_1169, n_1170, n_1171, n_1172, n_1173, n_1174, n_1175, n_1176, n_1177, 
      n_1178, n_1179, n_1180, n_1181, n_1182, n_1183, n_1184, n_1185, n_1186, 
      n_1187, n_1188, n_1189, n_1190, n_1191, n_1192, n_1193, n_1194, n_1195, 
      n_1196, n_1197, n_1198, n_1199, n_1200, n_1201, n_1202, n_1203, n_1204, 
      n_1205, n_1206, n_1207, n_1208, n_1209, n_1210, n_1211, n_1212, n_1213, 
      n_1214, n_1215, n_1216, n_1217, n_1218, n_1219, n_1220, n_1221, n_1222, 
      n_1223, n_1224, n_1225, n_1226, n_1227, n_1228, n_1229, n_1230, n_1231, 
      n_1232, n_1233, n_1234, n_1235, n_1236, n_1237, n_1238, n_1239, n_1240, 
      n_1241, n_1242, n_1243, n_1244, n_1245, n_1246, n_1247, n_1248, n_1249, 
      n_1250, n_1251, n_1252, n_1253, n_1254, n_1255, n_1256, n_1257, n_1258, 
      n_1259, n_1260, n_1261, n_1262, n_1263, n_1264, n_1265, n_1266, n_1267, 
      n_1268, n_1269, n_1270, n_1271, n_1272, n_1273, n_1274, n_1275, n_1276, 
      n_1277, n_1278, n_1279, n_1280, n_1281, n_1282, n_1283, n_1284, n_1285, 
      n_1286, n_1287, n_1288, n_1289, n_1290, n_1291, n_1292, n_1293, n_1294, 
      n_1295, n_1296, n_1297, n_1298, n_1299, n_1300, n_1301, n_1302, n_1303, 
      n_1304, n_1305, n_1306, n_1307, n_1308, n_1309, n_1310, n_1311, n_1312, 
      n_1313, n_1314, n_1315, n_1316, n_1317, n_1318, n_1319, n_1320, n_1321, 
      n_1322, n_1323, n_1324, n_1325, n_1326, n_1327, n_1328, n_1329, n_1330, 
      n_1331, n_1332, n_1333, n_1334, n_1335, n_1336, n_1337, n_1338, n_1339, 
      n_1340, n_1341, n_1342, n_1343, n_1344, n_1345, n_1346, n_1347, n_1348, 
      n_1349, n_1350, n_1351, n_1352, n_1353, n_1354, n_1355, n_1356, n_1357, 
      n_1358, n_1359, n_1360, n_1361, n_1362, n_1363, n_1364, n_1365, n_1366, 
      n_1367, n_1368, n_1369, n_1370, n_1371, n_1372, n_1373, n_1374, n_1375, 
      n_1376, n_1377, n_1378, n_1379, n_1380, n_1381, n_1382, n_1383, n_1384, 
      n_1385, n_1386, n_1387, n_1388, n_1389, n_1390, n_1391, n_1392, n_1393, 
      n_1394, n_1395, n_1396, n_1397, n_1398, n_1399, n_1400, n_1401, n_1402, 
      n_1403, n_1404, n_1405, n_1406, n_1407, n_1408, n_1409, n_1410, n_1411, 
      n_1412, n_1413, n_1414, n_1415, n_1416, n_1417, n_1418, n_1419, n_1420, 
      n_1421, n_1422, n_1423, n_1424, n_1425, n_1426, n_1427, n_1428, n_1429, 
      n_1430, n_1431, n_1432, n_1433, n_1434, n_1435, n_1436, n_1437, n_1438, 
      n_1439, n_1440, n_1441, n_1442, n_1443, n_1444, n_1445, n_1446, n_1447, 
      n_1448, n_1449, n_1450, n_1451, n_1452, n_1453, n_1454, n_1455, n_1456, 
      n_1457, n_1458, n_1459, n_1460, n_1461, n_1462, n_1463, n_1464, n_1465, 
      n_1466, n_1467, n_1468, n_1469, n_1470, n_1471, n_1472, n_1473, n_1474, 
      n_1475, n_1476, n_1477, n_1478, n_1479, n_1480, n_1481, n_1482, n_1483, 
      n_1484, n_1485, n_1486, n_1487, n_1488, n_1489, n_1490, n_1491, n_1492, 
      n_1493, n_1494, n_1495, n_1496, n_1497, n_1498, n_1499, n_1500, n_1501, 
      n_1502, n_1503, n_1504, n_1505, n_1506, n_1507, n_1508, n_1509, n_1510, 
      n_1511 : std_logic;

begin
   
   OUT1_reg_31_inst : DFF_X1 port map( D => n1610, CK => CLK, Q => n11163, QN 
                           => n4869);
   OUT1_tri_enable_reg_31_inst : DFF_X1 port map( D => n1609, CK => CLK, Q => 
                           n4870, QN => n4868);
   OUT1_reg_30_inst : DFF_X1 port map( D => n1608, CK => CLK, Q => n11162, QN 
                           => n4867);
   OUT1_tri_enable_reg_30_inst : DFF_X1 port map( D => n1607, CK => CLK, Q => 
                           n4871, QN => n4866);
   OUT1_reg_29_inst : DFF_X1 port map( D => n1606, CK => CLK, Q => n11161, QN 
                           => n4865);
   OUT1_tri_enable_reg_29_inst : DFF_X1 port map( D => n1605, CK => CLK, Q => 
                           n4872, QN => n4864);
   OUT1_reg_28_inst : DFF_X1 port map( D => n1604, CK => CLK, Q => n11160, QN 
                           => n4863);
   OUT1_tri_enable_reg_28_inst : DFF_X1 port map( D => n1603, CK => CLK, Q => 
                           n4873, QN => n4862);
   OUT1_reg_27_inst : DFF_X1 port map( D => n1602, CK => CLK, Q => n11159, QN 
                           => n4861);
   OUT1_tri_enable_reg_27_inst : DFF_X1 port map( D => n1601, CK => CLK, Q => 
                           n4874, QN => n4860);
   OUT1_reg_26_inst : DFF_X1 port map( D => n1600, CK => CLK, Q => n11158, QN 
                           => n4859);
   OUT1_tri_enable_reg_26_inst : DFF_X1 port map( D => n1599, CK => CLK, Q => 
                           n4875, QN => n4858);
   OUT1_reg_25_inst : DFF_X1 port map( D => n1598, CK => CLK, Q => n11157, QN 
                           => n4857);
   OUT1_tri_enable_reg_25_inst : DFF_X1 port map( D => n1597, CK => CLK, Q => 
                           n4876, QN => n4856);
   OUT1_reg_24_inst : DFF_X1 port map( D => n1596, CK => CLK, Q => n11156, QN 
                           => n4855);
   OUT1_tri_enable_reg_24_inst : DFF_X1 port map( D => n1595, CK => CLK, Q => 
                           n4877, QN => n4854);
   OUT1_reg_23_inst : DFF_X1 port map( D => n1594, CK => CLK, Q => n11155, QN 
                           => n4853);
   OUT1_tri_enable_reg_23_inst : DFF_X1 port map( D => n1593, CK => CLK, Q => 
                           n4878, QN => n4852);
   OUT1_reg_22_inst : DFF_X1 port map( D => n1592, CK => CLK, Q => n11154, QN 
                           => n4851);
   OUT1_tri_enable_reg_22_inst : DFF_X1 port map( D => n1591, CK => CLK, Q => 
                           n4879, QN => n4850);
   OUT1_reg_21_inst : DFF_X1 port map( D => n1590, CK => CLK, Q => n11153, QN 
                           => n4849);
   OUT1_tri_enable_reg_21_inst : DFF_X1 port map( D => n1589, CK => CLK, Q => 
                           n4880, QN => n4848);
   OUT1_reg_20_inst : DFF_X1 port map( D => n1588, CK => CLK, Q => n11152, QN 
                           => n4847);
   OUT1_tri_enable_reg_20_inst : DFF_X1 port map( D => n1587, CK => CLK, Q => 
                           n4881, QN => n4846);
   OUT1_reg_19_inst : DFF_X1 port map( D => n1586, CK => CLK, Q => n11151, QN 
                           => n4845);
   OUT1_tri_enable_reg_19_inst : DFF_X1 port map( D => n1585, CK => CLK, Q => 
                           n4882, QN => n4844);
   OUT1_reg_18_inst : DFF_X1 port map( D => n1584, CK => CLK, Q => n11150, QN 
                           => n4843);
   OUT1_tri_enable_reg_18_inst : DFF_X1 port map( D => n1583, CK => CLK, Q => 
                           n4883, QN => n4842);
   OUT1_reg_17_inst : DFF_X1 port map( D => n1582, CK => CLK, Q => n11149, QN 
                           => n4841);
   OUT1_tri_enable_reg_17_inst : DFF_X1 port map( D => n1581, CK => CLK, Q => 
                           n4884, QN => n4840);
   OUT1_reg_16_inst : DFF_X1 port map( D => n1580, CK => CLK, Q => n11148, QN 
                           => n4839);
   OUT1_tri_enable_reg_16_inst : DFF_X1 port map( D => n1579, CK => CLK, Q => 
                           n4885, QN => n4838);
   OUT1_reg_15_inst : DFF_X1 port map( D => n1578, CK => CLK, Q => n11147, QN 
                           => n4837);
   OUT1_tri_enable_reg_15_inst : DFF_X1 port map( D => n1577, CK => CLK, Q => 
                           n4886, QN => n4836);
   OUT1_reg_14_inst : DFF_X1 port map( D => n1576, CK => CLK, Q => n11146, QN 
                           => n4835);
   OUT1_tri_enable_reg_14_inst : DFF_X1 port map( D => n1575, CK => CLK, Q => 
                           n4887, QN => n4834);
   OUT1_reg_13_inst : DFF_X1 port map( D => n1574, CK => CLK, Q => n11145, QN 
                           => n4833);
   OUT1_tri_enable_reg_13_inst : DFF_X1 port map( D => n1573, CK => CLK, Q => 
                           n4888, QN => n4832);
   OUT1_reg_12_inst : DFF_X1 port map( D => n1572, CK => CLK, Q => n11144, QN 
                           => n4831);
   OUT1_tri_enable_reg_12_inst : DFF_X1 port map( D => n1571, CK => CLK, Q => 
                           n4889, QN => n4830);
   OUT1_reg_11_inst : DFF_X1 port map( D => n1570, CK => CLK, Q => n11143, QN 
                           => n4829);
   OUT1_tri_enable_reg_11_inst : DFF_X1 port map( D => n1569, CK => CLK, Q => 
                           n4890, QN => n4828);
   OUT1_reg_10_inst : DFF_X1 port map( D => n1568, CK => CLK, Q => n11142, QN 
                           => n4827);
   OUT1_tri_enable_reg_10_inst : DFF_X1 port map( D => n1567, CK => CLK, Q => 
                           n4891, QN => n4826);
   OUT1_reg_9_inst : DFF_X1 port map( D => n1566, CK => CLK, Q => n11141, QN =>
                           n4825);
   OUT1_tri_enable_reg_9_inst : DFF_X1 port map( D => n1565, CK => CLK, Q => 
                           n4892, QN => n4824);
   OUT1_reg_8_inst : DFF_X1 port map( D => n1564, CK => CLK, Q => n11140, QN =>
                           n4823);
   OUT1_tri_enable_reg_8_inst : DFF_X1 port map( D => n1563, CK => CLK, Q => 
                           n4893, QN => n4822);
   OUT1_reg_7_inst : DFF_X1 port map( D => n1562, CK => CLK, Q => n11139, QN =>
                           n4821);
   OUT1_tri_enable_reg_7_inst : DFF_X1 port map( D => n1561, CK => CLK, Q => 
                           n4894, QN => n4820);
   OUT1_reg_6_inst : DFF_X1 port map( D => n1560, CK => CLK, Q => n11138, QN =>
                           n4819);
   OUT1_tri_enable_reg_6_inst : DFF_X1 port map( D => n1559, CK => CLK, Q => 
                           n4895, QN => n4818);
   OUT1_reg_5_inst : DFF_X1 port map( D => n1558, CK => CLK, Q => n11137, QN =>
                           n4817);
   OUT1_tri_enable_reg_5_inst : DFF_X1 port map( D => n1557, CK => CLK, Q => 
                           n4896, QN => n4816);
   OUT1_reg_4_inst : DFF_X1 port map( D => n1556, CK => CLK, Q => n11136, QN =>
                           n4815);
   OUT1_tri_enable_reg_4_inst : DFF_X1 port map( D => n1555, CK => CLK, Q => 
                           n4897, QN => n4814);
   OUT1_reg_3_inst : DFF_X1 port map( D => n1554, CK => CLK, Q => n11135, QN =>
                           n4813);
   OUT1_tri_enable_reg_3_inst : DFF_X1 port map( D => n1553, CK => CLK, Q => 
                           n4898, QN => n4812);
   OUT1_reg_2_inst : DFF_X1 port map( D => n1552, CK => CLK, Q => n11134, QN =>
                           n4811);
   OUT1_tri_enable_reg_2_inst : DFF_X1 port map( D => n1551, CK => CLK, Q => 
                           n4899, QN => n4810);
   OUT1_reg_1_inst : DFF_X1 port map( D => n1550, CK => CLK, Q => n11133, QN =>
                           n4809);
   OUT1_tri_enable_reg_1_inst : DFF_X1 port map( D => n1549, CK => CLK, Q => 
                           n4900, QN => n4808);
   OUT1_reg_0_inst : DFF_X1 port map( D => n1548, CK => CLK, Q => n11132, QN =>
                           n4807);
   OUT1_tri_enable_reg_0_inst : DFF_X1 port map( D => n1547, CK => CLK, Q => 
                           n4901, QN => n4806);
   OUT2_reg_31_inst : DFF_X1 port map( D => n1546, CK => CLK, Q => n11131, QN 
                           => n4805);
   OUT2_tri_enable_reg_31_inst : DFF_X1 port map( D => n1545, CK => CLK, Q => 
                           n4902, QN => n4804);
   OUT2_reg_30_inst : DFF_X1 port map( D => n1544, CK => CLK, Q => n11130, QN 
                           => n4803);
   OUT2_tri_enable_reg_30_inst : DFF_X1 port map( D => n1543, CK => CLK, Q => 
                           n4903, QN => n4802);
   OUT2_reg_29_inst : DFF_X1 port map( D => n1542, CK => CLK, Q => n11129, QN 
                           => n4801);
   OUT2_tri_enable_reg_29_inst : DFF_X1 port map( D => n1541, CK => CLK, Q => 
                           n4904, QN => n4800);
   OUT2_reg_28_inst : DFF_X1 port map( D => n1540, CK => CLK, Q => n11128, QN 
                           => n4799);
   OUT2_tri_enable_reg_28_inst : DFF_X1 port map( D => n1539, CK => CLK, Q => 
                           n4905, QN => n4798);
   OUT2_reg_27_inst : DFF_X1 port map( D => n1538, CK => CLK, Q => n11127, QN 
                           => n4797);
   OUT2_tri_enable_reg_27_inst : DFF_X1 port map( D => n1537, CK => CLK, Q => 
                           n4906, QN => n4796);
   OUT2_reg_26_inst : DFF_X1 port map( D => n1536, CK => CLK, Q => n11126, QN 
                           => n4795);
   OUT2_tri_enable_reg_26_inst : DFF_X1 port map( D => n1535, CK => CLK, Q => 
                           n4907, QN => n4794);
   OUT2_reg_25_inst : DFF_X1 port map( D => n1534, CK => CLK, Q => n11125, QN 
                           => n4793);
   OUT2_tri_enable_reg_25_inst : DFF_X1 port map( D => n1533, CK => CLK, Q => 
                           n4908, QN => n4792);
   OUT2_reg_24_inst : DFF_X1 port map( D => n1532, CK => CLK, Q => n11124, QN 
                           => n4791);
   OUT2_tri_enable_reg_24_inst : DFF_X1 port map( D => n1531, CK => CLK, Q => 
                           n4909, QN => n4790);
   OUT2_reg_23_inst : DFF_X1 port map( D => n1530, CK => CLK, Q => n11123, QN 
                           => n4789);
   OUT2_tri_enable_reg_23_inst : DFF_X1 port map( D => n1529, CK => CLK, Q => 
                           n4910, QN => n4788);
   OUT2_reg_22_inst : DFF_X1 port map( D => n1528, CK => CLK, Q => n11122, QN 
                           => n4787);
   OUT2_tri_enable_reg_22_inst : DFF_X1 port map( D => n1527, CK => CLK, Q => 
                           n4911, QN => n4786);
   OUT2_reg_21_inst : DFF_X1 port map( D => n1526, CK => CLK, Q => n11121, QN 
                           => n4785);
   OUT2_tri_enable_reg_21_inst : DFF_X1 port map( D => n1525, CK => CLK, Q => 
                           n4912, QN => n4784);
   OUT2_reg_20_inst : DFF_X1 port map( D => n1524, CK => CLK, Q => n11120, QN 
                           => n4783);
   OUT2_tri_enable_reg_20_inst : DFF_X1 port map( D => n1523, CK => CLK, Q => 
                           n4913, QN => n4782);
   OUT2_reg_19_inst : DFF_X1 port map( D => n1522, CK => CLK, Q => n11119, QN 
                           => n4781);
   OUT2_tri_enable_reg_19_inst : DFF_X1 port map( D => n1521, CK => CLK, Q => 
                           n4914, QN => n4780);
   OUT2_reg_18_inst : DFF_X1 port map( D => n1520, CK => CLK, Q => n11118, QN 
                           => n4779);
   OUT2_tri_enable_reg_18_inst : DFF_X1 port map( D => n1519, CK => CLK, Q => 
                           n4915, QN => n4778);
   OUT2_reg_17_inst : DFF_X1 port map( D => n1518, CK => CLK, Q => n11117, QN 
                           => n4777);
   OUT2_tri_enable_reg_17_inst : DFF_X1 port map( D => n1517, CK => CLK, Q => 
                           n4916, QN => n4776);
   OUT2_reg_16_inst : DFF_X1 port map( D => n1516, CK => CLK, Q => n11116, QN 
                           => n4775);
   OUT2_tri_enable_reg_16_inst : DFF_X1 port map( D => n1515, CK => CLK, Q => 
                           n4917, QN => n4774);
   OUT2_reg_15_inst : DFF_X1 port map( D => n1514, CK => CLK, Q => n11115, QN 
                           => n4773);
   OUT2_tri_enable_reg_15_inst : DFF_X1 port map( D => n1513, CK => CLK, Q => 
                           n4918, QN => n4772);
   OUT2_reg_14_inst : DFF_X1 port map( D => n1512, CK => CLK, Q => n11114, QN 
                           => n4771);
   OUT2_tri_enable_reg_14_inst : DFF_X1 port map( D => n1511, CK => CLK, Q => 
                           n4919, QN => n4770);
   OUT2_reg_13_inst : DFF_X1 port map( D => n1510, CK => CLK, Q => n11113, QN 
                           => n4769);
   OUT2_tri_enable_reg_13_inst : DFF_X1 port map( D => n1509, CK => CLK, Q => 
                           n4920, QN => n4768);
   OUT2_reg_12_inst : DFF_X1 port map( D => n1508, CK => CLK, Q => n11112, QN 
                           => n4767);
   OUT2_tri_enable_reg_12_inst : DFF_X1 port map( D => n1507, CK => CLK, Q => 
                           n4921, QN => n4766);
   OUT2_reg_11_inst : DFF_X1 port map( D => n1506, CK => CLK, Q => n11111, QN 
                           => n4765);
   OUT2_tri_enable_reg_11_inst : DFF_X1 port map( D => n1505, CK => CLK, Q => 
                           n4922, QN => n4764);
   OUT2_reg_10_inst : DFF_X1 port map( D => n1504, CK => CLK, Q => n11110, QN 
                           => n4763);
   OUT2_tri_enable_reg_10_inst : DFF_X1 port map( D => n1503, CK => CLK, Q => 
                           n4923, QN => n4762);
   OUT2_reg_9_inst : DFF_X1 port map( D => n1502, CK => CLK, Q => n11109, QN =>
                           n4761);
   OUT2_tri_enable_reg_9_inst : DFF_X1 port map( D => n1501, CK => CLK, Q => 
                           n4924, QN => n4760);
   OUT2_reg_8_inst : DFF_X1 port map( D => n1500, CK => CLK, Q => n11108, QN =>
                           n4759);
   OUT2_tri_enable_reg_8_inst : DFF_X1 port map( D => n1499, CK => CLK, Q => 
                           n4925, QN => n4758);
   OUT2_reg_7_inst : DFF_X1 port map( D => n1498, CK => CLK, Q => n11107, QN =>
                           n4757);
   OUT2_tri_enable_reg_7_inst : DFF_X1 port map( D => n1497, CK => CLK, Q => 
                           n4926, QN => n4756);
   OUT2_reg_6_inst : DFF_X1 port map( D => n1496, CK => CLK, Q => n11106, QN =>
                           n4755);
   OUT2_tri_enable_reg_6_inst : DFF_X1 port map( D => n1495, CK => CLK, Q => 
                           n4927, QN => n4754);
   OUT2_reg_5_inst : DFF_X1 port map( D => n1494, CK => CLK, Q => n11105, QN =>
                           n4753);
   OUT2_tri_enable_reg_5_inst : DFF_X1 port map( D => n1493, CK => CLK, Q => 
                           n4928, QN => n4752);
   OUT2_reg_4_inst : DFF_X1 port map( D => n1492, CK => CLK, Q => n11104, QN =>
                           n4751);
   OUT2_tri_enable_reg_4_inst : DFF_X1 port map( D => n1491, CK => CLK, Q => 
                           n4929, QN => n4750);
   OUT2_reg_3_inst : DFF_X1 port map( D => n1490, CK => CLK, Q => n11103, QN =>
                           n4749);
   OUT2_tri_enable_reg_3_inst : DFF_X1 port map( D => n1489, CK => CLK, Q => 
                           n4930, QN => n4748);
   OUT2_reg_2_inst : DFF_X1 port map( D => n1488, CK => CLK, Q => n11102, QN =>
                           n4747);
   OUT2_tri_enable_reg_2_inst : DFF_X1 port map( D => n1487, CK => CLK, Q => 
                           n4931, QN => n4746);
   OUT2_reg_1_inst : DFF_X1 port map( D => n1486, CK => CLK, Q => n11101, QN =>
                           n4745);
   OUT2_tri_enable_reg_1_inst : DFF_X1 port map( D => n1485, CK => CLK, Q => 
                           n4932, QN => n4744);
   OUT2_reg_0_inst : DFF_X1 port map( D => n1484, CK => CLK, Q => n11100, QN =>
                           n4743);
   OUT2_tri_enable_reg_0_inst : DFF_X1 port map( D => n1483, CK => CLK, Q => 
                           n4933, QN => n4742);
   U1645 : TINV_X1 port map( I => n4869, EN => n4870, ZN => OUT1(31));
   U1646 : TINV_X1 port map( I => n4867, EN => n4871, ZN => OUT1(30));
   U1647 : TINV_X1 port map( I => n4865, EN => n4872, ZN => OUT1(29));
   U1648 : TINV_X1 port map( I => n4863, EN => n4873, ZN => OUT1(28));
   U1649 : TINV_X1 port map( I => n4861, EN => n4874, ZN => OUT1(27));
   U1650 : TINV_X1 port map( I => n4859, EN => n4875, ZN => OUT1(26));
   U1651 : TINV_X1 port map( I => n4857, EN => n4876, ZN => OUT1(25));
   U1652 : TINV_X1 port map( I => n4855, EN => n4877, ZN => OUT1(24));
   U1653 : TINV_X1 port map( I => n4853, EN => n4878, ZN => OUT1(23));
   U1654 : TINV_X1 port map( I => n4851, EN => n4879, ZN => OUT1(22));
   U1655 : TINV_X1 port map( I => n4849, EN => n4880, ZN => OUT1(21));
   U1656 : TINV_X1 port map( I => n4847, EN => n4881, ZN => OUT1(20));
   U1657 : TINV_X1 port map( I => n4845, EN => n4882, ZN => OUT1(19));
   U1658 : TINV_X1 port map( I => n4843, EN => n4883, ZN => OUT1(18));
   U1659 : TINV_X1 port map( I => n4841, EN => n4884, ZN => OUT1(17));
   U1660 : TINV_X1 port map( I => n4839, EN => n4885, ZN => OUT1(16));
   U1661 : TINV_X1 port map( I => n4837, EN => n4886, ZN => OUT1(15));
   U1662 : TINV_X1 port map( I => n4835, EN => n4887, ZN => OUT1(14));
   U1663 : TINV_X1 port map( I => n4833, EN => n4888, ZN => OUT1(13));
   U1664 : TINV_X1 port map( I => n4831, EN => n4889, ZN => OUT1(12));
   U1665 : TINV_X1 port map( I => n4829, EN => n4890, ZN => OUT1(11));
   U1666 : TINV_X1 port map( I => n4827, EN => n4891, ZN => OUT1(10));
   U1667 : TINV_X1 port map( I => n4825, EN => n4892, ZN => OUT1(9));
   U1668 : TINV_X1 port map( I => n4823, EN => n4893, ZN => OUT1(8));
   U1669 : TINV_X1 port map( I => n4821, EN => n4894, ZN => OUT1(7));
   U1670 : TINV_X1 port map( I => n4819, EN => n4895, ZN => OUT1(6));
   U1671 : TINV_X1 port map( I => n4817, EN => n4896, ZN => OUT1(5));
   U1672 : TINV_X1 port map( I => n4815, EN => n4897, ZN => OUT1(4));
   U1673 : TINV_X1 port map( I => n4813, EN => n4898, ZN => OUT1(3));
   U1674 : TINV_X1 port map( I => n4811, EN => n4899, ZN => OUT1(2));
   U1675 : TINV_X1 port map( I => n4809, EN => n4900, ZN => OUT1(1));
   U1676 : TINV_X1 port map( I => n4807, EN => n4901, ZN => OUT1(0));
   U1677 : TINV_X1 port map( I => n4805, EN => n4902, ZN => OUT2(31));
   U1678 : TINV_X1 port map( I => n4803, EN => n4903, ZN => OUT2(30));
   U1679 : TINV_X1 port map( I => n4801, EN => n4904, ZN => OUT2(29));
   U1680 : TINV_X1 port map( I => n4799, EN => n4905, ZN => OUT2(28));
   U1681 : TINV_X1 port map( I => n4797, EN => n4906, ZN => OUT2(27));
   U1682 : TINV_X1 port map( I => n4795, EN => n4907, ZN => OUT2(26));
   U1683 : TINV_X1 port map( I => n4793, EN => n4908, ZN => OUT2(25));
   U1684 : TINV_X1 port map( I => n4791, EN => n4909, ZN => OUT2(24));
   U1685 : TINV_X1 port map( I => n4789, EN => n4910, ZN => OUT2(23));
   U1686 : TINV_X1 port map( I => n4787, EN => n4911, ZN => OUT2(22));
   U1687 : TINV_X1 port map( I => n4785, EN => n4912, ZN => OUT2(21));
   U1688 : TINV_X1 port map( I => n4783, EN => n4913, ZN => OUT2(20));
   U1689 : TINV_X1 port map( I => n4781, EN => n4914, ZN => OUT2(19));
   U1690 : TINV_X1 port map( I => n4779, EN => n4915, ZN => OUT2(18));
   U1691 : TINV_X1 port map( I => n4777, EN => n4916, ZN => OUT2(17));
   U1692 : TINV_X1 port map( I => n4775, EN => n4917, ZN => OUT2(16));
   U1693 : TINV_X1 port map( I => n4773, EN => n4918, ZN => OUT2(15));
   U1694 : TINV_X1 port map( I => n4771, EN => n4919, ZN => OUT2(14));
   U1695 : TINV_X1 port map( I => n4769, EN => n4920, ZN => OUT2(13));
   U1696 : TINV_X1 port map( I => n4767, EN => n4921, ZN => OUT2(12));
   U1697 : TINV_X1 port map( I => n4765, EN => n4922, ZN => OUT2(11));
   U1698 : TINV_X1 port map( I => n4763, EN => n4923, ZN => OUT2(10));
   U1699 : TINV_X1 port map( I => n4761, EN => n4924, ZN => OUT2(9));
   U1700 : TINV_X1 port map( I => n4759, EN => n4925, ZN => OUT2(8));
   U1701 : TINV_X1 port map( I => n4757, EN => n4926, ZN => OUT2(7));
   U1702 : TINV_X1 port map( I => n4755, EN => n4927, ZN => OUT2(6));
   U1703 : TINV_X1 port map( I => n4753, EN => n4928, ZN => OUT2(5));
   U1704 : TINV_X1 port map( I => n4751, EN => n4929, ZN => OUT2(4));
   U1705 : TINV_X1 port map( I => n4749, EN => n4930, ZN => OUT2(3));
   U1706 : TINV_X1 port map( I => n4747, EN => n4931, ZN => OUT2(2));
   U1707 : TINV_X1 port map( I => n4745, EN => n4932, ZN => OUT2(1));
   U1708 : TINV_X1 port map( I => n4743, EN => n4933, ZN => OUT2(0));
   U7967 : NAND3_X1 port map( A1 => n8785, A2 => n8784, A3 => n9863, ZN => 
                           n9855);
   U7968 : NAND3_X1 port map( A1 => n9863, A2 => n8784, A3 => ADD_WR(2), ZN => 
                           n9865);
   U7969 : NAND3_X1 port map( A1 => n9863, A2 => n8785, A3 => ADD_WR(3), ZN => 
                           n9870);
   U7970 : NAND3_X1 port map( A1 => ADD_WR(2), A2 => n9863, A3 => ADD_WR(3), ZN
                           => n9875);
   U7971 : NAND3_X1 port map( A1 => n8785, A2 => n8784, A3 => n9884, ZN => 
                           n9880);
   U7972 : NAND3_X1 port map( A1 => ADD_WR(2), A2 => n8784, A3 => n9884, ZN => 
                           n9886);
   U7973 : NAND3_X1 port map( A1 => ADD_WR(3), A2 => n8785, A3 => n9884, ZN => 
                           n9891);
   U7974 : NAND3_X1 port map( A1 => ADD_WR(3), A2 => ADD_WR(2), A3 => n9884, ZN
                           => n9896);
   U7975 : NAND3_X1 port map( A1 => n10468, A2 => n12199, A3 => n10469, ZN => 
                           n9909);
   U7976 : NAND3_X1 port map( A1 => n10468, A2 => n12199, A3 => n10470, ZN => 
                           n9908);
   U7977 : NAND3_X1 port map( A1 => n10468, A2 => n12199, A3 => n10471, ZN => 
                           n9907);
   U7978 : NAND3_X1 port map( A1 => n10468, A2 => n12199, A3 => n10475, ZN => 
                           n9914);
   U7979 : NAND3_X1 port map( A1 => n10476, A2 => n12199, A3 => n10477, ZN => 
                           n9913);
   U7980 : NAND3_X1 port map( A1 => n10471, A2 => n12199, A3 => n10477, ZN => 
                           n9919);
   U7981 : NAND3_X1 port map( A1 => n10475, A2 => n12199, A3 => n10477, ZN => 
                           n9918);
   U7982 : NAND3_X1 port map( A1 => n10469, A2 => n12199, A3 => n10477, ZN => 
                           n9925);
   U7984 : XOR2_X1 port map( A => ADD_RD1(3), B => ADD_WR(3), Z => n10486);
   U7985 : XOR2_X1 port map( A => ADD_WR(1), B => ADD_RD1(1), Z => n10487);
   U7986 : XOR2_X1 port map( A => n8791, B => ADD_WR(2), Z => n10484);
   U7987 : NAND3_X1 port map( A1 => n11068, A2 => n12055, A3 => n11069, ZN => 
                           n10509);
   U7988 : NAND3_X1 port map( A1 => n11068, A2 => n12055, A3 => n11070, ZN => 
                           n10508);
   U7989 : NAND3_X1 port map( A1 => n11068, A2 => n12055, A3 => n11071, ZN => 
                           n10507);
   U7990 : NAND3_X1 port map( A1 => n11068, A2 => n12055, A3 => n11075, ZN => 
                           n10514);
   U7991 : NAND3_X1 port map( A1 => n11076, A2 => n12055, A3 => n11077, ZN => 
                           n10513);
   U7992 : NAND3_X1 port map( A1 => n11071, A2 => n12055, A3 => n11077, ZN => 
                           n10519);
   U7993 : NAND3_X1 port map( A1 => n11075, A2 => n12055, A3 => n11077, ZN => 
                           n10518);
   U7994 : NAND3_X1 port map( A1 => n11069, A2 => n12055, A3 => n11077, ZN => 
                           n10525);
   U7996 : XOR2_X1 port map( A => ADD_RD2(3), B => ADD_WR(3), Z => n11086);
   U7997 : XOR2_X1 port map( A => ADD_WR(1), B => ADD_RD2(1), Z => n11087);
   U7998 : XOR2_X1 port map( A => n8795, B => ADD_WR(2), Z => n11084);
   REGISTERS_reg_31_7_inst : DFF_X1 port map( D => n1618, CK => CLK, Q => 
                           n11843, QN => n9814);
   REGISTERS_reg_31_6_inst : DFF_X1 port map( D => n1617, CK => CLK, Q => 
                           n11842, QN => n9815);
   REGISTERS_reg_31_5_inst : DFF_X1 port map( D => n1616, CK => CLK, Q => 
                           n11841, QN => n9816);
   REGISTERS_reg_31_4_inst : DFF_X1 port map( D => n1615, CK => CLK, Q => 
                           n11840, QN => n9817);
   REGISTERS_reg_31_3_inst : DFF_X1 port map( D => n1614, CK => CLK, Q => 
                           n11839, QN => n9818);
   REGISTERS_reg_31_2_inst : DFF_X1 port map( D => n1613, CK => CLK, Q => 
                           n11838, QN => n9819);
   REGISTERS_reg_31_1_inst : DFF_X1 port map( D => n1612, CK => CLK, Q => 
                           n11837, QN => n9820);
   REGISTERS_reg_31_0_inst : DFF_X1 port map( D => n1611, CK => CLK, Q => 
                           n11516, QN => n9821);
   REGISTERS_reg_31_31_inst : DFF_X1 port map( D => n1642, CK => CLK, Q => 
                           n11867, QN => n9790);
   REGISTERS_reg_31_30_inst : DFF_X1 port map( D => n1641, CK => CLK, Q => 
                           n11866, QN => n9791);
   REGISTERS_reg_31_29_inst : DFF_X1 port map( D => n1640, CK => CLK, Q => 
                           n11865, QN => n9792);
   REGISTERS_reg_31_28_inst : DFF_X1 port map( D => n1639, CK => CLK, Q => 
                           n11864, QN => n9793);
   REGISTERS_reg_31_27_inst : DFF_X1 port map( D => n1638, CK => CLK, Q => 
                           n11863, QN => n9794);
   REGISTERS_reg_31_26_inst : DFF_X1 port map( D => n1637, CK => CLK, Q => 
                           n11862, QN => n9795);
   REGISTERS_reg_31_25_inst : DFF_X1 port map( D => n1636, CK => CLK, Q => 
                           n11861, QN => n9796);
   REGISTERS_reg_31_24_inst : DFF_X1 port map( D => n1635, CK => CLK, Q => 
                           n11860, QN => n9797);
   REGISTERS_reg_31_23_inst : DFF_X1 port map( D => n1634, CK => CLK, Q => 
                           n11859, QN => n9798);
   REGISTERS_reg_31_22_inst : DFF_X1 port map( D => n1633, CK => CLK, Q => 
                           n11858, QN => n9799);
   REGISTERS_reg_31_21_inst : DFF_X1 port map( D => n1632, CK => CLK, Q => 
                           n11857, QN => n9800);
   REGISTERS_reg_31_20_inst : DFF_X1 port map( D => n1631, CK => CLK, Q => 
                           n11856, QN => n9801);
   REGISTERS_reg_31_19_inst : DFF_X1 port map( D => n1630, CK => CLK, Q => 
                           n11855, QN => n9802);
   REGISTERS_reg_31_18_inst : DFF_X1 port map( D => n1629, CK => CLK, Q => 
                           n11854, QN => n9803);
   REGISTERS_reg_31_17_inst : DFF_X1 port map( D => n1628, CK => CLK, Q => 
                           n11853, QN => n9804);
   REGISTERS_reg_31_16_inst : DFF_X1 port map( D => n1627, CK => CLK, Q => 
                           n11852, QN => n9805);
   REGISTERS_reg_31_15_inst : DFF_X1 port map( D => n1626, CK => CLK, Q => 
                           n11851, QN => n9806);
   REGISTERS_reg_31_14_inst : DFF_X1 port map( D => n1625, CK => CLK, Q => 
                           n11850, QN => n9807);
   REGISTERS_reg_31_13_inst : DFF_X1 port map( D => n1624, CK => CLK, Q => 
                           n11849, QN => n9808);
   REGISTERS_reg_31_12_inst : DFF_X1 port map( D => n1623, CK => CLK, Q => 
                           n11848, QN => n9809);
   REGISTERS_reg_31_11_inst : DFF_X1 port map( D => n1622, CK => CLK, Q => 
                           n11847, QN => n9810);
   REGISTERS_reg_31_10_inst : DFF_X1 port map( D => n1621, CK => CLK, Q => 
                           n11846, QN => n9811);
   REGISTERS_reg_31_9_inst : DFF_X1 port map( D => n1620, CK => CLK, Q => 
                           n11845, QN => n9812);
   REGISTERS_reg_31_8_inst : DFF_X1 port map( D => n1619, CK => CLK, Q => 
                           n11844, QN => n9813);
   REGISTERS_reg_20_31_inst : DFF_X1 port map( D => n1994, CK => CLK, Q => 
                           n_1000, QN => n9438);
   REGISTERS_reg_20_30_inst : DFF_X1 port map( D => n1993, CK => CLK, Q => 
                           n_1001, QN => n9439);
   REGISTERS_reg_20_29_inst : DFF_X1 port map( D => n1992, CK => CLK, Q => 
                           n_1002, QN => n9440);
   REGISTERS_reg_20_28_inst : DFF_X1 port map( D => n1991, CK => CLK, Q => 
                           n_1003, QN => n9441);
   REGISTERS_reg_20_27_inst : DFF_X1 port map( D => n1990, CK => CLK, Q => 
                           n_1004, QN => n9442);
   REGISTERS_reg_20_26_inst : DFF_X1 port map( D => n1989, CK => CLK, Q => 
                           n_1005, QN => n9443);
   REGISTERS_reg_20_25_inst : DFF_X1 port map( D => n1988, CK => CLK, Q => 
                           n_1006, QN => n9444);
   REGISTERS_reg_20_24_inst : DFF_X1 port map( D => n1987, CK => CLK, Q => 
                           n_1007, QN => n9445);
   REGISTERS_reg_28_31_inst : DFF_X1 port map( D => n1738, CK => CLK, Q => 
                           n_1008, QN => n9694);
   REGISTERS_reg_28_30_inst : DFF_X1 port map( D => n1737, CK => CLK, Q => 
                           n_1009, QN => n9695);
   REGISTERS_reg_28_29_inst : DFF_X1 port map( D => n1736, CK => CLK, Q => 
                           n_1010, QN => n9696);
   REGISTERS_reg_28_28_inst : DFF_X1 port map( D => n1735, CK => CLK, Q => 
                           n_1011, QN => n9697);
   REGISTERS_reg_28_27_inst : DFF_X1 port map( D => n1734, CK => CLK, Q => 
                           n_1012, QN => n9698);
   REGISTERS_reg_28_26_inst : DFF_X1 port map( D => n1733, CK => CLK, Q => 
                           n_1013, QN => n9699);
   REGISTERS_reg_28_25_inst : DFF_X1 port map( D => n1732, CK => CLK, Q => 
                           n_1014, QN => n9700);
   REGISTERS_reg_28_24_inst : DFF_X1 port map( D => n1731, CK => CLK, Q => 
                           n_1015, QN => n9701);
   REGISTERS_reg_24_31_inst : DFF_X1 port map( D => n1866, CK => CLK, Q => 
                           n_1016, QN => n9566);
   REGISTERS_reg_24_30_inst : DFF_X1 port map( D => n1865, CK => CLK, Q => 
                           n_1017, QN => n9567);
   REGISTERS_reg_24_29_inst : DFF_X1 port map( D => n1864, CK => CLK, Q => 
                           n_1018, QN => n9568);
   REGISTERS_reg_24_28_inst : DFF_X1 port map( D => n1863, CK => CLK, Q => 
                           n_1019, QN => n9569);
   REGISTERS_reg_24_27_inst : DFF_X1 port map( D => n1862, CK => CLK, Q => 
                           n_1020, QN => n9570);
   REGISTERS_reg_24_26_inst : DFF_X1 port map( D => n1861, CK => CLK, Q => 
                           n_1021, QN => n9571);
   REGISTERS_reg_24_25_inst : DFF_X1 port map( D => n1860, CK => CLK, Q => 
                           n_1022, QN => n9572);
   REGISTERS_reg_24_24_inst : DFF_X1 port map( D => n1859, CK => CLK, Q => 
                           n_1023, QN => n9573);
   REGISTERS_reg_18_31_inst : DFF_X1 port map( D => n2058, CK => CLK, Q => 
                           n_1024, QN => n9374);
   REGISTERS_reg_18_30_inst : DFF_X1 port map( D => n2057, CK => CLK, Q => 
                           n_1025, QN => n9375);
   REGISTERS_reg_18_29_inst : DFF_X1 port map( D => n2056, CK => CLK, Q => 
                           n_1026, QN => n9376);
   REGISTERS_reg_18_28_inst : DFF_X1 port map( D => n2055, CK => CLK, Q => 
                           n_1027, QN => n9377);
   REGISTERS_reg_18_27_inst : DFF_X1 port map( D => n2054, CK => CLK, Q => 
                           n_1028, QN => n9378);
   REGISTERS_reg_18_26_inst : DFF_X1 port map( D => n2053, CK => CLK, Q => 
                           n_1029, QN => n9379);
   REGISTERS_reg_18_25_inst : DFF_X1 port map( D => n2052, CK => CLK, Q => 
                           n_1030, QN => n9380);
   REGISTERS_reg_18_24_inst : DFF_X1 port map( D => n2051, CK => CLK, Q => 
                           n_1031, QN => n9381);
   REGISTERS_reg_15_31_inst : DFF_X1 port map( D => n2154, CK => CLK, Q => 
                           n_1032, QN => n9278);
   REGISTERS_reg_15_30_inst : DFF_X1 port map( D => n2153, CK => CLK, Q => 
                           n_1033, QN => n9279);
   REGISTERS_reg_15_29_inst : DFF_X1 port map( D => n2152, CK => CLK, Q => 
                           n_1034, QN => n9280);
   REGISTERS_reg_15_28_inst : DFF_X1 port map( D => n2151, CK => CLK, Q => 
                           n_1035, QN => n9281);
   REGISTERS_reg_15_27_inst : DFF_X1 port map( D => n2150, CK => CLK, Q => 
                           n_1036, QN => n9282);
   REGISTERS_reg_15_26_inst : DFF_X1 port map( D => n2149, CK => CLK, Q => 
                           n_1037, QN => n9283);
   REGISTERS_reg_15_25_inst : DFF_X1 port map( D => n2148, CK => CLK, Q => 
                           n_1038, QN => n9284);
   REGISTERS_reg_15_24_inst : DFF_X1 port map( D => n2147, CK => CLK, Q => 
                           n_1039, QN => n9285);
   REGISTERS_reg_8_31_inst : DFF_X1 port map( D => n2378, CK => CLK, Q => 
                           n_1040, QN => n9054);
   REGISTERS_reg_8_30_inst : DFF_X1 port map( D => n2377, CK => CLK, Q => 
                           n_1041, QN => n9055);
   REGISTERS_reg_8_29_inst : DFF_X1 port map( D => n2376, CK => CLK, Q => 
                           n_1042, QN => n9056);
   REGISTERS_reg_8_28_inst : DFF_X1 port map( D => n2375, CK => CLK, Q => 
                           n_1043, QN => n9057);
   REGISTERS_reg_8_27_inst : DFF_X1 port map( D => n2374, CK => CLK, Q => 
                           n_1044, QN => n9058);
   REGISTERS_reg_8_26_inst : DFF_X1 port map( D => n2373, CK => CLK, Q => 
                           n_1045, QN => n9059);
   REGISTERS_reg_8_25_inst : DFF_X1 port map( D => n2372, CK => CLK, Q => 
                           n_1046, QN => n9060);
   REGISTERS_reg_8_24_inst : DFF_X1 port map( D => n2371, CK => CLK, Q => 
                           n_1047, QN => n9061);
   REGISTERS_reg_4_31_inst : DFF_X1 port map( D => n2506, CK => CLK, Q => 
                           n_1048, QN => n8926);
   REGISTERS_reg_4_30_inst : DFF_X1 port map( D => n2505, CK => CLK, Q => 
                           n_1049, QN => n8927);
   REGISTERS_reg_4_29_inst : DFF_X1 port map( D => n2504, CK => CLK, Q => 
                           n_1050, QN => n8928);
   REGISTERS_reg_4_28_inst : DFF_X1 port map( D => n2503, CK => CLK, Q => 
                           n_1051, QN => n8929);
   REGISTERS_reg_4_27_inst : DFF_X1 port map( D => n2502, CK => CLK, Q => 
                           n_1052, QN => n8930);
   REGISTERS_reg_4_26_inst : DFF_X1 port map( D => n2501, CK => CLK, Q => 
                           n_1053, QN => n8931);
   REGISTERS_reg_4_25_inst : DFF_X1 port map( D => n2500, CK => CLK, Q => 
                           n_1054, QN => n8932);
   REGISTERS_reg_4_24_inst : DFF_X1 port map( D => n2499, CK => CLK, Q => 
                           n_1055, QN => n8933);
   REGISTERS_reg_3_31_inst : DFF_X1 port map( D => n2538, CK => CLK, Q => 
                           n_1056, QN => n8894);
   REGISTERS_reg_3_30_inst : DFF_X1 port map( D => n2537, CK => CLK, Q => 
                           n_1057, QN => n8895);
   REGISTERS_reg_3_29_inst : DFF_X1 port map( D => n2536, CK => CLK, Q => 
                           n_1058, QN => n8896);
   REGISTERS_reg_3_28_inst : DFF_X1 port map( D => n2535, CK => CLK, Q => 
                           n_1059, QN => n8897);
   REGISTERS_reg_3_27_inst : DFF_X1 port map( D => n2534, CK => CLK, Q => 
                           n_1060, QN => n8898);
   REGISTERS_reg_3_26_inst : DFF_X1 port map( D => n2533, CK => CLK, Q => 
                           n_1061, QN => n8899);
   REGISTERS_reg_3_25_inst : DFF_X1 port map( D => n2532, CK => CLK, Q => 
                           n_1062, QN => n8900);
   REGISTERS_reg_3_24_inst : DFF_X1 port map( D => n2531, CK => CLK, Q => 
                           n_1063, QN => n8901);
   REGISTERS_reg_12_31_inst : DFF_X1 port map( D => n2250, CK => CLK, Q => 
                           n_1064, QN => n9182);
   REGISTERS_reg_12_30_inst : DFF_X1 port map( D => n2249, CK => CLK, Q => 
                           n_1065, QN => n9183);
   REGISTERS_reg_12_29_inst : DFF_X1 port map( D => n2248, CK => CLK, Q => 
                           n_1066, QN => n9184);
   REGISTERS_reg_12_28_inst : DFF_X1 port map( D => n2247, CK => CLK, Q => 
                           n_1067, QN => n9185);
   REGISTERS_reg_12_27_inst : DFF_X1 port map( D => n2246, CK => CLK, Q => 
                           n_1068, QN => n9186);
   REGISTERS_reg_12_26_inst : DFF_X1 port map( D => n2245, CK => CLK, Q => 
                           n_1069, QN => n9187);
   REGISTERS_reg_12_25_inst : DFF_X1 port map( D => n2244, CK => CLK, Q => 
                           n_1070, QN => n9188);
   REGISTERS_reg_12_24_inst : DFF_X1 port map( D => n2243, CK => CLK, Q => 
                           n_1071, QN => n9189);
   REGISTERS_reg_11_31_inst : DFF_X1 port map( D => n2282, CK => CLK, Q => 
                           n_1072, QN => n9150);
   REGISTERS_reg_11_30_inst : DFF_X1 port map( D => n2281, CK => CLK, Q => 
                           n_1073, QN => n9151);
   REGISTERS_reg_11_29_inst : DFF_X1 port map( D => n2280, CK => CLK, Q => 
                           n_1074, QN => n9152);
   REGISTERS_reg_11_28_inst : DFF_X1 port map( D => n2279, CK => CLK, Q => 
                           n_1075, QN => n9153);
   REGISTERS_reg_11_27_inst : DFF_X1 port map( D => n2278, CK => CLK, Q => 
                           n_1076, QN => n9154);
   REGISTERS_reg_11_26_inst : DFF_X1 port map( D => n2277, CK => CLK, Q => 
                           n_1077, QN => n9155);
   REGISTERS_reg_11_25_inst : DFF_X1 port map( D => n2276, CK => CLK, Q => 
                           n_1078, QN => n9156);
   REGISTERS_reg_11_24_inst : DFF_X1 port map( D => n2275, CK => CLK, Q => 
                           n_1079, QN => n9157);
   REGISTERS_reg_2_31_inst : DFF_X1 port map( D => n2570, CK => CLK, Q => 
                           n_1080, QN => n8862);
   REGISTERS_reg_2_30_inst : DFF_X1 port map( D => n2569, CK => CLK, Q => 
                           n_1081, QN => n8863);
   REGISTERS_reg_2_29_inst : DFF_X1 port map( D => n2568, CK => CLK, Q => 
                           n_1082, QN => n8864);
   REGISTERS_reg_2_28_inst : DFF_X1 port map( D => n2567, CK => CLK, Q => 
                           n_1083, QN => n8865);
   REGISTERS_reg_2_27_inst : DFF_X1 port map( D => n2566, CK => CLK, Q => 
                           n_1084, QN => n8866);
   REGISTERS_reg_2_26_inst : DFF_X1 port map( D => n2565, CK => CLK, Q => 
                           n_1085, QN => n8867);
   REGISTERS_reg_2_25_inst : DFF_X1 port map( D => n2564, CK => CLK, Q => 
                           n_1086, QN => n8868);
   REGISTERS_reg_2_24_inst : DFF_X1 port map( D => n2563, CK => CLK, Q => 
                           n_1087, QN => n8869);
   REGISTERS_reg_1_31_inst : DFF_X1 port map( D => n2602, CK => CLK, Q => 
                           n_1088, QN => n8830);
   REGISTERS_reg_1_30_inst : DFF_X1 port map( D => n2601, CK => CLK, Q => 
                           n_1089, QN => n8831);
   REGISTERS_reg_1_29_inst : DFF_X1 port map( D => n2600, CK => CLK, Q => 
                           n_1090, QN => n8832);
   REGISTERS_reg_1_28_inst : DFF_X1 port map( D => n2599, CK => CLK, Q => 
                           n_1091, QN => n8833);
   REGISTERS_reg_1_27_inst : DFF_X1 port map( D => n2598, CK => CLK, Q => 
                           n_1092, QN => n8834);
   REGISTERS_reg_1_26_inst : DFF_X1 port map( D => n2597, CK => CLK, Q => 
                           n_1093, QN => n8835);
   REGISTERS_reg_1_25_inst : DFF_X1 port map( D => n2596, CK => CLK, Q => 
                           n_1094, QN => n8836);
   REGISTERS_reg_1_24_inst : DFF_X1 port map( D => n2595, CK => CLK, Q => 
                           n_1095, QN => n8837);
   REGISTERS_reg_20_23_inst : DFF_X1 port map( D => n1986, CK => CLK, Q => 
                           n_1096, QN => n9446);
   REGISTERS_reg_20_22_inst : DFF_X1 port map( D => n1985, CK => CLK, Q => 
                           n_1097, QN => n9447);
   REGISTERS_reg_20_21_inst : DFF_X1 port map( D => n1984, CK => CLK, Q => 
                           n_1098, QN => n9448);
   REGISTERS_reg_20_20_inst : DFF_X1 port map( D => n1983, CK => CLK, Q => 
                           n_1099, QN => n9449);
   REGISTERS_reg_20_19_inst : DFF_X1 port map( D => n1982, CK => CLK, Q => 
                           n_1100, QN => n9450);
   REGISTERS_reg_20_18_inst : DFF_X1 port map( D => n1981, CK => CLK, Q => 
                           n_1101, QN => n9451);
   REGISTERS_reg_20_17_inst : DFF_X1 port map( D => n1980, CK => CLK, Q => 
                           n_1102, QN => n9452);
   REGISTERS_reg_20_16_inst : DFF_X1 port map( D => n1979, CK => CLK, Q => 
                           n_1103, QN => n9453);
   REGISTERS_reg_20_15_inst : DFF_X1 port map( D => n1978, CK => CLK, Q => 
                           n_1104, QN => n9454);
   REGISTERS_reg_20_14_inst : DFF_X1 port map( D => n1977, CK => CLK, Q => 
                           n_1105, QN => n9455);
   REGISTERS_reg_20_13_inst : DFF_X1 port map( D => n1976, CK => CLK, Q => 
                           n_1106, QN => n9456);
   REGISTERS_reg_20_12_inst : DFF_X1 port map( D => n1975, CK => CLK, Q => 
                           n_1107, QN => n9457);
   REGISTERS_reg_20_11_inst : DFF_X1 port map( D => n1974, CK => CLK, Q => 
                           n_1108, QN => n9458);
   REGISTERS_reg_20_10_inst : DFF_X1 port map( D => n1973, CK => CLK, Q => 
                           n_1109, QN => n9459);
   REGISTERS_reg_20_9_inst : DFF_X1 port map( D => n1972, CK => CLK, Q => 
                           n_1110, QN => n9460);
   REGISTERS_reg_20_8_inst : DFF_X1 port map( D => n1971, CK => CLK, Q => 
                           n_1111, QN => n9461);
   REGISTERS_reg_20_7_inst : DFF_X1 port map( D => n1970, CK => CLK, Q => 
                           n_1112, QN => n9462);
   REGISTERS_reg_20_6_inst : DFF_X1 port map( D => n1969, CK => CLK, Q => 
                           n_1113, QN => n9463);
   REGISTERS_reg_20_5_inst : DFF_X1 port map( D => n1968, CK => CLK, Q => 
                           n_1114, QN => n9464);
   REGISTERS_reg_20_4_inst : DFF_X1 port map( D => n1967, CK => CLK, Q => 
                           n_1115, QN => n9465);
   REGISTERS_reg_20_3_inst : DFF_X1 port map( D => n1966, CK => CLK, Q => 
                           n_1116, QN => n9466);
   REGISTERS_reg_20_2_inst : DFF_X1 port map( D => n1965, CK => CLK, Q => 
                           n_1117, QN => n9467);
   REGISTERS_reg_20_1_inst : DFF_X1 port map( D => n1964, CK => CLK, Q => 
                           n_1118, QN => n9468);
   REGISTERS_reg_20_0_inst : DFF_X1 port map( D => n1963, CK => CLK, Q => 
                           n_1119, QN => n9469);
   REGISTERS_reg_16_31_inst : DFF_X1 port map( D => n2122, CK => CLK, Q => 
                           n_1120, QN => n9310);
   REGISTERS_reg_16_30_inst : DFF_X1 port map( D => n2121, CK => CLK, Q => 
                           n_1121, QN => n9311);
   REGISTERS_reg_16_29_inst : DFF_X1 port map( D => n2120, CK => CLK, Q => 
                           n_1122, QN => n9312);
   REGISTERS_reg_16_28_inst : DFF_X1 port map( D => n2119, CK => CLK, Q => 
                           n_1123, QN => n9313);
   REGISTERS_reg_16_27_inst : DFF_X1 port map( D => n2118, CK => CLK, Q => 
                           n_1124, QN => n9314);
   REGISTERS_reg_16_26_inst : DFF_X1 port map( D => n2117, CK => CLK, Q => 
                           n_1125, QN => n9315);
   REGISTERS_reg_16_25_inst : DFF_X1 port map( D => n2116, CK => CLK, Q => 
                           n_1126, QN => n9316);
   REGISTERS_reg_16_24_inst : DFF_X1 port map( D => n2115, CK => CLK, Q => 
                           n_1127, QN => n9317);
   REGISTERS_reg_22_31_inst : DFF_X1 port map( D => n1930, CK => CLK, Q => 
                           n_1128, QN => n9502);
   REGISTERS_reg_22_30_inst : DFF_X1 port map( D => n1929, CK => CLK, Q => 
                           n_1129, QN => n9503);
   REGISTERS_reg_22_29_inst : DFF_X1 port map( D => n1928, CK => CLK, Q => 
                           n_1130, QN => n9504);
   REGISTERS_reg_22_28_inst : DFF_X1 port map( D => n1927, CK => CLK, Q => 
                           n_1131, QN => n9505);
   REGISTERS_reg_22_27_inst : DFF_X1 port map( D => n1926, CK => CLK, Q => 
                           n_1132, QN => n9506);
   REGISTERS_reg_22_26_inst : DFF_X1 port map( D => n1925, CK => CLK, Q => 
                           n_1133, QN => n9507);
   REGISTERS_reg_22_25_inst : DFF_X1 port map( D => n1924, CK => CLK, Q => 
                           n_1134, QN => n9508);
   REGISTERS_reg_22_24_inst : DFF_X1 port map( D => n1923, CK => CLK, Q => 
                           n_1135, QN => n9509);
   REGISTERS_reg_29_31_inst : DFF_X1 port map( D => n1706, CK => CLK, Q => 
                           n_1136, QN => n9726);
   REGISTERS_reg_29_30_inst : DFF_X1 port map( D => n1705, CK => CLK, Q => 
                           n_1137, QN => n9727);
   REGISTERS_reg_29_29_inst : DFF_X1 port map( D => n1704, CK => CLK, Q => 
                           n_1138, QN => n9728);
   REGISTERS_reg_29_28_inst : DFF_X1 port map( D => n1703, CK => CLK, Q => 
                           n_1139, QN => n9729);
   REGISTERS_reg_29_27_inst : DFF_X1 port map( D => n1702, CK => CLK, Q => 
                           n_1140, QN => n9730);
   REGISTERS_reg_29_26_inst : DFF_X1 port map( D => n1701, CK => CLK, Q => 
                           n_1141, QN => n9731);
   REGISTERS_reg_29_25_inst : DFF_X1 port map( D => n1700, CK => CLK, Q => 
                           n_1142, QN => n9732);
   REGISTERS_reg_29_24_inst : DFF_X1 port map( D => n1699, CK => CLK, Q => 
                           n_1143, QN => n9733);
   REGISTERS_reg_26_31_inst : DFF_X1 port map( D => n1802, CK => CLK, Q => 
                           n_1144, QN => n9630);
   REGISTERS_reg_26_30_inst : DFF_X1 port map( D => n1801, CK => CLK, Q => 
                           n_1145, QN => n9631);
   REGISTERS_reg_26_29_inst : DFF_X1 port map( D => n1800, CK => CLK, Q => 
                           n_1146, QN => n9632);
   REGISTERS_reg_26_28_inst : DFF_X1 port map( D => n1799, CK => CLK, Q => 
                           n_1147, QN => n9633);
   REGISTERS_reg_26_27_inst : DFF_X1 port map( D => n1798, CK => CLK, Q => 
                           n_1148, QN => n9634);
   REGISTERS_reg_26_26_inst : DFF_X1 port map( D => n1797, CK => CLK, Q => 
                           n_1149, QN => n9635);
   REGISTERS_reg_26_25_inst : DFF_X1 port map( D => n1796, CK => CLK, Q => 
                           n_1150, QN => n9636);
   REGISTERS_reg_26_24_inst : DFF_X1 port map( D => n1795, CK => CLK, Q => 
                           n_1151, QN => n9637);
   REGISTERS_reg_28_23_inst : DFF_X1 port map( D => n1730, CK => CLK, Q => 
                           n_1152, QN => n9702);
   REGISTERS_reg_28_22_inst : DFF_X1 port map( D => n1729, CK => CLK, Q => 
                           n_1153, QN => n9703);
   REGISTERS_reg_28_21_inst : DFF_X1 port map( D => n1728, CK => CLK, Q => 
                           n_1154, QN => n9704);
   REGISTERS_reg_28_20_inst : DFF_X1 port map( D => n1727, CK => CLK, Q => 
                           n_1155, QN => n9705);
   REGISTERS_reg_28_19_inst : DFF_X1 port map( D => n1726, CK => CLK, Q => 
                           n_1156, QN => n9706);
   REGISTERS_reg_28_18_inst : DFF_X1 port map( D => n1725, CK => CLK, Q => 
                           n_1157, QN => n9707);
   REGISTERS_reg_28_17_inst : DFF_X1 port map( D => n1724, CK => CLK, Q => 
                           n_1158, QN => n9708);
   REGISTERS_reg_28_16_inst : DFF_X1 port map( D => n1723, CK => CLK, Q => 
                           n_1159, QN => n9709);
   REGISTERS_reg_28_15_inst : DFF_X1 port map( D => n1722, CK => CLK, Q => 
                           n_1160, QN => n9710);
   REGISTERS_reg_28_14_inst : DFF_X1 port map( D => n1721, CK => CLK, Q => 
                           n_1161, QN => n9711);
   REGISTERS_reg_28_13_inst : DFF_X1 port map( D => n1720, CK => CLK, Q => 
                           n_1162, QN => n9712);
   REGISTERS_reg_28_12_inst : DFF_X1 port map( D => n1719, CK => CLK, Q => 
                           n_1163, QN => n9713);
   REGISTERS_reg_28_11_inst : DFF_X1 port map( D => n1718, CK => CLK, Q => 
                           n_1164, QN => n9714);
   REGISTERS_reg_28_10_inst : DFF_X1 port map( D => n1717, CK => CLK, Q => 
                           n_1165, QN => n9715);
   REGISTERS_reg_28_9_inst : DFF_X1 port map( D => n1716, CK => CLK, Q => 
                           n_1166, QN => n9716);
   REGISTERS_reg_28_8_inst : DFF_X1 port map( D => n1715, CK => CLK, Q => 
                           n_1167, QN => n9717);
   REGISTERS_reg_28_7_inst : DFF_X1 port map( D => n1714, CK => CLK, Q => 
                           n_1168, QN => n9718);
   REGISTERS_reg_28_6_inst : DFF_X1 port map( D => n1713, CK => CLK, Q => 
                           n_1169, QN => n9719);
   REGISTERS_reg_28_5_inst : DFF_X1 port map( D => n1712, CK => CLK, Q => 
                           n_1170, QN => n9720);
   REGISTERS_reg_28_4_inst : DFF_X1 port map( D => n1711, CK => CLK, Q => 
                           n_1171, QN => n9721);
   REGISTERS_reg_28_3_inst : DFF_X1 port map( D => n1710, CK => CLK, Q => 
                           n_1172, QN => n9722);
   REGISTERS_reg_28_2_inst : DFF_X1 port map( D => n1709, CK => CLK, Q => 
                           n_1173, QN => n9723);
   REGISTERS_reg_28_1_inst : DFF_X1 port map( D => n1708, CK => CLK, Q => 
                           n_1174, QN => n9724);
   REGISTERS_reg_28_0_inst : DFF_X1 port map( D => n1707, CK => CLK, Q => 
                           n_1175, QN => n9725);
   REGISTERS_reg_24_23_inst : DFF_X1 port map( D => n1858, CK => CLK, Q => 
                           n_1176, QN => n9574);
   REGISTERS_reg_24_22_inst : DFF_X1 port map( D => n1857, CK => CLK, Q => 
                           n_1177, QN => n9575);
   REGISTERS_reg_24_21_inst : DFF_X1 port map( D => n1856, CK => CLK, Q => 
                           n_1178, QN => n9576);
   REGISTERS_reg_24_20_inst : DFF_X1 port map( D => n1855, CK => CLK, Q => 
                           n_1179, QN => n9577);
   REGISTERS_reg_24_19_inst : DFF_X1 port map( D => n1854, CK => CLK, Q => 
                           n_1180, QN => n9578);
   REGISTERS_reg_24_18_inst : DFF_X1 port map( D => n1853, CK => CLK, Q => 
                           n_1181, QN => n9579);
   REGISTERS_reg_24_17_inst : DFF_X1 port map( D => n1852, CK => CLK, Q => 
                           n_1182, QN => n9580);
   REGISTERS_reg_24_16_inst : DFF_X1 port map( D => n1851, CK => CLK, Q => 
                           n_1183, QN => n9581);
   REGISTERS_reg_24_15_inst : DFF_X1 port map( D => n1850, CK => CLK, Q => 
                           n_1184, QN => n9582);
   REGISTERS_reg_24_14_inst : DFF_X1 port map( D => n1849, CK => CLK, Q => 
                           n_1185, QN => n9583);
   REGISTERS_reg_24_13_inst : DFF_X1 port map( D => n1848, CK => CLK, Q => 
                           n_1186, QN => n9584);
   REGISTERS_reg_24_12_inst : DFF_X1 port map( D => n1847, CK => CLK, Q => 
                           n_1187, QN => n9585);
   REGISTERS_reg_24_11_inst : DFF_X1 port map( D => n1846, CK => CLK, Q => 
                           n_1188, QN => n9586);
   REGISTERS_reg_24_10_inst : DFF_X1 port map( D => n1845, CK => CLK, Q => 
                           n_1189, QN => n9587);
   REGISTERS_reg_24_9_inst : DFF_X1 port map( D => n1844, CK => CLK, Q => 
                           n_1190, QN => n9588);
   REGISTERS_reg_24_8_inst : DFF_X1 port map( D => n1843, CK => CLK, Q => 
                           n_1191, QN => n9589);
   REGISTERS_reg_24_7_inst : DFF_X1 port map( D => n1842, CK => CLK, Q => 
                           n_1192, QN => n9590);
   REGISTERS_reg_24_6_inst : DFF_X1 port map( D => n1841, CK => CLK, Q => 
                           n_1193, QN => n9591);
   REGISTERS_reg_24_5_inst : DFF_X1 port map( D => n1840, CK => CLK, Q => 
                           n_1194, QN => n9592);
   REGISTERS_reg_24_4_inst : DFF_X1 port map( D => n1839, CK => CLK, Q => 
                           n_1195, QN => n9593);
   REGISTERS_reg_24_3_inst : DFF_X1 port map( D => n1838, CK => CLK, Q => 
                           n_1196, QN => n9594);
   REGISTERS_reg_24_2_inst : DFF_X1 port map( D => n1837, CK => CLK, Q => 
                           n_1197, QN => n9595);
   REGISTERS_reg_24_1_inst : DFF_X1 port map( D => n1836, CK => CLK, Q => 
                           n_1198, QN => n9596);
   REGISTERS_reg_24_0_inst : DFF_X1 port map( D => n1835, CK => CLK, Q => 
                           n_1199, QN => n9597);
   REGISTERS_reg_18_23_inst : DFF_X1 port map( D => n2050, CK => CLK, Q => 
                           n_1200, QN => n9382);
   REGISTERS_reg_18_22_inst : DFF_X1 port map( D => n2049, CK => CLK, Q => 
                           n_1201, QN => n9383);
   REGISTERS_reg_18_21_inst : DFF_X1 port map( D => n2048, CK => CLK, Q => 
                           n_1202, QN => n9384);
   REGISTERS_reg_18_20_inst : DFF_X1 port map( D => n2047, CK => CLK, Q => 
                           n_1203, QN => n9385);
   REGISTERS_reg_18_19_inst : DFF_X1 port map( D => n2046, CK => CLK, Q => 
                           n_1204, QN => n9386);
   REGISTERS_reg_18_18_inst : DFF_X1 port map( D => n2045, CK => CLK, Q => 
                           n_1205, QN => n9387);
   REGISTERS_reg_18_17_inst : DFF_X1 port map( D => n2044, CK => CLK, Q => 
                           n_1206, QN => n9388);
   REGISTERS_reg_18_16_inst : DFF_X1 port map( D => n2043, CK => CLK, Q => 
                           n_1207, QN => n9389);
   REGISTERS_reg_18_15_inst : DFF_X1 port map( D => n2042, CK => CLK, Q => 
                           n_1208, QN => n9390);
   REGISTERS_reg_18_14_inst : DFF_X1 port map( D => n2041, CK => CLK, Q => 
                           n_1209, QN => n9391);
   REGISTERS_reg_18_13_inst : DFF_X1 port map( D => n2040, CK => CLK, Q => 
                           n_1210, QN => n9392);
   REGISTERS_reg_18_12_inst : DFF_X1 port map( D => n2039, CK => CLK, Q => 
                           n_1211, QN => n9393);
   REGISTERS_reg_18_11_inst : DFF_X1 port map( D => n2038, CK => CLK, Q => 
                           n_1212, QN => n9394);
   REGISTERS_reg_18_10_inst : DFF_X1 port map( D => n2037, CK => CLK, Q => 
                           n_1213, QN => n9395);
   REGISTERS_reg_18_9_inst : DFF_X1 port map( D => n2036, CK => CLK, Q => 
                           n_1214, QN => n9396);
   REGISTERS_reg_18_8_inst : DFF_X1 port map( D => n2035, CK => CLK, Q => 
                           n_1215, QN => n9397);
   REGISTERS_reg_18_7_inst : DFF_X1 port map( D => n2034, CK => CLK, Q => 
                           n_1216, QN => n9398);
   REGISTERS_reg_18_6_inst : DFF_X1 port map( D => n2033, CK => CLK, Q => 
                           n_1217, QN => n9399);
   REGISTERS_reg_18_5_inst : DFF_X1 port map( D => n2032, CK => CLK, Q => 
                           n_1218, QN => n9400);
   REGISTERS_reg_18_4_inst : DFF_X1 port map( D => n2031, CK => CLK, Q => 
                           n_1219, QN => n9401);
   REGISTERS_reg_18_3_inst : DFF_X1 port map( D => n2030, CK => CLK, Q => 
                           n_1220, QN => n9402);
   REGISTERS_reg_18_2_inst : DFF_X1 port map( D => n2029, CK => CLK, Q => 
                           n_1221, QN => n9403);
   REGISTERS_reg_18_1_inst : DFF_X1 port map( D => n2028, CK => CLK, Q => 
                           n_1222, QN => n9404);
   REGISTERS_reg_18_0_inst : DFF_X1 port map( D => n2027, CK => CLK, Q => 
                           n_1223, QN => n9405);
   REGISTERS_reg_15_23_inst : DFF_X1 port map( D => n2146, CK => CLK, Q => 
                           n_1224, QN => n9286);
   REGISTERS_reg_15_22_inst : DFF_X1 port map( D => n2145, CK => CLK, Q => 
                           n_1225, QN => n9287);
   REGISTERS_reg_15_21_inst : DFF_X1 port map( D => n2144, CK => CLK, Q => 
                           n_1226, QN => n9288);
   REGISTERS_reg_15_20_inst : DFF_X1 port map( D => n2143, CK => CLK, Q => 
                           n_1227, QN => n9289);
   REGISTERS_reg_15_19_inst : DFF_X1 port map( D => n2142, CK => CLK, Q => 
                           n_1228, QN => n9290);
   REGISTERS_reg_15_18_inst : DFF_X1 port map( D => n2141, CK => CLK, Q => 
                           n_1229, QN => n9291);
   REGISTERS_reg_15_17_inst : DFF_X1 port map( D => n2140, CK => CLK, Q => 
                           n_1230, QN => n9292);
   REGISTERS_reg_15_16_inst : DFF_X1 port map( D => n2139, CK => CLK, Q => 
                           n_1231, QN => n9293);
   REGISTERS_reg_15_15_inst : DFF_X1 port map( D => n2138, CK => CLK, Q => 
                           n_1232, QN => n9294);
   REGISTERS_reg_15_14_inst : DFF_X1 port map( D => n2137, CK => CLK, Q => 
                           n_1233, QN => n9295);
   REGISTERS_reg_15_13_inst : DFF_X1 port map( D => n2136, CK => CLK, Q => 
                           n_1234, QN => n9296);
   REGISTERS_reg_15_12_inst : DFF_X1 port map( D => n2135, CK => CLK, Q => 
                           n_1235, QN => n9297);
   REGISTERS_reg_15_11_inst : DFF_X1 port map( D => n2134, CK => CLK, Q => 
                           n_1236, QN => n9298);
   REGISTERS_reg_15_10_inst : DFF_X1 port map( D => n2133, CK => CLK, Q => 
                           n_1237, QN => n9299);
   REGISTERS_reg_15_9_inst : DFF_X1 port map( D => n2132, CK => CLK, Q => 
                           n_1238, QN => n9300);
   REGISTERS_reg_15_8_inst : DFF_X1 port map( D => n2131, CK => CLK, Q => 
                           n_1239, QN => n9301);
   REGISTERS_reg_15_7_inst : DFF_X1 port map( D => n2130, CK => CLK, Q => 
                           n_1240, QN => n9302);
   REGISTERS_reg_15_6_inst : DFF_X1 port map( D => n2129, CK => CLK, Q => 
                           n_1241, QN => n9303);
   REGISTERS_reg_15_5_inst : DFF_X1 port map( D => n2128, CK => CLK, Q => 
                           n_1242, QN => n9304);
   REGISTERS_reg_15_4_inst : DFF_X1 port map( D => n2127, CK => CLK, Q => 
                           n_1243, QN => n9305);
   REGISTERS_reg_15_3_inst : DFF_X1 port map( D => n2126, CK => CLK, Q => 
                           n_1244, QN => n9306);
   REGISTERS_reg_15_2_inst : DFF_X1 port map( D => n2125, CK => CLK, Q => 
                           n_1245, QN => n9307);
   REGISTERS_reg_15_1_inst : DFF_X1 port map( D => n2124, CK => CLK, Q => 
                           n_1246, QN => n9308);
   REGISTERS_reg_15_0_inst : DFF_X1 port map( D => n2123, CK => CLK, Q => 
                           n_1247, QN => n9309);
   REGISTERS_reg_8_23_inst : DFF_X1 port map( D => n2370, CK => CLK, Q => 
                           n_1248, QN => n9062);
   REGISTERS_reg_8_22_inst : DFF_X1 port map( D => n2369, CK => CLK, Q => 
                           n_1249, QN => n9063);
   REGISTERS_reg_8_21_inst : DFF_X1 port map( D => n2368, CK => CLK, Q => 
                           n_1250, QN => n9064);
   REGISTERS_reg_8_20_inst : DFF_X1 port map( D => n2367, CK => CLK, Q => 
                           n_1251, QN => n9065);
   REGISTERS_reg_8_19_inst : DFF_X1 port map( D => n2366, CK => CLK, Q => 
                           n_1252, QN => n9066);
   REGISTERS_reg_8_18_inst : DFF_X1 port map( D => n2365, CK => CLK, Q => 
                           n_1253, QN => n9067);
   REGISTERS_reg_8_17_inst : DFF_X1 port map( D => n2364, CK => CLK, Q => 
                           n_1254, QN => n9068);
   REGISTERS_reg_8_16_inst : DFF_X1 port map( D => n2363, CK => CLK, Q => 
                           n_1255, QN => n9069);
   REGISTERS_reg_8_15_inst : DFF_X1 port map( D => n2362, CK => CLK, Q => 
                           n_1256, QN => n9070);
   REGISTERS_reg_8_14_inst : DFF_X1 port map( D => n2361, CK => CLK, Q => 
                           n_1257, QN => n9071);
   REGISTERS_reg_8_13_inst : DFF_X1 port map( D => n2360, CK => CLK, Q => 
                           n_1258, QN => n9072);
   REGISTERS_reg_8_12_inst : DFF_X1 port map( D => n2359, CK => CLK, Q => 
                           n_1259, QN => n9073);
   REGISTERS_reg_8_11_inst : DFF_X1 port map( D => n2358, CK => CLK, Q => 
                           n_1260, QN => n9074);
   REGISTERS_reg_8_10_inst : DFF_X1 port map( D => n2357, CK => CLK, Q => 
                           n_1261, QN => n9075);
   REGISTERS_reg_8_9_inst : DFF_X1 port map( D => n2356, CK => CLK, Q => n_1262
                           , QN => n9076);
   REGISTERS_reg_8_8_inst : DFF_X1 port map( D => n2355, CK => CLK, Q => n_1263
                           , QN => n9077);
   REGISTERS_reg_8_7_inst : DFF_X1 port map( D => n2354, CK => CLK, Q => n_1264
                           , QN => n9078);
   REGISTERS_reg_8_6_inst : DFF_X1 port map( D => n2353, CK => CLK, Q => n_1265
                           , QN => n9079);
   REGISTERS_reg_8_5_inst : DFF_X1 port map( D => n2352, CK => CLK, Q => n_1266
                           , QN => n9080);
   REGISTERS_reg_8_4_inst : DFF_X1 port map( D => n2351, CK => CLK, Q => n_1267
                           , QN => n9081);
   REGISTERS_reg_8_3_inst : DFF_X1 port map( D => n2350, CK => CLK, Q => n_1268
                           , QN => n9082);
   REGISTERS_reg_8_2_inst : DFF_X1 port map( D => n2349, CK => CLK, Q => n_1269
                           , QN => n9083);
   REGISTERS_reg_8_1_inst : DFF_X1 port map( D => n2348, CK => CLK, Q => n_1270
                           , QN => n9084);
   REGISTERS_reg_8_0_inst : DFF_X1 port map( D => n2347, CK => CLK, Q => n_1271
                           , QN => n9085);
   REGISTERS_reg_4_23_inst : DFF_X1 port map( D => n2498, CK => CLK, Q => 
                           n_1272, QN => n8934);
   REGISTERS_reg_4_22_inst : DFF_X1 port map( D => n2497, CK => CLK, Q => 
                           n_1273, QN => n8935);
   REGISTERS_reg_4_21_inst : DFF_X1 port map( D => n2496, CK => CLK, Q => 
                           n_1274, QN => n8936);
   REGISTERS_reg_4_20_inst : DFF_X1 port map( D => n2495, CK => CLK, Q => 
                           n_1275, QN => n8937);
   REGISTERS_reg_4_19_inst : DFF_X1 port map( D => n2494, CK => CLK, Q => 
                           n_1276, QN => n8938);
   REGISTERS_reg_4_18_inst : DFF_X1 port map( D => n2493, CK => CLK, Q => 
                           n_1277, QN => n8939);
   REGISTERS_reg_4_17_inst : DFF_X1 port map( D => n2492, CK => CLK, Q => 
                           n_1278, QN => n8940);
   REGISTERS_reg_4_16_inst : DFF_X1 port map( D => n2491, CK => CLK, Q => 
                           n_1279, QN => n8941);
   REGISTERS_reg_4_15_inst : DFF_X1 port map( D => n2490, CK => CLK, Q => 
                           n_1280, QN => n8942);
   REGISTERS_reg_4_14_inst : DFF_X1 port map( D => n2489, CK => CLK, Q => 
                           n_1281, QN => n8943);
   REGISTERS_reg_4_13_inst : DFF_X1 port map( D => n2488, CK => CLK, Q => 
                           n_1282, QN => n8944);
   REGISTERS_reg_4_12_inst : DFF_X1 port map( D => n2487, CK => CLK, Q => 
                           n_1283, QN => n8945);
   REGISTERS_reg_4_11_inst : DFF_X1 port map( D => n2486, CK => CLK, Q => 
                           n_1284, QN => n8946);
   REGISTERS_reg_4_10_inst : DFF_X1 port map( D => n2485, CK => CLK, Q => 
                           n_1285, QN => n8947);
   REGISTERS_reg_4_9_inst : DFF_X1 port map( D => n2484, CK => CLK, Q => n_1286
                           , QN => n8948);
   REGISTERS_reg_4_8_inst : DFF_X1 port map( D => n2483, CK => CLK, Q => n_1287
                           , QN => n8949);
   REGISTERS_reg_4_7_inst : DFF_X1 port map( D => n2482, CK => CLK, Q => n_1288
                           , QN => n8950);
   REGISTERS_reg_4_6_inst : DFF_X1 port map( D => n2481, CK => CLK, Q => n_1289
                           , QN => n8951);
   REGISTERS_reg_4_5_inst : DFF_X1 port map( D => n2480, CK => CLK, Q => n_1290
                           , QN => n8952);
   REGISTERS_reg_4_4_inst : DFF_X1 port map( D => n2479, CK => CLK, Q => n_1291
                           , QN => n8953);
   REGISTERS_reg_4_3_inst : DFF_X1 port map( D => n2478, CK => CLK, Q => n_1292
                           , QN => n8954);
   REGISTERS_reg_4_2_inst : DFF_X1 port map( D => n2477, CK => CLK, Q => n_1293
                           , QN => n8955);
   REGISTERS_reg_4_1_inst : DFF_X1 port map( D => n2476, CK => CLK, Q => n_1294
                           , QN => n8956);
   REGISTERS_reg_4_0_inst : DFF_X1 port map( D => n2475, CK => CLK, Q => n_1295
                           , QN => n8957);
   REGISTERS_reg_3_23_inst : DFF_X1 port map( D => n2530, CK => CLK, Q => 
                           n_1296, QN => n8902);
   REGISTERS_reg_3_22_inst : DFF_X1 port map( D => n2529, CK => CLK, Q => 
                           n_1297, QN => n8903);
   REGISTERS_reg_3_21_inst : DFF_X1 port map( D => n2528, CK => CLK, Q => 
                           n_1298, QN => n8904);
   REGISTERS_reg_3_20_inst : DFF_X1 port map( D => n2527, CK => CLK, Q => 
                           n_1299, QN => n8905);
   REGISTERS_reg_3_19_inst : DFF_X1 port map( D => n2526, CK => CLK, Q => 
                           n_1300, QN => n8906);
   REGISTERS_reg_3_18_inst : DFF_X1 port map( D => n2525, CK => CLK, Q => 
                           n_1301, QN => n8907);
   REGISTERS_reg_3_17_inst : DFF_X1 port map( D => n2524, CK => CLK, Q => 
                           n_1302, QN => n8908);
   REGISTERS_reg_3_16_inst : DFF_X1 port map( D => n2523, CK => CLK, Q => 
                           n_1303, QN => n8909);
   REGISTERS_reg_3_15_inst : DFF_X1 port map( D => n2522, CK => CLK, Q => 
                           n_1304, QN => n8910);
   REGISTERS_reg_3_14_inst : DFF_X1 port map( D => n2521, CK => CLK, Q => 
                           n_1305, QN => n8911);
   REGISTERS_reg_3_13_inst : DFF_X1 port map( D => n2520, CK => CLK, Q => 
                           n_1306, QN => n8912);
   REGISTERS_reg_3_12_inst : DFF_X1 port map( D => n2519, CK => CLK, Q => 
                           n_1307, QN => n8913);
   REGISTERS_reg_3_11_inst : DFF_X1 port map( D => n2518, CK => CLK, Q => 
                           n_1308, QN => n8914);
   REGISTERS_reg_3_10_inst : DFF_X1 port map( D => n2517, CK => CLK, Q => 
                           n_1309, QN => n8915);
   REGISTERS_reg_3_9_inst : DFF_X1 port map( D => n2516, CK => CLK, Q => n_1310
                           , QN => n8916);
   REGISTERS_reg_3_8_inst : DFF_X1 port map( D => n2515, CK => CLK, Q => n_1311
                           , QN => n8917);
   REGISTERS_reg_3_7_inst : DFF_X1 port map( D => n2514, CK => CLK, Q => n_1312
                           , QN => n8918);
   REGISTERS_reg_3_6_inst : DFF_X1 port map( D => n2513, CK => CLK, Q => n_1313
                           , QN => n8919);
   REGISTERS_reg_3_5_inst : DFF_X1 port map( D => n2512, CK => CLK, Q => n_1314
                           , QN => n8920);
   REGISTERS_reg_3_4_inst : DFF_X1 port map( D => n2511, CK => CLK, Q => n_1315
                           , QN => n8921);
   REGISTERS_reg_3_3_inst : DFF_X1 port map( D => n2510, CK => CLK, Q => n_1316
                           , QN => n8922);
   REGISTERS_reg_3_2_inst : DFF_X1 port map( D => n2509, CK => CLK, Q => n_1317
                           , QN => n8923);
   REGISTERS_reg_3_1_inst : DFF_X1 port map( D => n2508, CK => CLK, Q => n_1318
                           , QN => n8924);
   REGISTERS_reg_3_0_inst : DFF_X1 port map( D => n2507, CK => CLK, Q => n_1319
                           , QN => n8925);
   REGISTERS_reg_12_23_inst : DFF_X1 port map( D => n2242, CK => CLK, Q => 
                           n_1320, QN => n9190);
   REGISTERS_reg_12_22_inst : DFF_X1 port map( D => n2241, CK => CLK, Q => 
                           n_1321, QN => n9191);
   REGISTERS_reg_12_21_inst : DFF_X1 port map( D => n2240, CK => CLK, Q => 
                           n_1322, QN => n9192);
   REGISTERS_reg_12_20_inst : DFF_X1 port map( D => n2239, CK => CLK, Q => 
                           n_1323, QN => n9193);
   REGISTERS_reg_12_19_inst : DFF_X1 port map( D => n2238, CK => CLK, Q => 
                           n_1324, QN => n9194);
   REGISTERS_reg_12_18_inst : DFF_X1 port map( D => n2237, CK => CLK, Q => 
                           n_1325, QN => n9195);
   REGISTERS_reg_12_17_inst : DFF_X1 port map( D => n2236, CK => CLK, Q => 
                           n_1326, QN => n9196);
   REGISTERS_reg_12_16_inst : DFF_X1 port map( D => n2235, CK => CLK, Q => 
                           n_1327, QN => n9197);
   REGISTERS_reg_12_15_inst : DFF_X1 port map( D => n2234, CK => CLK, Q => 
                           n_1328, QN => n9198);
   REGISTERS_reg_12_14_inst : DFF_X1 port map( D => n2233, CK => CLK, Q => 
                           n_1329, QN => n9199);
   REGISTERS_reg_12_13_inst : DFF_X1 port map( D => n2232, CK => CLK, Q => 
                           n_1330, QN => n9200);
   REGISTERS_reg_12_12_inst : DFF_X1 port map( D => n2231, CK => CLK, Q => 
                           n_1331, QN => n9201);
   REGISTERS_reg_12_11_inst : DFF_X1 port map( D => n2230, CK => CLK, Q => 
                           n_1332, QN => n9202);
   REGISTERS_reg_12_10_inst : DFF_X1 port map( D => n2229, CK => CLK, Q => 
                           n_1333, QN => n9203);
   REGISTERS_reg_12_9_inst : DFF_X1 port map( D => n2228, CK => CLK, Q => 
                           n_1334, QN => n9204);
   REGISTERS_reg_12_8_inst : DFF_X1 port map( D => n2227, CK => CLK, Q => 
                           n_1335, QN => n9205);
   REGISTERS_reg_12_7_inst : DFF_X1 port map( D => n2226, CK => CLK, Q => 
                           n_1336, QN => n9206);
   REGISTERS_reg_12_6_inst : DFF_X1 port map( D => n2225, CK => CLK, Q => 
                           n_1337, QN => n9207);
   REGISTERS_reg_12_5_inst : DFF_X1 port map( D => n2224, CK => CLK, Q => 
                           n_1338, QN => n9208);
   REGISTERS_reg_12_4_inst : DFF_X1 port map( D => n2223, CK => CLK, Q => 
                           n_1339, QN => n9209);
   REGISTERS_reg_12_3_inst : DFF_X1 port map( D => n2222, CK => CLK, Q => 
                           n_1340, QN => n9210);
   REGISTERS_reg_12_2_inst : DFF_X1 port map( D => n2221, CK => CLK, Q => 
                           n_1341, QN => n9211);
   REGISTERS_reg_12_1_inst : DFF_X1 port map( D => n2220, CK => CLK, Q => 
                           n_1342, QN => n9212);
   REGISTERS_reg_12_0_inst : DFF_X1 port map( D => n2219, CK => CLK, Q => 
                           n_1343, QN => n9213);
   REGISTERS_reg_11_23_inst : DFF_X1 port map( D => n2274, CK => CLK, Q => 
                           n_1344, QN => n9158);
   REGISTERS_reg_11_22_inst : DFF_X1 port map( D => n2273, CK => CLK, Q => 
                           n_1345, QN => n9159);
   REGISTERS_reg_11_21_inst : DFF_X1 port map( D => n2272, CK => CLK, Q => 
                           n_1346, QN => n9160);
   REGISTERS_reg_11_20_inst : DFF_X1 port map( D => n2271, CK => CLK, Q => 
                           n_1347, QN => n9161);
   REGISTERS_reg_11_19_inst : DFF_X1 port map( D => n2270, CK => CLK, Q => 
                           n_1348, QN => n9162);
   REGISTERS_reg_11_18_inst : DFF_X1 port map( D => n2269, CK => CLK, Q => 
                           n_1349, QN => n9163);
   REGISTERS_reg_11_17_inst : DFF_X1 port map( D => n2268, CK => CLK, Q => 
                           n_1350, QN => n9164);
   REGISTERS_reg_11_16_inst : DFF_X1 port map( D => n2267, CK => CLK, Q => 
                           n_1351, QN => n9165);
   REGISTERS_reg_11_15_inst : DFF_X1 port map( D => n2266, CK => CLK, Q => 
                           n_1352, QN => n9166);
   REGISTERS_reg_11_14_inst : DFF_X1 port map( D => n2265, CK => CLK, Q => 
                           n_1353, QN => n9167);
   REGISTERS_reg_11_13_inst : DFF_X1 port map( D => n2264, CK => CLK, Q => 
                           n_1354, QN => n9168);
   REGISTERS_reg_11_12_inst : DFF_X1 port map( D => n2263, CK => CLK, Q => 
                           n_1355, QN => n9169);
   REGISTERS_reg_11_11_inst : DFF_X1 port map( D => n2262, CK => CLK, Q => 
                           n_1356, QN => n9170);
   REGISTERS_reg_11_10_inst : DFF_X1 port map( D => n2261, CK => CLK, Q => 
                           n_1357, QN => n9171);
   REGISTERS_reg_11_9_inst : DFF_X1 port map( D => n2260, CK => CLK, Q => 
                           n_1358, QN => n9172);
   REGISTERS_reg_11_8_inst : DFF_X1 port map( D => n2259, CK => CLK, Q => 
                           n_1359, QN => n9173);
   REGISTERS_reg_11_7_inst : DFF_X1 port map( D => n2258, CK => CLK, Q => 
                           n_1360, QN => n9174);
   REGISTERS_reg_11_6_inst : DFF_X1 port map( D => n2257, CK => CLK, Q => 
                           n_1361, QN => n9175);
   REGISTERS_reg_11_5_inst : DFF_X1 port map( D => n2256, CK => CLK, Q => 
                           n_1362, QN => n9176);
   REGISTERS_reg_11_4_inst : DFF_X1 port map( D => n2255, CK => CLK, Q => 
                           n_1363, QN => n9177);
   REGISTERS_reg_11_3_inst : DFF_X1 port map( D => n2254, CK => CLK, Q => 
                           n_1364, QN => n9178);
   REGISTERS_reg_11_2_inst : DFF_X1 port map( D => n2253, CK => CLK, Q => 
                           n_1365, QN => n9179);
   REGISTERS_reg_11_1_inst : DFF_X1 port map( D => n2252, CK => CLK, Q => 
                           n_1366, QN => n9180);
   REGISTERS_reg_11_0_inst : DFF_X1 port map( D => n2251, CK => CLK, Q => 
                           n_1367, QN => n9181);
   REGISTERS_reg_2_23_inst : DFF_X1 port map( D => n2562, CK => CLK, Q => 
                           n_1368, QN => n8870);
   REGISTERS_reg_2_22_inst : DFF_X1 port map( D => n2561, CK => CLK, Q => 
                           n_1369, QN => n8871);
   REGISTERS_reg_2_21_inst : DFF_X1 port map( D => n2560, CK => CLK, Q => 
                           n_1370, QN => n8872);
   REGISTERS_reg_2_20_inst : DFF_X1 port map( D => n2559, CK => CLK, Q => 
                           n_1371, QN => n8873);
   REGISTERS_reg_2_19_inst : DFF_X1 port map( D => n2558, CK => CLK, Q => 
                           n_1372, QN => n8874);
   REGISTERS_reg_2_18_inst : DFF_X1 port map( D => n2557, CK => CLK, Q => 
                           n_1373, QN => n8875);
   REGISTERS_reg_2_17_inst : DFF_X1 port map( D => n2556, CK => CLK, Q => 
                           n_1374, QN => n8876);
   REGISTERS_reg_2_16_inst : DFF_X1 port map( D => n2555, CK => CLK, Q => 
                           n_1375, QN => n8877);
   REGISTERS_reg_2_15_inst : DFF_X1 port map( D => n2554, CK => CLK, Q => 
                           n_1376, QN => n8878);
   REGISTERS_reg_2_14_inst : DFF_X1 port map( D => n2553, CK => CLK, Q => 
                           n_1377, QN => n8879);
   REGISTERS_reg_2_13_inst : DFF_X1 port map( D => n2552, CK => CLK, Q => 
                           n_1378, QN => n8880);
   REGISTERS_reg_2_12_inst : DFF_X1 port map( D => n2551, CK => CLK, Q => 
                           n_1379, QN => n8881);
   REGISTERS_reg_2_11_inst : DFF_X1 port map( D => n2550, CK => CLK, Q => 
                           n_1380, QN => n8882);
   REGISTERS_reg_2_10_inst : DFF_X1 port map( D => n2549, CK => CLK, Q => 
                           n_1381, QN => n8883);
   REGISTERS_reg_2_9_inst : DFF_X1 port map( D => n2548, CK => CLK, Q => n_1382
                           , QN => n8884);
   REGISTERS_reg_2_8_inst : DFF_X1 port map( D => n2547, CK => CLK, Q => n_1383
                           , QN => n8885);
   REGISTERS_reg_2_7_inst : DFF_X1 port map( D => n2546, CK => CLK, Q => n_1384
                           , QN => n8886);
   REGISTERS_reg_2_6_inst : DFF_X1 port map( D => n2545, CK => CLK, Q => n_1385
                           , QN => n8887);
   REGISTERS_reg_2_5_inst : DFF_X1 port map( D => n2544, CK => CLK, Q => n_1386
                           , QN => n8888);
   REGISTERS_reg_2_4_inst : DFF_X1 port map( D => n2543, CK => CLK, Q => n_1387
                           , QN => n8889);
   REGISTERS_reg_2_3_inst : DFF_X1 port map( D => n2542, CK => CLK, Q => n_1388
                           , QN => n8890);
   REGISTERS_reg_2_2_inst : DFF_X1 port map( D => n2541, CK => CLK, Q => n_1389
                           , QN => n8891);
   REGISTERS_reg_2_1_inst : DFF_X1 port map( D => n2540, CK => CLK, Q => n_1390
                           , QN => n8892);
   REGISTERS_reg_2_0_inst : DFF_X1 port map( D => n2539, CK => CLK, Q => n_1391
                           , QN => n8893);
   REGISTERS_reg_1_23_inst : DFF_X1 port map( D => n2594, CK => CLK, Q => 
                           n_1392, QN => n8838);
   REGISTERS_reg_1_22_inst : DFF_X1 port map( D => n2593, CK => CLK, Q => 
                           n_1393, QN => n8839);
   REGISTERS_reg_1_21_inst : DFF_X1 port map( D => n2592, CK => CLK, Q => 
                           n_1394, QN => n8840);
   REGISTERS_reg_1_20_inst : DFF_X1 port map( D => n2591, CK => CLK, Q => 
                           n_1395, QN => n8841);
   REGISTERS_reg_1_19_inst : DFF_X1 port map( D => n2590, CK => CLK, Q => 
                           n_1396, QN => n8842);
   REGISTERS_reg_1_18_inst : DFF_X1 port map( D => n2589, CK => CLK, Q => 
                           n_1397, QN => n8843);
   REGISTERS_reg_1_17_inst : DFF_X1 port map( D => n2588, CK => CLK, Q => 
                           n_1398, QN => n8844);
   REGISTERS_reg_1_16_inst : DFF_X1 port map( D => n2587, CK => CLK, Q => 
                           n_1399, QN => n8845);
   REGISTERS_reg_1_15_inst : DFF_X1 port map( D => n2586, CK => CLK, Q => 
                           n_1400, QN => n8846);
   REGISTERS_reg_1_14_inst : DFF_X1 port map( D => n2585, CK => CLK, Q => 
                           n_1401, QN => n8847);
   REGISTERS_reg_1_13_inst : DFF_X1 port map( D => n2584, CK => CLK, Q => 
                           n_1402, QN => n8848);
   REGISTERS_reg_1_12_inst : DFF_X1 port map( D => n2583, CK => CLK, Q => 
                           n_1403, QN => n8849);
   REGISTERS_reg_1_11_inst : DFF_X1 port map( D => n2582, CK => CLK, Q => 
                           n_1404, QN => n8850);
   REGISTERS_reg_1_10_inst : DFF_X1 port map( D => n2581, CK => CLK, Q => 
                           n_1405, QN => n8851);
   REGISTERS_reg_1_9_inst : DFF_X1 port map( D => n2580, CK => CLK, Q => n_1406
                           , QN => n8852);
   REGISTERS_reg_1_8_inst : DFF_X1 port map( D => n2579, CK => CLK, Q => n_1407
                           , QN => n8853);
   REGISTERS_reg_1_7_inst : DFF_X1 port map( D => n2578, CK => CLK, Q => n_1408
                           , QN => n8854);
   REGISTERS_reg_1_6_inst : DFF_X1 port map( D => n2577, CK => CLK, Q => n_1409
                           , QN => n8855);
   REGISTERS_reg_1_5_inst : DFF_X1 port map( D => n2576, CK => CLK, Q => n_1410
                           , QN => n8856);
   REGISTERS_reg_1_4_inst : DFF_X1 port map( D => n2575, CK => CLK, Q => n_1411
                           , QN => n8857);
   REGISTERS_reg_1_3_inst : DFF_X1 port map( D => n2574, CK => CLK, Q => n_1412
                           , QN => n8858);
   REGISTERS_reg_1_2_inst : DFF_X1 port map( D => n2573, CK => CLK, Q => n_1413
                           , QN => n8859);
   REGISTERS_reg_1_1_inst : DFF_X1 port map( D => n2572, CK => CLK, Q => n_1414
                           , QN => n8860);
   REGISTERS_reg_1_0_inst : DFF_X1 port map( D => n2571, CK => CLK, Q => n_1415
                           , QN => n8861);
   REGISTERS_reg_16_23_inst : DFF_X1 port map( D => n2114, CK => CLK, Q => 
                           n_1416, QN => n9318);
   REGISTERS_reg_16_22_inst : DFF_X1 port map( D => n2113, CK => CLK, Q => 
                           n_1417, QN => n9319);
   REGISTERS_reg_16_21_inst : DFF_X1 port map( D => n2112, CK => CLK, Q => 
                           n_1418, QN => n9320);
   REGISTERS_reg_16_20_inst : DFF_X1 port map( D => n2111, CK => CLK, Q => 
                           n_1419, QN => n9321);
   REGISTERS_reg_16_19_inst : DFF_X1 port map( D => n2110, CK => CLK, Q => 
                           n_1420, QN => n9322);
   REGISTERS_reg_16_18_inst : DFF_X1 port map( D => n2109, CK => CLK, Q => 
                           n_1421, QN => n9323);
   REGISTERS_reg_16_17_inst : DFF_X1 port map( D => n2108, CK => CLK, Q => 
                           n_1422, QN => n9324);
   REGISTERS_reg_16_16_inst : DFF_X1 port map( D => n2107, CK => CLK, Q => 
                           n_1423, QN => n9325);
   REGISTERS_reg_16_15_inst : DFF_X1 port map( D => n2106, CK => CLK, Q => 
                           n_1424, QN => n9326);
   REGISTERS_reg_16_14_inst : DFF_X1 port map( D => n2105, CK => CLK, Q => 
                           n_1425, QN => n9327);
   REGISTERS_reg_16_13_inst : DFF_X1 port map( D => n2104, CK => CLK, Q => 
                           n_1426, QN => n9328);
   REGISTERS_reg_16_12_inst : DFF_X1 port map( D => n2103, CK => CLK, Q => 
                           n_1427, QN => n9329);
   REGISTERS_reg_16_11_inst : DFF_X1 port map( D => n2102, CK => CLK, Q => 
                           n_1428, QN => n9330);
   REGISTERS_reg_16_10_inst : DFF_X1 port map( D => n2101, CK => CLK, Q => 
                           n_1429, QN => n9331);
   REGISTERS_reg_16_9_inst : DFF_X1 port map( D => n2100, CK => CLK, Q => 
                           n_1430, QN => n9332);
   REGISTERS_reg_16_8_inst : DFF_X1 port map( D => n2099, CK => CLK, Q => 
                           n_1431, QN => n9333);
   REGISTERS_reg_16_7_inst : DFF_X1 port map( D => n2098, CK => CLK, Q => 
                           n_1432, QN => n9334);
   REGISTERS_reg_16_6_inst : DFF_X1 port map( D => n2097, CK => CLK, Q => 
                           n_1433, QN => n9335);
   REGISTERS_reg_16_5_inst : DFF_X1 port map( D => n2096, CK => CLK, Q => 
                           n_1434, QN => n9336);
   REGISTERS_reg_16_4_inst : DFF_X1 port map( D => n2095, CK => CLK, Q => 
                           n_1435, QN => n9337);
   REGISTERS_reg_16_3_inst : DFF_X1 port map( D => n2094, CK => CLK, Q => 
                           n_1436, QN => n9338);
   REGISTERS_reg_16_2_inst : DFF_X1 port map( D => n2093, CK => CLK, Q => 
                           n_1437, QN => n9339);
   REGISTERS_reg_16_1_inst : DFF_X1 port map( D => n2092, CK => CLK, Q => 
                           n_1438, QN => n9340);
   REGISTERS_reg_16_0_inst : DFF_X1 port map( D => n2091, CK => CLK, Q => 
                           n_1439, QN => n9341);
   REGISTERS_reg_22_23_inst : DFF_X1 port map( D => n1922, CK => CLK, Q => 
                           n_1440, QN => n9510);
   REGISTERS_reg_22_22_inst : DFF_X1 port map( D => n1921, CK => CLK, Q => 
                           n_1441, QN => n9511);
   REGISTERS_reg_22_21_inst : DFF_X1 port map( D => n1920, CK => CLK, Q => 
                           n_1442, QN => n9512);
   REGISTERS_reg_22_20_inst : DFF_X1 port map( D => n1919, CK => CLK, Q => 
                           n_1443, QN => n9513);
   REGISTERS_reg_22_19_inst : DFF_X1 port map( D => n1918, CK => CLK, Q => 
                           n_1444, QN => n9514);
   REGISTERS_reg_22_18_inst : DFF_X1 port map( D => n1917, CK => CLK, Q => 
                           n_1445, QN => n9515);
   REGISTERS_reg_22_17_inst : DFF_X1 port map( D => n1916, CK => CLK, Q => 
                           n_1446, QN => n9516);
   REGISTERS_reg_22_16_inst : DFF_X1 port map( D => n1915, CK => CLK, Q => 
                           n_1447, QN => n9517);
   REGISTERS_reg_22_15_inst : DFF_X1 port map( D => n1914, CK => CLK, Q => 
                           n_1448, QN => n9518);
   REGISTERS_reg_22_14_inst : DFF_X1 port map( D => n1913, CK => CLK, Q => 
                           n_1449, QN => n9519);
   REGISTERS_reg_22_13_inst : DFF_X1 port map( D => n1912, CK => CLK, Q => 
                           n_1450, QN => n9520);
   REGISTERS_reg_22_12_inst : DFF_X1 port map( D => n1911, CK => CLK, Q => 
                           n_1451, QN => n9521);
   REGISTERS_reg_22_11_inst : DFF_X1 port map( D => n1910, CK => CLK, Q => 
                           n_1452, QN => n9522);
   REGISTERS_reg_22_10_inst : DFF_X1 port map( D => n1909, CK => CLK, Q => 
                           n_1453, QN => n9523);
   REGISTERS_reg_22_9_inst : DFF_X1 port map( D => n1908, CK => CLK, Q => 
                           n_1454, QN => n9524);
   REGISTERS_reg_22_8_inst : DFF_X1 port map( D => n1907, CK => CLK, Q => 
                           n_1455, QN => n9525);
   REGISTERS_reg_22_7_inst : DFF_X1 port map( D => n1906, CK => CLK, Q => 
                           n_1456, QN => n9526);
   REGISTERS_reg_22_6_inst : DFF_X1 port map( D => n1905, CK => CLK, Q => 
                           n_1457, QN => n9527);
   REGISTERS_reg_22_5_inst : DFF_X1 port map( D => n1904, CK => CLK, Q => 
                           n_1458, QN => n9528);
   REGISTERS_reg_22_4_inst : DFF_X1 port map( D => n1903, CK => CLK, Q => 
                           n_1459, QN => n9529);
   REGISTERS_reg_22_3_inst : DFF_X1 port map( D => n1902, CK => CLK, Q => 
                           n_1460, QN => n9530);
   REGISTERS_reg_22_2_inst : DFF_X1 port map( D => n1901, CK => CLK, Q => 
                           n_1461, QN => n9531);
   REGISTERS_reg_22_1_inst : DFF_X1 port map( D => n1900, CK => CLK, Q => 
                           n_1462, QN => n9532);
   REGISTERS_reg_22_0_inst : DFF_X1 port map( D => n1899, CK => CLK, Q => 
                           n_1463, QN => n9533);
   REGISTERS_reg_29_23_inst : DFF_X1 port map( D => n1698, CK => CLK, Q => 
                           n_1464, QN => n9734);
   REGISTERS_reg_29_22_inst : DFF_X1 port map( D => n1697, CK => CLK, Q => 
                           n_1465, QN => n9735);
   REGISTERS_reg_29_21_inst : DFF_X1 port map( D => n1696, CK => CLK, Q => 
                           n_1466, QN => n9736);
   REGISTERS_reg_29_20_inst : DFF_X1 port map( D => n1695, CK => CLK, Q => 
                           n_1467, QN => n9737);
   REGISTERS_reg_29_19_inst : DFF_X1 port map( D => n1694, CK => CLK, Q => 
                           n_1468, QN => n9738);
   REGISTERS_reg_29_18_inst : DFF_X1 port map( D => n1693, CK => CLK, Q => 
                           n_1469, QN => n9739);
   REGISTERS_reg_29_17_inst : DFF_X1 port map( D => n1692, CK => CLK, Q => 
                           n_1470, QN => n9740);
   REGISTERS_reg_29_16_inst : DFF_X1 port map( D => n1691, CK => CLK, Q => 
                           n_1471, QN => n9741);
   REGISTERS_reg_29_15_inst : DFF_X1 port map( D => n1690, CK => CLK, Q => 
                           n_1472, QN => n9742);
   REGISTERS_reg_29_14_inst : DFF_X1 port map( D => n1689, CK => CLK, Q => 
                           n_1473, QN => n9743);
   REGISTERS_reg_29_13_inst : DFF_X1 port map( D => n1688, CK => CLK, Q => 
                           n_1474, QN => n9744);
   REGISTERS_reg_29_12_inst : DFF_X1 port map( D => n1687, CK => CLK, Q => 
                           n_1475, QN => n9745);
   REGISTERS_reg_29_11_inst : DFF_X1 port map( D => n1686, CK => CLK, Q => 
                           n_1476, QN => n9746);
   REGISTERS_reg_29_10_inst : DFF_X1 port map( D => n1685, CK => CLK, Q => 
                           n_1477, QN => n9747);
   REGISTERS_reg_29_9_inst : DFF_X1 port map( D => n1684, CK => CLK, Q => 
                           n_1478, QN => n9748);
   REGISTERS_reg_29_8_inst : DFF_X1 port map( D => n1683, CK => CLK, Q => 
                           n_1479, QN => n9749);
   REGISTERS_reg_29_7_inst : DFF_X1 port map( D => n1682, CK => CLK, Q => 
                           n_1480, QN => n9750);
   REGISTERS_reg_29_6_inst : DFF_X1 port map( D => n1681, CK => CLK, Q => 
                           n_1481, QN => n9751);
   REGISTERS_reg_29_5_inst : DFF_X1 port map( D => n1680, CK => CLK, Q => 
                           n_1482, QN => n9752);
   REGISTERS_reg_29_4_inst : DFF_X1 port map( D => n1679, CK => CLK, Q => 
                           n_1483, QN => n9753);
   REGISTERS_reg_29_3_inst : DFF_X1 port map( D => n1678, CK => CLK, Q => 
                           n_1484, QN => n9754);
   REGISTERS_reg_29_2_inst : DFF_X1 port map( D => n1677, CK => CLK, Q => 
                           n_1485, QN => n9755);
   REGISTERS_reg_29_1_inst : DFF_X1 port map( D => n1676, CK => CLK, Q => 
                           n_1486, QN => n9756);
   REGISTERS_reg_29_0_inst : DFF_X1 port map( D => n1675, CK => CLK, Q => 
                           n_1487, QN => n9757);
   REGISTERS_reg_26_23_inst : DFF_X1 port map( D => n1794, CK => CLK, Q => 
                           n_1488, QN => n9638);
   REGISTERS_reg_26_22_inst : DFF_X1 port map( D => n1793, CK => CLK, Q => 
                           n_1489, QN => n9639);
   REGISTERS_reg_26_21_inst : DFF_X1 port map( D => n1792, CK => CLK, Q => 
                           n_1490, QN => n9640);
   REGISTERS_reg_26_20_inst : DFF_X1 port map( D => n1791, CK => CLK, Q => 
                           n_1491, QN => n9641);
   REGISTERS_reg_26_19_inst : DFF_X1 port map( D => n1790, CK => CLK, Q => 
                           n_1492, QN => n9642);
   REGISTERS_reg_26_18_inst : DFF_X1 port map( D => n1789, CK => CLK, Q => 
                           n_1493, QN => n9643);
   REGISTERS_reg_26_17_inst : DFF_X1 port map( D => n1788, CK => CLK, Q => 
                           n_1494, QN => n9644);
   REGISTERS_reg_26_16_inst : DFF_X1 port map( D => n1787, CK => CLK, Q => 
                           n_1495, QN => n9645);
   REGISTERS_reg_26_15_inst : DFF_X1 port map( D => n1786, CK => CLK, Q => 
                           n_1496, QN => n9646);
   REGISTERS_reg_26_14_inst : DFF_X1 port map( D => n1785, CK => CLK, Q => 
                           n_1497, QN => n9647);
   REGISTERS_reg_26_13_inst : DFF_X1 port map( D => n1784, CK => CLK, Q => 
                           n_1498, QN => n9648);
   REGISTERS_reg_26_12_inst : DFF_X1 port map( D => n1783, CK => CLK, Q => 
                           n_1499, QN => n9649);
   REGISTERS_reg_26_11_inst : DFF_X1 port map( D => n1782, CK => CLK, Q => 
                           n_1500, QN => n9650);
   REGISTERS_reg_26_10_inst : DFF_X1 port map( D => n1781, CK => CLK, Q => 
                           n_1501, QN => n9651);
   REGISTERS_reg_26_9_inst : DFF_X1 port map( D => n1780, CK => CLK, Q => 
                           n_1502, QN => n9652);
   REGISTERS_reg_26_8_inst : DFF_X1 port map( D => n1779, CK => CLK, Q => 
                           n_1503, QN => n9653);
   REGISTERS_reg_26_7_inst : DFF_X1 port map( D => n1778, CK => CLK, Q => 
                           n_1504, QN => n9654);
   REGISTERS_reg_26_6_inst : DFF_X1 port map( D => n1777, CK => CLK, Q => 
                           n_1505, QN => n9655);
   REGISTERS_reg_26_5_inst : DFF_X1 port map( D => n1776, CK => CLK, Q => 
                           n_1506, QN => n9656);
   REGISTERS_reg_26_4_inst : DFF_X1 port map( D => n1775, CK => CLK, Q => 
                           n_1507, QN => n9657);
   REGISTERS_reg_26_3_inst : DFF_X1 port map( D => n1774, CK => CLK, Q => 
                           n_1508, QN => n9658);
   REGISTERS_reg_26_2_inst : DFF_X1 port map( D => n1773, CK => CLK, Q => 
                           n_1509, QN => n9659);
   REGISTERS_reg_26_1_inst : DFF_X1 port map( D => n1772, CK => CLK, Q => 
                           n_1510, QN => n9660);
   REGISTERS_reg_26_0_inst : DFF_X1 port map( D => n1771, CK => CLK, Q => 
                           n_1511, QN => n9661);
   REGISTERS_reg_13_31_inst : DFF_X1 port map( D => n2218, CK => CLK, Q => 
                           n11291, QN => n9214);
   REGISTERS_reg_13_30_inst : DFF_X1 port map( D => n2217, CK => CLK, Q => 
                           n11290, QN => n9215);
   REGISTERS_reg_13_29_inst : DFF_X1 port map( D => n2216, CK => CLK, Q => 
                           n11289, QN => n9216);
   REGISTERS_reg_13_28_inst : DFF_X1 port map( D => n2215, CK => CLK, Q => 
                           n11288, QN => n9217);
   REGISTERS_reg_13_27_inst : DFF_X1 port map( D => n2214, CK => CLK, Q => 
                           n11287, QN => n9218);
   REGISTERS_reg_13_26_inst : DFF_X1 port map( D => n2213, CK => CLK, Q => 
                           n11286, QN => n9219);
   REGISTERS_reg_13_25_inst : DFF_X1 port map( D => n2212, CK => CLK, Q => 
                           n11285, QN => n9220);
   REGISTERS_reg_13_24_inst : DFF_X1 port map( D => n2211, CK => CLK, Q => 
                           n11284, QN => n9221);
   REGISTERS_reg_6_31_inst : DFF_X1 port map( D => n2442, CK => CLK, Q => 
                           n11772, QN => n8990);
   REGISTERS_reg_6_30_inst : DFF_X1 port map( D => n2441, CK => CLK, Q => 
                           n11771, QN => n8991);
   REGISTERS_reg_6_29_inst : DFF_X1 port map( D => n2440, CK => CLK, Q => 
                           n11770, QN => n8992);
   REGISTERS_reg_6_28_inst : DFF_X1 port map( D => n2439, CK => CLK, Q => 
                           n11769, QN => n8993);
   REGISTERS_reg_6_27_inst : DFF_X1 port map( D => n2438, CK => CLK, Q => 
                           n11768, QN => n8994);
   REGISTERS_reg_6_26_inst : DFF_X1 port map( D => n2437, CK => CLK, Q => 
                           n11767, QN => n8995);
   REGISTERS_reg_6_25_inst : DFF_X1 port map( D => n2436, CK => CLK, Q => 
                           n11766, QN => n8996);
   REGISTERS_reg_6_24_inst : DFF_X1 port map( D => n2435, CK => CLK, Q => 
                           n11765, QN => n8997);
   REGISTERS_reg_13_23_inst : DFF_X1 port map( D => n2210, CK => CLK, Q => 
                           n11283, QN => n9222);
   REGISTERS_reg_13_22_inst : DFF_X1 port map( D => n2209, CK => CLK, Q => 
                           n11282, QN => n9223);
   REGISTERS_reg_13_21_inst : DFF_X1 port map( D => n2208, CK => CLK, Q => 
                           n11281, QN => n9224);
   REGISTERS_reg_13_20_inst : DFF_X1 port map( D => n2207, CK => CLK, Q => 
                           n11280, QN => n9225);
   REGISTERS_reg_13_19_inst : DFF_X1 port map( D => n2206, CK => CLK, Q => 
                           n11279, QN => n9226);
   REGISTERS_reg_13_18_inst : DFF_X1 port map( D => n2205, CK => CLK, Q => 
                           n11278, QN => n9227);
   REGISTERS_reg_13_17_inst : DFF_X1 port map( D => n2204, CK => CLK, Q => 
                           n11277, QN => n9228);
   REGISTERS_reg_13_16_inst : DFF_X1 port map( D => n2203, CK => CLK, Q => 
                           n11276, QN => n9229);
   REGISTERS_reg_13_15_inst : DFF_X1 port map( D => n2202, CK => CLK, Q => 
                           n11275, QN => n9230);
   REGISTERS_reg_13_14_inst : DFF_X1 port map( D => n2201, CK => CLK, Q => 
                           n11274, QN => n9231);
   REGISTERS_reg_13_13_inst : DFF_X1 port map( D => n2200, CK => CLK, Q => 
                           n11273, QN => n9232);
   REGISTERS_reg_13_12_inst : DFF_X1 port map( D => n2199, CK => CLK, Q => 
                           n11272, QN => n9233);
   REGISTERS_reg_13_11_inst : DFF_X1 port map( D => n2198, CK => CLK, Q => 
                           n11271, QN => n9234);
   REGISTERS_reg_13_10_inst : DFF_X1 port map( D => n2197, CK => CLK, Q => 
                           n11270, QN => n9235);
   REGISTERS_reg_13_9_inst : DFF_X1 port map( D => n2196, CK => CLK, Q => 
                           n11269, QN => n9236);
   REGISTERS_reg_13_8_inst : DFF_X1 port map( D => n2195, CK => CLK, Q => 
                           n11268, QN => n9237);
   REGISTERS_reg_13_7_inst : DFF_X1 port map( D => n2194, CK => CLK, Q => 
                           n11267, QN => n9238);
   REGISTERS_reg_13_6_inst : DFF_X1 port map( D => n2193, CK => CLK, Q => 
                           n11266, QN => n9239);
   REGISTERS_reg_13_5_inst : DFF_X1 port map( D => n2192, CK => CLK, Q => 
                           n11265, QN => n9240);
   REGISTERS_reg_13_4_inst : DFF_X1 port map( D => n2191, CK => CLK, Q => 
                           n11264, QN => n9241);
   REGISTERS_reg_13_3_inst : DFF_X1 port map( D => n2190, CK => CLK, Q => 
                           n11263, QN => n9242);
   REGISTERS_reg_13_2_inst : DFF_X1 port map( D => n2189, CK => CLK, Q => 
                           n11262, QN => n9243);
   REGISTERS_reg_13_1_inst : DFF_X1 port map( D => n2188, CK => CLK, Q => 
                           n11261, QN => n9244);
   REGISTERS_reg_13_0_inst : DFF_X1 port map( D => n2187, CK => CLK, Q => 
                           n11260, QN => n9245);
   REGISTERS_reg_6_23_inst : DFF_X1 port map( D => n2434, CK => CLK, Q => 
                           n11764, QN => n8998);
   REGISTERS_reg_6_22_inst : DFF_X1 port map( D => n2433, CK => CLK, Q => 
                           n11763, QN => n8999);
   REGISTERS_reg_6_21_inst : DFF_X1 port map( D => n2432, CK => CLK, Q => 
                           n11762, QN => n9000);
   REGISTERS_reg_6_20_inst : DFF_X1 port map( D => n2431, CK => CLK, Q => 
                           n11761, QN => n9001);
   REGISTERS_reg_6_19_inst : DFF_X1 port map( D => n2430, CK => CLK, Q => 
                           n11760, QN => n9002);
   REGISTERS_reg_6_18_inst : DFF_X1 port map( D => n2429, CK => CLK, Q => 
                           n11759, QN => n9003);
   REGISTERS_reg_6_17_inst : DFF_X1 port map( D => n2428, CK => CLK, Q => 
                           n11758, QN => n9004);
   REGISTERS_reg_6_16_inst : DFF_X1 port map( D => n2427, CK => CLK, Q => 
                           n11757, QN => n9005);
   REGISTERS_reg_6_15_inst : DFF_X1 port map( D => n2426, CK => CLK, Q => 
                           n11756, QN => n9006);
   REGISTERS_reg_6_14_inst : DFF_X1 port map( D => n2425, CK => CLK, Q => 
                           n11755, QN => n9007);
   REGISTERS_reg_6_13_inst : DFF_X1 port map( D => n2424, CK => CLK, Q => 
                           n11754, QN => n9008);
   REGISTERS_reg_6_12_inst : DFF_X1 port map( D => n2423, CK => CLK, Q => 
                           n11753, QN => n9009);
   REGISTERS_reg_6_11_inst : DFF_X1 port map( D => n2422, CK => CLK, Q => 
                           n11752, QN => n9010);
   REGISTERS_reg_6_10_inst : DFF_X1 port map( D => n2421, CK => CLK, Q => 
                           n11751, QN => n9011);
   REGISTERS_reg_6_9_inst : DFF_X1 port map( D => n2420, CK => CLK, Q => n11750
                           , QN => n9012);
   REGISTERS_reg_6_8_inst : DFF_X1 port map( D => n2419, CK => CLK, Q => n11749
                           , QN => n9013);
   REGISTERS_reg_6_7_inst : DFF_X1 port map( D => n2418, CK => CLK, Q => n11748
                           , QN => n9014);
   REGISTERS_reg_6_6_inst : DFF_X1 port map( D => n2417, CK => CLK, Q => n11747
                           , QN => n9015);
   REGISTERS_reg_6_5_inst : DFF_X1 port map( D => n2416, CK => CLK, Q => n11746
                           , QN => n9016);
   REGISTERS_reg_6_4_inst : DFF_X1 port map( D => n2415, CK => CLK, Q => n11745
                           , QN => n9017);
   REGISTERS_reg_6_3_inst : DFF_X1 port map( D => n2414, CK => CLK, Q => n11744
                           , QN => n9018);
   REGISTERS_reg_6_2_inst : DFF_X1 port map( D => n2413, CK => CLK, Q => n11743
                           , QN => n9019);
   REGISTERS_reg_6_1_inst : DFF_X1 port map( D => n2412, CK => CLK, Q => n11742
                           , QN => n9020);
   REGISTERS_reg_6_0_inst : DFF_X1 port map( D => n2411, CK => CLK, Q => n11741
                           , QN => n9021);
   REGISTERS_reg_10_31_inst : DFF_X1 port map( D => n2314, CK => CLK, Q => 
                           n11708, QN => n9118);
   REGISTERS_reg_10_30_inst : DFF_X1 port map( D => n2313, CK => CLK, Q => 
                           n11707, QN => n9119);
   REGISTERS_reg_10_29_inst : DFF_X1 port map( D => n2312, CK => CLK, Q => 
                           n11706, QN => n9120);
   REGISTERS_reg_10_28_inst : DFF_X1 port map( D => n2311, CK => CLK, Q => 
                           n11705, QN => n9121);
   REGISTERS_reg_10_27_inst : DFF_X1 port map( D => n2310, CK => CLK, Q => 
                           n11704, QN => n9122);
   REGISTERS_reg_10_26_inst : DFF_X1 port map( D => n2309, CK => CLK, Q => 
                           n11703, QN => n9123);
   REGISTERS_reg_10_25_inst : DFF_X1 port map( D => n2308, CK => CLK, Q => 
                           n11702, QN => n9124);
   REGISTERS_reg_10_24_inst : DFF_X1 port map( D => n2307, CK => CLK, Q => 
                           n11701, QN => n9125);
   REGISTERS_reg_5_31_inst : DFF_X1 port map( D => n2474, CK => CLK, Q => 
                           n11419, QN => n8958);
   REGISTERS_reg_5_30_inst : DFF_X1 port map( D => n2473, CK => CLK, Q => 
                           n11418, QN => n8959);
   REGISTERS_reg_5_29_inst : DFF_X1 port map( D => n2472, CK => CLK, Q => 
                           n11417, QN => n8960);
   REGISTERS_reg_5_28_inst : DFF_X1 port map( D => n2471, CK => CLK, Q => 
                           n11416, QN => n8961);
   REGISTERS_reg_5_27_inst : DFF_X1 port map( D => n2470, CK => CLK, Q => 
                           n11415, QN => n8962);
   REGISTERS_reg_5_26_inst : DFF_X1 port map( D => n2469, CK => CLK, Q => 
                           n11414, QN => n8963);
   REGISTERS_reg_5_25_inst : DFF_X1 port map( D => n2468, CK => CLK, Q => 
                           n11413, QN => n8964);
   REGISTERS_reg_5_24_inst : DFF_X1 port map( D => n2467, CK => CLK, Q => 
                           n11412, QN => n8965);
   REGISTERS_reg_23_31_inst : DFF_X1 port map( D => n1898, CK => CLK, Q => 
                           n8006, QN => n9534);
   REGISTERS_reg_23_30_inst : DFF_X1 port map( D => n1897, CK => CLK, Q => 
                           n8005, QN => n9535);
   REGISTERS_reg_23_29_inst : DFF_X1 port map( D => n1896, CK => CLK, Q => 
                           n8004, QN => n9536);
   REGISTERS_reg_23_28_inst : DFF_X1 port map( D => n1895, CK => CLK, Q => 
                           n8003, QN => n9537);
   REGISTERS_reg_23_27_inst : DFF_X1 port map( D => n1894, CK => CLK, Q => 
                           n8002, QN => n9538);
   REGISTERS_reg_23_26_inst : DFF_X1 port map( D => n1893, CK => CLK, Q => 
                           n8001, QN => n9539);
   REGISTERS_reg_23_25_inst : DFF_X1 port map( D => n1892, CK => CLK, Q => 
                           n8000, QN => n9540);
   REGISTERS_reg_23_24_inst : DFF_X1 port map( D => n1891, CK => CLK, Q => 
                           n7999, QN => n9541);
   REGISTERS_reg_0_31_inst : DFF_X1 port map( D => n2634, CK => CLK, Q => 
                           n11515, QN => n8798);
   REGISTERS_reg_0_30_inst : DFF_X1 port map( D => n2633, CK => CLK, Q => 
                           n11514, QN => n8799);
   REGISTERS_reg_0_29_inst : DFF_X1 port map( D => n2632, CK => CLK, Q => 
                           n11513, QN => n8800);
   REGISTERS_reg_0_28_inst : DFF_X1 port map( D => n2631, CK => CLK, Q => 
                           n11512, QN => n8801);
   REGISTERS_reg_0_27_inst : DFF_X1 port map( D => n2630, CK => CLK, Q => 
                           n11511, QN => n8802);
   REGISTERS_reg_0_26_inst : DFF_X1 port map( D => n2629, CK => CLK, Q => 
                           n11510, QN => n8803);
   REGISTERS_reg_0_25_inst : DFF_X1 port map( D => n2628, CK => CLK, Q => 
                           n11509, QN => n8804);
   REGISTERS_reg_0_24_inst : DFF_X1 port map( D => n2627, CK => CLK, Q => 
                           n11508, QN => n8805);
   REGISTERS_reg_30_31_inst : DFF_X1 port map( D => n1674, CK => CLK, Q => 
                           n8038, QN => n9758);
   REGISTERS_reg_30_30_inst : DFF_X1 port map( D => n1673, CK => CLK, Q => 
                           n8037, QN => n9759);
   REGISTERS_reg_30_29_inst : DFF_X1 port map( D => n1672, CK => CLK, Q => 
                           n8036, QN => n9760);
   REGISTERS_reg_30_28_inst : DFF_X1 port map( D => n1671, CK => CLK, Q => 
                           n8035, QN => n9761);
   REGISTERS_reg_30_27_inst : DFF_X1 port map( D => n1670, CK => CLK, Q => 
                           n8034, QN => n9762);
   REGISTERS_reg_30_26_inst : DFF_X1 port map( D => n1669, CK => CLK, Q => 
                           n8033, QN => n9763);
   REGISTERS_reg_30_25_inst : DFF_X1 port map( D => n1668, CK => CLK, Q => 
                           n8032, QN => n9764);
   REGISTERS_reg_30_24_inst : DFF_X1 port map( D => n1667, CK => CLK, Q => 
                           n8031, QN => n9765);
   REGISTERS_reg_17_31_inst : DFF_X1 port map( D => n2090, CK => CLK, Q => 
                           n11580, QN => n9342);
   REGISTERS_reg_17_30_inst : DFF_X1 port map( D => n2089, CK => CLK, Q => 
                           n11579, QN => n9343);
   REGISTERS_reg_17_29_inst : DFF_X1 port map( D => n2088, CK => CLK, Q => 
                           n11578, QN => n9344);
   REGISTERS_reg_17_28_inst : DFF_X1 port map( D => n2087, CK => CLK, Q => 
                           n11577, QN => n9345);
   REGISTERS_reg_17_27_inst : DFF_X1 port map( D => n2086, CK => CLK, Q => 
                           n11576, QN => n9346);
   REGISTERS_reg_17_26_inst : DFF_X1 port map( D => n2085, CK => CLK, Q => 
                           n11575, QN => n9347);
   REGISTERS_reg_17_25_inst : DFF_X1 port map( D => n2084, CK => CLK, Q => 
                           n11574, QN => n9348);
   REGISTERS_reg_17_24_inst : DFF_X1 port map( D => n2083, CK => CLK, Q => 
                           n11573, QN => n9349);
   REGISTERS_reg_10_23_inst : DFF_X1 port map( D => n2306, CK => CLK, Q => 
                           n11700, QN => n9126);
   REGISTERS_reg_10_22_inst : DFF_X1 port map( D => n2305, CK => CLK, Q => 
                           n11699, QN => n9127);
   REGISTERS_reg_10_21_inst : DFF_X1 port map( D => n2304, CK => CLK, Q => 
                           n11698, QN => n9128);
   REGISTERS_reg_10_20_inst : DFF_X1 port map( D => n2303, CK => CLK, Q => 
                           n11697, QN => n9129);
   REGISTERS_reg_10_19_inst : DFF_X1 port map( D => n2302, CK => CLK, Q => 
                           n11696, QN => n9130);
   REGISTERS_reg_10_18_inst : DFF_X1 port map( D => n2301, CK => CLK, Q => 
                           n11695, QN => n9131);
   REGISTERS_reg_10_17_inst : DFF_X1 port map( D => n2300, CK => CLK, Q => 
                           n11694, QN => n9132);
   REGISTERS_reg_10_16_inst : DFF_X1 port map( D => n2299, CK => CLK, Q => 
                           n11693, QN => n9133);
   REGISTERS_reg_10_15_inst : DFF_X1 port map( D => n2298, CK => CLK, Q => 
                           n11692, QN => n9134);
   REGISTERS_reg_10_14_inst : DFF_X1 port map( D => n2297, CK => CLK, Q => 
                           n11691, QN => n9135);
   REGISTERS_reg_10_13_inst : DFF_X1 port map( D => n2296, CK => CLK, Q => 
                           n11690, QN => n9136);
   REGISTERS_reg_10_12_inst : DFF_X1 port map( D => n2295, CK => CLK, Q => 
                           n11689, QN => n9137);
   REGISTERS_reg_10_11_inst : DFF_X1 port map( D => n2294, CK => CLK, Q => 
                           n11688, QN => n9138);
   REGISTERS_reg_10_10_inst : DFF_X1 port map( D => n2293, CK => CLK, Q => 
                           n11687, QN => n9139);
   REGISTERS_reg_10_9_inst : DFF_X1 port map( D => n2292, CK => CLK, Q => 
                           n11686, QN => n9140);
   REGISTERS_reg_10_8_inst : DFF_X1 port map( D => n2291, CK => CLK, Q => 
                           n11685, QN => n9141);
   REGISTERS_reg_10_7_inst : DFF_X1 port map( D => n2290, CK => CLK, Q => 
                           n11684, QN => n9142);
   REGISTERS_reg_10_6_inst : DFF_X1 port map( D => n2289, CK => CLK, Q => 
                           n11683, QN => n9143);
   REGISTERS_reg_10_5_inst : DFF_X1 port map( D => n2288, CK => CLK, Q => 
                           n11682, QN => n9144);
   REGISTERS_reg_10_4_inst : DFF_X1 port map( D => n2287, CK => CLK, Q => 
                           n11681, QN => n9145);
   REGISTERS_reg_10_3_inst : DFF_X1 port map( D => n2286, CK => CLK, Q => 
                           n11680, QN => n9146);
   REGISTERS_reg_10_2_inst : DFF_X1 port map( D => n2285, CK => CLK, Q => 
                           n11679, QN => n9147);
   REGISTERS_reg_10_1_inst : DFF_X1 port map( D => n2284, CK => CLK, Q => 
                           n11678, QN => n9148);
   REGISTERS_reg_10_0_inst : DFF_X1 port map( D => n2283, CK => CLK, Q => 
                           n11677, QN => n9149);
   REGISTERS_reg_5_23_inst : DFF_X1 port map( D => n2466, CK => CLK, Q => 
                           n11411, QN => n8966);
   REGISTERS_reg_5_22_inst : DFF_X1 port map( D => n2465, CK => CLK, Q => 
                           n11410, QN => n8967);
   REGISTERS_reg_5_21_inst : DFF_X1 port map( D => n2464, CK => CLK, Q => 
                           n11409, QN => n8968);
   REGISTERS_reg_5_20_inst : DFF_X1 port map( D => n2463, CK => CLK, Q => 
                           n11408, QN => n8969);
   REGISTERS_reg_5_19_inst : DFF_X1 port map( D => n2462, CK => CLK, Q => 
                           n11407, QN => n8970);
   REGISTERS_reg_5_18_inst : DFF_X1 port map( D => n2461, CK => CLK, Q => 
                           n11406, QN => n8971);
   REGISTERS_reg_5_17_inst : DFF_X1 port map( D => n2460, CK => CLK, Q => 
                           n11405, QN => n8972);
   REGISTERS_reg_5_16_inst : DFF_X1 port map( D => n2459, CK => CLK, Q => 
                           n11404, QN => n8973);
   REGISTERS_reg_5_15_inst : DFF_X1 port map( D => n2458, CK => CLK, Q => 
                           n11403, QN => n8974);
   REGISTERS_reg_5_14_inst : DFF_X1 port map( D => n2457, CK => CLK, Q => 
                           n11402, QN => n8975);
   REGISTERS_reg_5_13_inst : DFF_X1 port map( D => n2456, CK => CLK, Q => 
                           n11401, QN => n8976);
   REGISTERS_reg_5_12_inst : DFF_X1 port map( D => n2455, CK => CLK, Q => 
                           n11400, QN => n8977);
   REGISTERS_reg_5_11_inst : DFF_X1 port map( D => n2454, CK => CLK, Q => 
                           n11399, QN => n8978);
   REGISTERS_reg_5_10_inst : DFF_X1 port map( D => n2453, CK => CLK, Q => 
                           n11398, QN => n8979);
   REGISTERS_reg_5_9_inst : DFF_X1 port map( D => n2452, CK => CLK, Q => n11397
                           , QN => n8980);
   REGISTERS_reg_5_8_inst : DFF_X1 port map( D => n2451, CK => CLK, Q => n11396
                           , QN => n8981);
   REGISTERS_reg_5_7_inst : DFF_X1 port map( D => n2450, CK => CLK, Q => n11395
                           , QN => n8982);
   REGISTERS_reg_5_6_inst : DFF_X1 port map( D => n2449, CK => CLK, Q => n11394
                           , QN => n8983);
   REGISTERS_reg_5_5_inst : DFF_X1 port map( D => n2448, CK => CLK, Q => n11393
                           , QN => n8984);
   REGISTERS_reg_5_4_inst : DFF_X1 port map( D => n2447, CK => CLK, Q => n11392
                           , QN => n8985);
   REGISTERS_reg_5_3_inst : DFF_X1 port map( D => n2446, CK => CLK, Q => n11391
                           , QN => n8986);
   REGISTERS_reg_5_2_inst : DFF_X1 port map( D => n2445, CK => CLK, Q => n11390
                           , QN => n8987);
   REGISTERS_reg_5_1_inst : DFF_X1 port map( D => n2444, CK => CLK, Q => n11389
                           , QN => n8988);
   REGISTERS_reg_5_0_inst : DFF_X1 port map( D => n2443, CK => CLK, Q => n11388
                           , QN => n8989);
   REGISTERS_reg_23_23_inst : DFF_X1 port map( D => n1890, CK => CLK, Q => 
                           n7998, QN => n9542);
   REGISTERS_reg_23_22_inst : DFF_X1 port map( D => n1889, CK => CLK, Q => 
                           n7997, QN => n9543);
   REGISTERS_reg_23_21_inst : DFF_X1 port map( D => n1888, CK => CLK, Q => 
                           n7996, QN => n9544);
   REGISTERS_reg_23_20_inst : DFF_X1 port map( D => n1887, CK => CLK, Q => 
                           n7995, QN => n9545);
   REGISTERS_reg_23_19_inst : DFF_X1 port map( D => n1886, CK => CLK, Q => 
                           n7994, QN => n9546);
   REGISTERS_reg_23_18_inst : DFF_X1 port map( D => n1885, CK => CLK, Q => 
                           n7993, QN => n9547);
   REGISTERS_reg_23_17_inst : DFF_X1 port map( D => n1884, CK => CLK, Q => 
                           n7992, QN => n9548);
   REGISTERS_reg_23_16_inst : DFF_X1 port map( D => n1883, CK => CLK, Q => 
                           n7991, QN => n9549);
   REGISTERS_reg_23_15_inst : DFF_X1 port map( D => n1882, CK => CLK, Q => 
                           n7990, QN => n9550);
   REGISTERS_reg_23_14_inst : DFF_X1 port map( D => n1881, CK => CLK, Q => 
                           n7989, QN => n9551);
   REGISTERS_reg_23_13_inst : DFF_X1 port map( D => n1880, CK => CLK, Q => 
                           n7988, QN => n9552);
   REGISTERS_reg_23_12_inst : DFF_X1 port map( D => n1879, CK => CLK, Q => 
                           n7987, QN => n9553);
   REGISTERS_reg_23_11_inst : DFF_X1 port map( D => n1878, CK => CLK, Q => 
                           n7986, QN => n9554);
   REGISTERS_reg_23_10_inst : DFF_X1 port map( D => n1877, CK => CLK, Q => 
                           n7985, QN => n9555);
   REGISTERS_reg_23_9_inst : DFF_X1 port map( D => n1876, CK => CLK, Q => n7984
                           , QN => n9556);
   REGISTERS_reg_23_8_inst : DFF_X1 port map( D => n1875, CK => CLK, Q => n7983
                           , QN => n9557);
   REGISTERS_reg_23_7_inst : DFF_X1 port map( D => n1874, CK => CLK, Q => n7982
                           , QN => n9558);
   REGISTERS_reg_23_6_inst : DFF_X1 port map( D => n1873, CK => CLK, Q => n7981
                           , QN => n9559);
   REGISTERS_reg_23_5_inst : DFF_X1 port map( D => n1872, CK => CLK, Q => n7980
                           , QN => n9560);
   REGISTERS_reg_23_4_inst : DFF_X1 port map( D => n1871, CK => CLK, Q => n7979
                           , QN => n9561);
   REGISTERS_reg_23_3_inst : DFF_X1 port map( D => n1870, CK => CLK, Q => n7978
                           , QN => n9562);
   REGISTERS_reg_23_2_inst : DFF_X1 port map( D => n1869, CK => CLK, Q => n7977
                           , QN => n9563);
   REGISTERS_reg_23_1_inst : DFF_X1 port map( D => n1868, CK => CLK, Q => n7976
                           , QN => n9564);
   REGISTERS_reg_23_0_inst : DFF_X1 port map( D => n1867, CK => CLK, Q => n7975
                           , QN => n9565);
   REGISTERS_reg_0_23_inst : DFF_X1 port map( D => n2626, CK => CLK, Q => 
                           n11507, QN => n8806);
   REGISTERS_reg_0_22_inst : DFF_X1 port map( D => n2625, CK => CLK, Q => 
                           n11506, QN => n8807);
   REGISTERS_reg_0_21_inst : DFF_X1 port map( D => n2624, CK => CLK, Q => 
                           n11505, QN => n8808);
   REGISTERS_reg_0_20_inst : DFF_X1 port map( D => n2623, CK => CLK, Q => 
                           n11504, QN => n8809);
   REGISTERS_reg_0_19_inst : DFF_X1 port map( D => n2622, CK => CLK, Q => 
                           n11503, QN => n8810);
   REGISTERS_reg_0_18_inst : DFF_X1 port map( D => n2621, CK => CLK, Q => 
                           n11502, QN => n8811);
   REGISTERS_reg_0_17_inst : DFF_X1 port map( D => n2620, CK => CLK, Q => 
                           n11501, QN => n8812);
   REGISTERS_reg_0_16_inst : DFF_X1 port map( D => n2619, CK => CLK, Q => 
                           n11500, QN => n8813);
   REGISTERS_reg_0_15_inst : DFF_X1 port map( D => n2618, CK => CLK, Q => 
                           n11499, QN => n8814);
   REGISTERS_reg_0_14_inst : DFF_X1 port map( D => n2617, CK => CLK, Q => 
                           n11498, QN => n8815);
   REGISTERS_reg_0_13_inst : DFF_X1 port map( D => n2616, CK => CLK, Q => 
                           n11497, QN => n8816);
   REGISTERS_reg_0_12_inst : DFF_X1 port map( D => n2615, CK => CLK, Q => 
                           n11496, QN => n8817);
   REGISTERS_reg_0_11_inst : DFF_X1 port map( D => n2614, CK => CLK, Q => 
                           n11495, QN => n8818);
   REGISTERS_reg_0_10_inst : DFF_X1 port map( D => n2613, CK => CLK, Q => 
                           n11494, QN => n8819);
   REGISTERS_reg_0_9_inst : DFF_X1 port map( D => n2612, CK => CLK, Q => n11493
                           , QN => n8820);
   REGISTERS_reg_0_8_inst : DFF_X1 port map( D => n2611, CK => CLK, Q => n11492
                           , QN => n8821);
   REGISTERS_reg_0_7_inst : DFF_X1 port map( D => n2610, CK => CLK, Q => n11491
                           , QN => n8822);
   REGISTERS_reg_0_6_inst : DFF_X1 port map( D => n2609, CK => CLK, Q => n11490
                           , QN => n8823);
   REGISTERS_reg_0_5_inst : DFF_X1 port map( D => n2608, CK => CLK, Q => n11489
                           , QN => n8824);
   REGISTERS_reg_0_4_inst : DFF_X1 port map( D => n2607, CK => CLK, Q => n11488
                           , QN => n8825);
   REGISTERS_reg_0_3_inst : DFF_X1 port map( D => n2606, CK => CLK, Q => n11487
                           , QN => n8826);
   REGISTERS_reg_0_2_inst : DFF_X1 port map( D => n2605, CK => CLK, Q => n11486
                           , QN => n8827);
   REGISTERS_reg_0_1_inst : DFF_X1 port map( D => n2604, CK => CLK, Q => n11485
                           , QN => n8828);
   REGISTERS_reg_0_0_inst : DFF_X1 port map( D => n2603, CK => CLK, Q => n11484
                           , QN => n8829);
   REGISTERS_reg_30_23_inst : DFF_X1 port map( D => n1666, CK => CLK, Q => 
                           n8030, QN => n9766);
   REGISTERS_reg_30_22_inst : DFF_X1 port map( D => n1665, CK => CLK, Q => 
                           n8029, QN => n9767);
   REGISTERS_reg_30_21_inst : DFF_X1 port map( D => n1664, CK => CLK, Q => 
                           n8028, QN => n9768);
   REGISTERS_reg_30_20_inst : DFF_X1 port map( D => n1663, CK => CLK, Q => 
                           n8027, QN => n9769);
   REGISTERS_reg_30_19_inst : DFF_X1 port map( D => n1662, CK => CLK, Q => 
                           n8026, QN => n9770);
   REGISTERS_reg_30_18_inst : DFF_X1 port map( D => n1661, CK => CLK, Q => 
                           n8025, QN => n9771);
   REGISTERS_reg_30_17_inst : DFF_X1 port map( D => n1660, CK => CLK, Q => 
                           n8024, QN => n9772);
   REGISTERS_reg_30_16_inst : DFF_X1 port map( D => n1659, CK => CLK, Q => 
                           n8023, QN => n9773);
   REGISTERS_reg_30_15_inst : DFF_X1 port map( D => n1658, CK => CLK, Q => 
                           n8022, QN => n9774);
   REGISTERS_reg_30_14_inst : DFF_X1 port map( D => n1657, CK => CLK, Q => 
                           n8021, QN => n9775);
   REGISTERS_reg_30_13_inst : DFF_X1 port map( D => n1656, CK => CLK, Q => 
                           n8020, QN => n9776);
   REGISTERS_reg_30_12_inst : DFF_X1 port map( D => n1655, CK => CLK, Q => 
                           n8019, QN => n9777);
   REGISTERS_reg_30_11_inst : DFF_X1 port map( D => n1654, CK => CLK, Q => 
                           n8018, QN => n9778);
   REGISTERS_reg_30_10_inst : DFF_X1 port map( D => n1653, CK => CLK, Q => 
                           n8017, QN => n9779);
   REGISTERS_reg_30_9_inst : DFF_X1 port map( D => n1652, CK => CLK, Q => n8016
                           , QN => n9780);
   REGISTERS_reg_30_8_inst : DFF_X1 port map( D => n1651, CK => CLK, Q => n8015
                           , QN => n9781);
   REGISTERS_reg_30_7_inst : DFF_X1 port map( D => n1650, CK => CLK, Q => n8014
                           , QN => n9782);
   REGISTERS_reg_30_6_inst : DFF_X1 port map( D => n1649, CK => CLK, Q => n8013
                           , QN => n9783);
   REGISTERS_reg_30_5_inst : DFF_X1 port map( D => n1648, CK => CLK, Q => n8012
                           , QN => n9784);
   REGISTERS_reg_30_4_inst : DFF_X1 port map( D => n1647, CK => CLK, Q => n8011
                           , QN => n9785);
   REGISTERS_reg_30_3_inst : DFF_X1 port map( D => n1646, CK => CLK, Q => n8010
                           , QN => n9786);
   REGISTERS_reg_30_2_inst : DFF_X1 port map( D => n1645, CK => CLK, Q => n8009
                           , QN => n9787);
   REGISTERS_reg_30_1_inst : DFF_X1 port map( D => n1644, CK => CLK, Q => n8008
                           , QN => n9788);
   REGISTERS_reg_30_0_inst : DFF_X1 port map( D => n1643, CK => CLK, Q => n8007
                           , QN => n9789);
   REGISTERS_reg_17_23_inst : DFF_X1 port map( D => n2082, CK => CLK, Q => 
                           n11572, QN => n9350);
   REGISTERS_reg_17_22_inst : DFF_X1 port map( D => n2081, CK => CLK, Q => 
                           n11571, QN => n9351);
   REGISTERS_reg_17_21_inst : DFF_X1 port map( D => n2080, CK => CLK, Q => 
                           n11570, QN => n9352);
   REGISTERS_reg_17_20_inst : DFF_X1 port map( D => n2079, CK => CLK, Q => 
                           n11569, QN => n9353);
   REGISTERS_reg_17_19_inst : DFF_X1 port map( D => n2078, CK => CLK, Q => 
                           n11568, QN => n9354);
   REGISTERS_reg_17_18_inst : DFF_X1 port map( D => n2077, CK => CLK, Q => 
                           n11567, QN => n9355);
   REGISTERS_reg_17_17_inst : DFF_X1 port map( D => n2076, CK => CLK, Q => 
                           n11566, QN => n9356);
   REGISTERS_reg_17_16_inst : DFF_X1 port map( D => n2075, CK => CLK, Q => 
                           n11565, QN => n9357);
   REGISTERS_reg_17_15_inst : DFF_X1 port map( D => n2074, CK => CLK, Q => 
                           n11564, QN => n9358);
   REGISTERS_reg_17_14_inst : DFF_X1 port map( D => n2073, CK => CLK, Q => 
                           n11563, QN => n9359);
   REGISTERS_reg_17_13_inst : DFF_X1 port map( D => n2072, CK => CLK, Q => 
                           n11562, QN => n9360);
   REGISTERS_reg_17_12_inst : DFF_X1 port map( D => n2071, CK => CLK, Q => 
                           n11561, QN => n9361);
   REGISTERS_reg_17_11_inst : DFF_X1 port map( D => n2070, CK => CLK, Q => 
                           n11560, QN => n9362);
   REGISTERS_reg_17_10_inst : DFF_X1 port map( D => n2069, CK => CLK, Q => 
                           n11559, QN => n9363);
   REGISTERS_reg_17_9_inst : DFF_X1 port map( D => n2068, CK => CLK, Q => 
                           n11558, QN => n9364);
   REGISTERS_reg_17_8_inst : DFF_X1 port map( D => n2067, CK => CLK, Q => 
                           n11557, QN => n9365);
   REGISTERS_reg_17_7_inst : DFF_X1 port map( D => n2066, CK => CLK, Q => 
                           n11556, QN => n9366);
   REGISTERS_reg_17_6_inst : DFF_X1 port map( D => n2065, CK => CLK, Q => 
                           n11555, QN => n9367);
   REGISTERS_reg_17_5_inst : DFF_X1 port map( D => n2064, CK => CLK, Q => 
                           n11554, QN => n9368);
   REGISTERS_reg_17_4_inst : DFF_X1 port map( D => n2063, CK => CLK, Q => 
                           n11553, QN => n9369);
   REGISTERS_reg_17_3_inst : DFF_X1 port map( D => n2062, CK => CLK, Q => 
                           n11552, QN => n9370);
   REGISTERS_reg_17_2_inst : DFF_X1 port map( D => n2061, CK => CLK, Q => 
                           n11551, QN => n9371);
   REGISTERS_reg_17_1_inst : DFF_X1 port map( D => n2060, CK => CLK, Q => 
                           n11550, QN => n9372);
   REGISTERS_reg_17_0_inst : DFF_X1 port map( D => n2059, CK => CLK, Q => 
                           n11549, QN => n9373);
   REGISTERS_reg_21_31_inst : DFF_X1 port map( D => n1962, CK => CLK, Q => 
                           n7910, QN => n9470);
   REGISTERS_reg_21_30_inst : DFF_X1 port map( D => n1961, CK => CLK, Q => 
                           n7909, QN => n9471);
   REGISTERS_reg_21_29_inst : DFF_X1 port map( D => n1960, CK => CLK, Q => 
                           n7908, QN => n9472);
   REGISTERS_reg_21_28_inst : DFF_X1 port map( D => n1959, CK => CLK, Q => 
                           n7907, QN => n9473);
   REGISTERS_reg_21_27_inst : DFF_X1 port map( D => n1958, CK => CLK, Q => 
                           n7906, QN => n9474);
   REGISTERS_reg_21_26_inst : DFF_X1 port map( D => n1957, CK => CLK, Q => 
                           n7905, QN => n9475);
   REGISTERS_reg_21_25_inst : DFF_X1 port map( D => n1956, CK => CLK, Q => 
                           n7904, QN => n9476);
   REGISTERS_reg_21_24_inst : DFF_X1 port map( D => n1955, CK => CLK, Q => 
                           n7903, QN => n9477);
   REGISTERS_reg_9_31_inst : DFF_X1 port map( D => n2346, CK => CLK, Q => 
                           n11355, QN => n9086);
   REGISTERS_reg_9_30_inst : DFF_X1 port map( D => n2345, CK => CLK, Q => 
                           n11354, QN => n9087);
   REGISTERS_reg_9_29_inst : DFF_X1 port map( D => n2344, CK => CLK, Q => 
                           n11353, QN => n9088);
   REGISTERS_reg_9_28_inst : DFF_X1 port map( D => n2343, CK => CLK, Q => 
                           n11352, QN => n9089);
   REGISTERS_reg_9_27_inst : DFF_X1 port map( D => n2342, CK => CLK, Q => 
                           n11351, QN => n9090);
   REGISTERS_reg_9_26_inst : DFF_X1 port map( D => n2341, CK => CLK, Q => 
                           n11350, QN => n9091);
   REGISTERS_reg_9_25_inst : DFF_X1 port map( D => n2340, CK => CLK, Q => 
                           n11349, QN => n9092);
   REGISTERS_reg_9_24_inst : DFF_X1 port map( D => n2339, CK => CLK, Q => 
                           n11348, QN => n9093);
   REGISTERS_reg_14_31_inst : DFF_X1 port map( D => n2186, CK => CLK, Q => 
                           n11644, QN => n9246);
   REGISTERS_reg_14_30_inst : DFF_X1 port map( D => n2185, CK => CLK, Q => 
                           n11643, QN => n9247);
   REGISTERS_reg_14_29_inst : DFF_X1 port map( D => n2184, CK => CLK, Q => 
                           n11642, QN => n9248);
   REGISTERS_reg_14_28_inst : DFF_X1 port map( D => n2183, CK => CLK, Q => 
                           n11641, QN => n9249);
   REGISTERS_reg_14_27_inst : DFF_X1 port map( D => n2182, CK => CLK, Q => 
                           n11640, QN => n9250);
   REGISTERS_reg_14_26_inst : DFF_X1 port map( D => n2181, CK => CLK, Q => 
                           n11639, QN => n9251);
   REGISTERS_reg_14_25_inst : DFF_X1 port map( D => n2180, CK => CLK, Q => 
                           n11638, QN => n9252);
   REGISTERS_reg_14_24_inst : DFF_X1 port map( D => n2179, CK => CLK, Q => 
                           n11637, QN => n9253);
   REGISTERS_reg_7_31_inst : DFF_X1 port map( D => n2410, CK => CLK, Q => 
                           n11740, QN => n9022);
   REGISTERS_reg_7_30_inst : DFF_X1 port map( D => n2409, CK => CLK, Q => 
                           n11739, QN => n9023);
   REGISTERS_reg_7_29_inst : DFF_X1 port map( D => n2408, CK => CLK, Q => 
                           n11738, QN => n9024);
   REGISTERS_reg_7_28_inst : DFF_X1 port map( D => n2407, CK => CLK, Q => 
                           n11737, QN => n9025);
   REGISTERS_reg_7_27_inst : DFF_X1 port map( D => n2406, CK => CLK, Q => 
                           n11736, QN => n9026);
   REGISTERS_reg_7_26_inst : DFF_X1 port map( D => n2405, CK => CLK, Q => 
                           n11735, QN => n9027);
   REGISTERS_reg_7_25_inst : DFF_X1 port map( D => n2404, CK => CLK, Q => 
                           n11734, QN => n9028);
   REGISTERS_reg_7_24_inst : DFF_X1 port map( D => n2403, CK => CLK, Q => 
                           n11733, QN => n9029);
   REGISTERS_reg_27_31_inst : DFF_X1 port map( D => n1770, CK => CLK, Q => 
                           n11548, QN => n9662);
   REGISTERS_reg_27_30_inst : DFF_X1 port map( D => n1769, CK => CLK, Q => 
                           n11547, QN => n9663);
   REGISTERS_reg_27_29_inst : DFF_X1 port map( D => n1768, CK => CLK, Q => 
                           n11546, QN => n9664);
   REGISTERS_reg_27_28_inst : DFF_X1 port map( D => n1767, CK => CLK, Q => 
                           n11545, QN => n9665);
   REGISTERS_reg_27_27_inst : DFF_X1 port map( D => n1766, CK => CLK, Q => 
                           n11544, QN => n9666);
   REGISTERS_reg_27_26_inst : DFF_X1 port map( D => n1765, CK => CLK, Q => 
                           n11543, QN => n9667);
   REGISTERS_reg_27_25_inst : DFF_X1 port map( D => n1764, CK => CLK, Q => 
                           n11542, QN => n9668);
   REGISTERS_reg_27_24_inst : DFF_X1 port map( D => n1763, CK => CLK, Q => 
                           n11541, QN => n9669);
   REGISTERS_reg_25_31_inst : DFF_X1 port map( D => n1834, CK => CLK, Q => 
                           n11227, QN => n9598);
   REGISTERS_reg_25_30_inst : DFF_X1 port map( D => n1833, CK => CLK, Q => 
                           n11226, QN => n9599);
   REGISTERS_reg_25_29_inst : DFF_X1 port map( D => n1832, CK => CLK, Q => 
                           n11225, QN => n9600);
   REGISTERS_reg_25_28_inst : DFF_X1 port map( D => n1831, CK => CLK, Q => 
                           n11224, QN => n9601);
   REGISTERS_reg_25_27_inst : DFF_X1 port map( D => n1830, CK => CLK, Q => 
                           n11223, QN => n9602);
   REGISTERS_reg_25_26_inst : DFF_X1 port map( D => n1829, CK => CLK, Q => 
                           n11222, QN => n9603);
   REGISTERS_reg_25_25_inst : DFF_X1 port map( D => n1828, CK => CLK, Q => 
                           n11221, QN => n9604);
   REGISTERS_reg_25_24_inst : DFF_X1 port map( D => n1827, CK => CLK, Q => 
                           n11220, QN => n9605);
   REGISTERS_reg_19_31_inst : DFF_X1 port map( D => n2026, CK => CLK, Q => 
                           n11259, QN => n9406);
   REGISTERS_reg_19_30_inst : DFF_X1 port map( D => n2025, CK => CLK, Q => 
                           n11258, QN => n9407);
   REGISTERS_reg_19_29_inst : DFF_X1 port map( D => n2024, CK => CLK, Q => 
                           n11257, QN => n9408);
   REGISTERS_reg_19_28_inst : DFF_X1 port map( D => n2023, CK => CLK, Q => 
                           n11256, QN => n9409);
   REGISTERS_reg_19_27_inst : DFF_X1 port map( D => n2022, CK => CLK, Q => 
                           n11255, QN => n9410);
   REGISTERS_reg_19_26_inst : DFF_X1 port map( D => n2021, CK => CLK, Q => 
                           n11254, QN => n9411);
   REGISTERS_reg_19_25_inst : DFF_X1 port map( D => n2020, CK => CLK, Q => 
                           n11253, QN => n9412);
   REGISTERS_reg_19_24_inst : DFF_X1 port map( D => n2019, CK => CLK, Q => 
                           n11252, QN => n9413);
   REGISTERS_reg_21_23_inst : DFF_X1 port map( D => n1954, CK => CLK, Q => 
                           n7902, QN => n9478);
   REGISTERS_reg_21_22_inst : DFF_X1 port map( D => n1953, CK => CLK, Q => 
                           n7901, QN => n9479);
   REGISTERS_reg_21_21_inst : DFF_X1 port map( D => n1952, CK => CLK, Q => 
                           n7900, QN => n9480);
   REGISTERS_reg_21_20_inst : DFF_X1 port map( D => n1951, CK => CLK, Q => 
                           n7899, QN => n9481);
   REGISTERS_reg_21_19_inst : DFF_X1 port map( D => n1950, CK => CLK, Q => 
                           n7898, QN => n9482);
   REGISTERS_reg_21_18_inst : DFF_X1 port map( D => n1949, CK => CLK, Q => 
                           n7897, QN => n9483);
   REGISTERS_reg_21_17_inst : DFF_X1 port map( D => n1948, CK => CLK, Q => 
                           n7896, QN => n9484);
   REGISTERS_reg_21_16_inst : DFF_X1 port map( D => n1947, CK => CLK, Q => 
                           n7895, QN => n9485);
   REGISTERS_reg_21_15_inst : DFF_X1 port map( D => n1946, CK => CLK, Q => 
                           n7894, QN => n9486);
   REGISTERS_reg_21_14_inst : DFF_X1 port map( D => n1945, CK => CLK, Q => 
                           n7893, QN => n9487);
   REGISTERS_reg_21_13_inst : DFF_X1 port map( D => n1944, CK => CLK, Q => 
                           n7892, QN => n9488);
   REGISTERS_reg_21_12_inst : DFF_X1 port map( D => n1943, CK => CLK, Q => 
                           n7891, QN => n9489);
   REGISTERS_reg_21_11_inst : DFF_X1 port map( D => n1942, CK => CLK, Q => 
                           n7890, QN => n9490);
   REGISTERS_reg_21_10_inst : DFF_X1 port map( D => n1941, CK => CLK, Q => 
                           n7889, QN => n9491);
   REGISTERS_reg_21_9_inst : DFF_X1 port map( D => n1940, CK => CLK, Q => n7888
                           , QN => n9492);
   REGISTERS_reg_21_8_inst : DFF_X1 port map( D => n1939, CK => CLK, Q => n7887
                           , QN => n9493);
   REGISTERS_reg_21_7_inst : DFF_X1 port map( D => n1938, CK => CLK, Q => n7886
                           , QN => n9494);
   REGISTERS_reg_21_6_inst : DFF_X1 port map( D => n1937, CK => CLK, Q => n7885
                           , QN => n9495);
   REGISTERS_reg_21_5_inst : DFF_X1 port map( D => n1936, CK => CLK, Q => n7884
                           , QN => n9496);
   REGISTERS_reg_21_4_inst : DFF_X1 port map( D => n1935, CK => CLK, Q => n7883
                           , QN => n9497);
   REGISTERS_reg_21_3_inst : DFF_X1 port map( D => n1934, CK => CLK, Q => n7882
                           , QN => n9498);
   REGISTERS_reg_21_2_inst : DFF_X1 port map( D => n1933, CK => CLK, Q => n7881
                           , QN => n9499);
   REGISTERS_reg_21_1_inst : DFF_X1 port map( D => n1932, CK => CLK, Q => n7880
                           , QN => n9500);
   REGISTERS_reg_21_0_inst : DFF_X1 port map( D => n1931, CK => CLK, Q => n7879
                           , QN => n9501);
   REGISTERS_reg_9_23_inst : DFF_X1 port map( D => n2338, CK => CLK, Q => 
                           n11347, QN => n9094);
   REGISTERS_reg_9_22_inst : DFF_X1 port map( D => n2337, CK => CLK, Q => 
                           n11346, QN => n9095);
   REGISTERS_reg_9_21_inst : DFF_X1 port map( D => n2336, CK => CLK, Q => 
                           n11345, QN => n9096);
   REGISTERS_reg_9_20_inst : DFF_X1 port map( D => n2335, CK => CLK, Q => 
                           n11344, QN => n9097);
   REGISTERS_reg_9_19_inst : DFF_X1 port map( D => n2334, CK => CLK, Q => 
                           n11343, QN => n9098);
   REGISTERS_reg_9_18_inst : DFF_X1 port map( D => n2333, CK => CLK, Q => 
                           n11342, QN => n9099);
   REGISTERS_reg_9_17_inst : DFF_X1 port map( D => n2332, CK => CLK, Q => 
                           n11341, QN => n9100);
   REGISTERS_reg_9_16_inst : DFF_X1 port map( D => n2331, CK => CLK, Q => 
                           n11340, QN => n9101);
   REGISTERS_reg_9_15_inst : DFF_X1 port map( D => n2330, CK => CLK, Q => 
                           n11339, QN => n9102);
   REGISTERS_reg_9_14_inst : DFF_X1 port map( D => n2329, CK => CLK, Q => 
                           n11338, QN => n9103);
   REGISTERS_reg_9_13_inst : DFF_X1 port map( D => n2328, CK => CLK, Q => 
                           n11337, QN => n9104);
   REGISTERS_reg_9_12_inst : DFF_X1 port map( D => n2327, CK => CLK, Q => 
                           n11336, QN => n9105);
   REGISTERS_reg_9_11_inst : DFF_X1 port map( D => n2326, CK => CLK, Q => 
                           n11335, QN => n9106);
   REGISTERS_reg_9_10_inst : DFF_X1 port map( D => n2325, CK => CLK, Q => 
                           n11334, QN => n9107);
   REGISTERS_reg_9_9_inst : DFF_X1 port map( D => n2324, CK => CLK, Q => n11333
                           , QN => n9108);
   REGISTERS_reg_9_8_inst : DFF_X1 port map( D => n2323, CK => CLK, Q => n11332
                           , QN => n9109);
   REGISTERS_reg_9_7_inst : DFF_X1 port map( D => n2322, CK => CLK, Q => n11331
                           , QN => n9110);
   REGISTERS_reg_9_6_inst : DFF_X1 port map( D => n2321, CK => CLK, Q => n11330
                           , QN => n9111);
   REGISTERS_reg_9_5_inst : DFF_X1 port map( D => n2320, CK => CLK, Q => n11329
                           , QN => n9112);
   REGISTERS_reg_9_4_inst : DFF_X1 port map( D => n2319, CK => CLK, Q => n11328
                           , QN => n9113);
   REGISTERS_reg_9_3_inst : DFF_X1 port map( D => n2318, CK => CLK, Q => n11327
                           , QN => n9114);
   REGISTERS_reg_9_2_inst : DFF_X1 port map( D => n2317, CK => CLK, Q => n11326
                           , QN => n9115);
   REGISTERS_reg_9_1_inst : DFF_X1 port map( D => n2316, CK => CLK, Q => n11325
                           , QN => n9116);
   REGISTERS_reg_9_0_inst : DFF_X1 port map( D => n2315, CK => CLK, Q => n11324
                           , QN => n9117);
   REGISTERS_reg_14_23_inst : DFF_X1 port map( D => n2178, CK => CLK, Q => 
                           n11636, QN => n9254);
   REGISTERS_reg_14_22_inst : DFF_X1 port map( D => n2177, CK => CLK, Q => 
                           n11635, QN => n9255);
   REGISTERS_reg_14_21_inst : DFF_X1 port map( D => n2176, CK => CLK, Q => 
                           n11634, QN => n9256);
   REGISTERS_reg_14_20_inst : DFF_X1 port map( D => n2175, CK => CLK, Q => 
                           n11633, QN => n9257);
   REGISTERS_reg_14_19_inst : DFF_X1 port map( D => n2174, CK => CLK, Q => 
                           n11632, QN => n9258);
   REGISTERS_reg_14_18_inst : DFF_X1 port map( D => n2173, CK => CLK, Q => 
                           n11631, QN => n9259);
   REGISTERS_reg_14_17_inst : DFF_X1 port map( D => n2172, CK => CLK, Q => 
                           n11630, QN => n9260);
   REGISTERS_reg_14_16_inst : DFF_X1 port map( D => n2171, CK => CLK, Q => 
                           n11629, QN => n9261);
   REGISTERS_reg_14_15_inst : DFF_X1 port map( D => n2170, CK => CLK, Q => 
                           n11628, QN => n9262);
   REGISTERS_reg_14_14_inst : DFF_X1 port map( D => n2169, CK => CLK, Q => 
                           n11627, QN => n9263);
   REGISTERS_reg_14_13_inst : DFF_X1 port map( D => n2168, CK => CLK, Q => 
                           n11626, QN => n9264);
   REGISTERS_reg_14_12_inst : DFF_X1 port map( D => n2167, CK => CLK, Q => 
                           n11625, QN => n9265);
   REGISTERS_reg_14_11_inst : DFF_X1 port map( D => n2166, CK => CLK, Q => 
                           n11624, QN => n9266);
   REGISTERS_reg_14_10_inst : DFF_X1 port map( D => n2165, CK => CLK, Q => 
                           n11623, QN => n9267);
   REGISTERS_reg_14_9_inst : DFF_X1 port map( D => n2164, CK => CLK, Q => 
                           n11622, QN => n9268);
   REGISTERS_reg_14_8_inst : DFF_X1 port map( D => n2163, CK => CLK, Q => 
                           n11621, QN => n9269);
   REGISTERS_reg_14_7_inst : DFF_X1 port map( D => n2162, CK => CLK, Q => 
                           n11620, QN => n9270);
   REGISTERS_reg_14_6_inst : DFF_X1 port map( D => n2161, CK => CLK, Q => 
                           n11619, QN => n9271);
   REGISTERS_reg_14_5_inst : DFF_X1 port map( D => n2160, CK => CLK, Q => 
                           n11618, QN => n9272);
   REGISTERS_reg_14_4_inst : DFF_X1 port map( D => n2159, CK => CLK, Q => 
                           n11617, QN => n9273);
   REGISTERS_reg_14_3_inst : DFF_X1 port map( D => n2158, CK => CLK, Q => 
                           n11616, QN => n9274);
   REGISTERS_reg_14_2_inst : DFF_X1 port map( D => n2157, CK => CLK, Q => 
                           n11615, QN => n9275);
   REGISTERS_reg_14_1_inst : DFF_X1 port map( D => n2156, CK => CLK, Q => 
                           n11614, QN => n9276);
   REGISTERS_reg_14_0_inst : DFF_X1 port map( D => n2155, CK => CLK, Q => 
                           n11613, QN => n9277);
   REGISTERS_reg_7_23_inst : DFF_X1 port map( D => n2402, CK => CLK, Q => 
                           n11732, QN => n9030);
   REGISTERS_reg_7_22_inst : DFF_X1 port map( D => n2401, CK => CLK, Q => 
                           n11731, QN => n9031);
   REGISTERS_reg_7_21_inst : DFF_X1 port map( D => n2400, CK => CLK, Q => 
                           n11730, QN => n9032);
   REGISTERS_reg_7_20_inst : DFF_X1 port map( D => n2399, CK => CLK, Q => 
                           n11729, QN => n9033);
   REGISTERS_reg_7_19_inst : DFF_X1 port map( D => n2398, CK => CLK, Q => 
                           n11728, QN => n9034);
   REGISTERS_reg_7_18_inst : DFF_X1 port map( D => n2397, CK => CLK, Q => 
                           n11727, QN => n9035);
   REGISTERS_reg_7_17_inst : DFF_X1 port map( D => n2396, CK => CLK, Q => 
                           n11726, QN => n9036);
   REGISTERS_reg_7_16_inst : DFF_X1 port map( D => n2395, CK => CLK, Q => 
                           n11725, QN => n9037);
   REGISTERS_reg_7_15_inst : DFF_X1 port map( D => n2394, CK => CLK, Q => 
                           n11724, QN => n9038);
   REGISTERS_reg_7_14_inst : DFF_X1 port map( D => n2393, CK => CLK, Q => 
                           n11723, QN => n9039);
   REGISTERS_reg_7_13_inst : DFF_X1 port map( D => n2392, CK => CLK, Q => 
                           n11722, QN => n9040);
   REGISTERS_reg_7_12_inst : DFF_X1 port map( D => n2391, CK => CLK, Q => 
                           n11721, QN => n9041);
   REGISTERS_reg_7_11_inst : DFF_X1 port map( D => n2390, CK => CLK, Q => 
                           n11720, QN => n9042);
   REGISTERS_reg_7_10_inst : DFF_X1 port map( D => n2389, CK => CLK, Q => 
                           n11719, QN => n9043);
   REGISTERS_reg_7_9_inst : DFF_X1 port map( D => n2388, CK => CLK, Q => n11718
                           , QN => n9044);
   REGISTERS_reg_7_8_inst : DFF_X1 port map( D => n2387, CK => CLK, Q => n11717
                           , QN => n9045);
   REGISTERS_reg_7_7_inst : DFF_X1 port map( D => n2386, CK => CLK, Q => n11716
                           , QN => n9046);
   REGISTERS_reg_7_6_inst : DFF_X1 port map( D => n2385, CK => CLK, Q => n11715
                           , QN => n9047);
   REGISTERS_reg_7_5_inst : DFF_X1 port map( D => n2384, CK => CLK, Q => n11714
                           , QN => n9048);
   REGISTERS_reg_7_4_inst : DFF_X1 port map( D => n2383, CK => CLK, Q => n11713
                           , QN => n9049);
   REGISTERS_reg_7_3_inst : DFF_X1 port map( D => n2382, CK => CLK, Q => n11712
                           , QN => n9050);
   REGISTERS_reg_7_2_inst : DFF_X1 port map( D => n2381, CK => CLK, Q => n11711
                           , QN => n9051);
   REGISTERS_reg_7_1_inst : DFF_X1 port map( D => n2380, CK => CLK, Q => n11710
                           , QN => n9052);
   REGISTERS_reg_7_0_inst : DFF_X1 port map( D => n2379, CK => CLK, Q => n11709
                           , QN => n9053);
   REGISTERS_reg_27_23_inst : DFF_X1 port map( D => n1762, CK => CLK, Q => 
                           n11540, QN => n9670);
   REGISTERS_reg_27_22_inst : DFF_X1 port map( D => n1761, CK => CLK, Q => 
                           n11539, QN => n9671);
   REGISTERS_reg_27_21_inst : DFF_X1 port map( D => n1760, CK => CLK, Q => 
                           n11538, QN => n9672);
   REGISTERS_reg_27_20_inst : DFF_X1 port map( D => n1759, CK => CLK, Q => 
                           n11537, QN => n9673);
   REGISTERS_reg_27_19_inst : DFF_X1 port map( D => n1758, CK => CLK, Q => 
                           n11536, QN => n9674);
   REGISTERS_reg_27_18_inst : DFF_X1 port map( D => n1757, CK => CLK, Q => 
                           n11535, QN => n9675);
   REGISTERS_reg_27_17_inst : DFF_X1 port map( D => n1756, CK => CLK, Q => 
                           n11534, QN => n9676);
   REGISTERS_reg_27_16_inst : DFF_X1 port map( D => n1755, CK => CLK, Q => 
                           n11533, QN => n9677);
   REGISTERS_reg_27_15_inst : DFF_X1 port map( D => n1754, CK => CLK, Q => 
                           n11532, QN => n9678);
   REGISTERS_reg_27_14_inst : DFF_X1 port map( D => n1753, CK => CLK, Q => 
                           n11531, QN => n9679);
   REGISTERS_reg_27_13_inst : DFF_X1 port map( D => n1752, CK => CLK, Q => 
                           n11530, QN => n9680);
   REGISTERS_reg_27_12_inst : DFF_X1 port map( D => n1751, CK => CLK, Q => 
                           n11529, QN => n9681);
   REGISTERS_reg_27_11_inst : DFF_X1 port map( D => n1750, CK => CLK, Q => 
                           n11528, QN => n9682);
   REGISTERS_reg_27_10_inst : DFF_X1 port map( D => n1749, CK => CLK, Q => 
                           n11527, QN => n9683);
   REGISTERS_reg_27_9_inst : DFF_X1 port map( D => n1748, CK => CLK, Q => 
                           n11526, QN => n9684);
   REGISTERS_reg_27_8_inst : DFF_X1 port map( D => n1747, CK => CLK, Q => 
                           n11525, QN => n9685);
   REGISTERS_reg_27_7_inst : DFF_X1 port map( D => n1746, CK => CLK, Q => 
                           n11524, QN => n9686);
   REGISTERS_reg_27_6_inst : DFF_X1 port map( D => n1745, CK => CLK, Q => 
                           n11523, QN => n9687);
   REGISTERS_reg_27_5_inst : DFF_X1 port map( D => n1744, CK => CLK, Q => 
                           n11522, QN => n9688);
   REGISTERS_reg_27_4_inst : DFF_X1 port map( D => n1743, CK => CLK, Q => 
                           n11521, QN => n9689);
   REGISTERS_reg_27_3_inst : DFF_X1 port map( D => n1742, CK => CLK, Q => 
                           n11520, QN => n9690);
   REGISTERS_reg_27_2_inst : DFF_X1 port map( D => n1741, CK => CLK, Q => 
                           n11519, QN => n9691);
   REGISTERS_reg_27_1_inst : DFF_X1 port map( D => n1740, CK => CLK, Q => 
                           n11518, QN => n9692);
   REGISTERS_reg_27_0_inst : DFF_X1 port map( D => n1739, CK => CLK, Q => 
                           n11517, QN => n9693);
   REGISTERS_reg_25_23_inst : DFF_X1 port map( D => n1826, CK => CLK, Q => 
                           n11219, QN => n9606);
   REGISTERS_reg_25_22_inst : DFF_X1 port map( D => n1825, CK => CLK, Q => 
                           n11218, QN => n9607);
   REGISTERS_reg_25_21_inst : DFF_X1 port map( D => n1824, CK => CLK, Q => 
                           n11217, QN => n9608);
   REGISTERS_reg_25_20_inst : DFF_X1 port map( D => n1823, CK => CLK, Q => 
                           n11216, QN => n9609);
   REGISTERS_reg_25_19_inst : DFF_X1 port map( D => n1822, CK => CLK, Q => 
                           n11215, QN => n9610);
   REGISTERS_reg_25_18_inst : DFF_X1 port map( D => n1821, CK => CLK, Q => 
                           n11214, QN => n9611);
   REGISTERS_reg_25_17_inst : DFF_X1 port map( D => n1820, CK => CLK, Q => 
                           n11213, QN => n9612);
   REGISTERS_reg_25_16_inst : DFF_X1 port map( D => n1819, CK => CLK, Q => 
                           n11212, QN => n9613);
   REGISTERS_reg_25_15_inst : DFF_X1 port map( D => n1818, CK => CLK, Q => 
                           n11211, QN => n9614);
   REGISTERS_reg_25_14_inst : DFF_X1 port map( D => n1817, CK => CLK, Q => 
                           n11210, QN => n9615);
   REGISTERS_reg_25_13_inst : DFF_X1 port map( D => n1816, CK => CLK, Q => 
                           n11209, QN => n9616);
   REGISTERS_reg_25_12_inst : DFF_X1 port map( D => n1815, CK => CLK, Q => 
                           n11208, QN => n9617);
   REGISTERS_reg_25_11_inst : DFF_X1 port map( D => n1814, CK => CLK, Q => 
                           n11207, QN => n9618);
   REGISTERS_reg_25_10_inst : DFF_X1 port map( D => n1813, CK => CLK, Q => 
                           n11206, QN => n9619);
   REGISTERS_reg_25_9_inst : DFF_X1 port map( D => n1812, CK => CLK, Q => 
                           n11205, QN => n9620);
   REGISTERS_reg_25_8_inst : DFF_X1 port map( D => n1811, CK => CLK, Q => 
                           n11204, QN => n9621);
   REGISTERS_reg_25_7_inst : DFF_X1 port map( D => n1810, CK => CLK, Q => 
                           n11203, QN => n9622);
   REGISTERS_reg_25_6_inst : DFF_X1 port map( D => n1809, CK => CLK, Q => 
                           n11202, QN => n9623);
   REGISTERS_reg_25_5_inst : DFF_X1 port map( D => n1808, CK => CLK, Q => 
                           n11201, QN => n9624);
   REGISTERS_reg_25_4_inst : DFF_X1 port map( D => n1807, CK => CLK, Q => 
                           n11200, QN => n9625);
   REGISTERS_reg_25_3_inst : DFF_X1 port map( D => n1806, CK => CLK, Q => 
                           n11199, QN => n9626);
   REGISTERS_reg_25_2_inst : DFF_X1 port map( D => n1805, CK => CLK, Q => 
                           n11198, QN => n9627);
   REGISTERS_reg_25_1_inst : DFF_X1 port map( D => n1804, CK => CLK, Q => 
                           n11197, QN => n9628);
   REGISTERS_reg_25_0_inst : DFF_X1 port map( D => n1803, CK => CLK, Q => 
                           n11196, QN => n9629);
   REGISTERS_reg_19_23_inst : DFF_X1 port map( D => n2018, CK => CLK, Q => 
                           n11251, QN => n9414);
   REGISTERS_reg_19_22_inst : DFF_X1 port map( D => n2017, CK => CLK, Q => 
                           n11250, QN => n9415);
   REGISTERS_reg_19_21_inst : DFF_X1 port map( D => n2016, CK => CLK, Q => 
                           n11249, QN => n9416);
   REGISTERS_reg_19_20_inst : DFF_X1 port map( D => n2015, CK => CLK, Q => 
                           n11248, QN => n9417);
   REGISTERS_reg_19_19_inst : DFF_X1 port map( D => n2014, CK => CLK, Q => 
                           n11247, QN => n9418);
   REGISTERS_reg_19_18_inst : DFF_X1 port map( D => n2013, CK => CLK, Q => 
                           n11246, QN => n9419);
   REGISTERS_reg_19_17_inst : DFF_X1 port map( D => n2012, CK => CLK, Q => 
                           n11245, QN => n9420);
   REGISTERS_reg_19_16_inst : DFF_X1 port map( D => n2011, CK => CLK, Q => 
                           n11244, QN => n9421);
   REGISTERS_reg_19_15_inst : DFF_X1 port map( D => n2010, CK => CLK, Q => 
                           n11243, QN => n9422);
   REGISTERS_reg_19_14_inst : DFF_X1 port map( D => n2009, CK => CLK, Q => 
                           n11242, QN => n9423);
   REGISTERS_reg_19_13_inst : DFF_X1 port map( D => n2008, CK => CLK, Q => 
                           n11241, QN => n9424);
   REGISTERS_reg_19_12_inst : DFF_X1 port map( D => n2007, CK => CLK, Q => 
                           n11240, QN => n9425);
   REGISTERS_reg_19_11_inst : DFF_X1 port map( D => n2006, CK => CLK, Q => 
                           n11239, QN => n9426);
   REGISTERS_reg_19_10_inst : DFF_X1 port map( D => n2005, CK => CLK, Q => 
                           n11238, QN => n9427);
   REGISTERS_reg_19_9_inst : DFF_X1 port map( D => n2004, CK => CLK, Q => 
                           n11237, QN => n9428);
   REGISTERS_reg_19_8_inst : DFF_X1 port map( D => n2003, CK => CLK, Q => 
                           n11236, QN => n9429);
   REGISTERS_reg_19_7_inst : DFF_X1 port map( D => n2002, CK => CLK, Q => 
                           n11235, QN => n9430);
   REGISTERS_reg_19_6_inst : DFF_X1 port map( D => n2001, CK => CLK, Q => 
                           n11234, QN => n9431);
   REGISTERS_reg_19_5_inst : DFF_X1 port map( D => n2000, CK => CLK, Q => 
                           n11233, QN => n9432);
   REGISTERS_reg_19_4_inst : DFF_X1 port map( D => n1999, CK => CLK, Q => 
                           n11232, QN => n9433);
   REGISTERS_reg_19_3_inst : DFF_X1 port map( D => n1998, CK => CLK, Q => 
                           n11231, QN => n9434);
   REGISTERS_reg_19_2_inst : DFF_X1 port map( D => n1997, CK => CLK, Q => 
                           n11230, QN => n9435);
   REGISTERS_reg_19_1_inst : DFF_X1 port map( D => n1996, CK => CLK, Q => 
                           n11229, QN => n9436);
   REGISTERS_reg_19_0_inst : DFF_X1 port map( D => n1995, CK => CLK, Q => 
                           n11228, QN => n9437);
   U7999 : AND3_X1 port map( A1 => n11872, A2 => n11082, A3 => RD2, ZN => 
                           n11868);
   U8000 : AND3_X1 port map( A1 => n11875, A2 => n10482, A3 => RD1, ZN => 
                           n11869);
   U8001 : BUF_X1 port map( A => n12324, Z => n12322);
   U8002 : BUF_X1 port map( A => n12512, Z => n12510);
   U8003 : BUF_X1 port map( A => n12324, Z => n12323);
   U8004 : BUF_X1 port map( A => n12512, Z => n12511);
   U8005 : BUF_X1 port map( A => n12264, Z => n12262);
   U8006 : BUF_X1 port map( A => n12268, Z => n12266);
   U8007 : BUF_X1 port map( A => n12272, Z => n12270);
   U8008 : BUF_X1 port map( A => n12276, Z => n12274);
   U8009 : BUF_X1 port map( A => n12280, Z => n12278);
   U8010 : BUF_X1 port map( A => n12284, Z => n12282);
   U8011 : BUF_X1 port map( A => n12288, Z => n12286);
   U8012 : BUF_X1 port map( A => n12292, Z => n12290);
   U8013 : BUF_X1 port map( A => n12296, Z => n12294);
   U8014 : BUF_X1 port map( A => n12300, Z => n12298);
   U8015 : BUF_X1 port map( A => n12304, Z => n12302);
   U8016 : BUF_X1 port map( A => n12308, Z => n12306);
   U8017 : BUF_X1 port map( A => n12312, Z => n12310);
   U8018 : BUF_X1 port map( A => n12316, Z => n12314);
   U8019 : BUF_X1 port map( A => n12320, Z => n12318);
   U8020 : BUF_X1 port map( A => n12328, Z => n12326);
   U8021 : BUF_X1 port map( A => n12332, Z => n12330);
   U8022 : BUF_X1 port map( A => n12336, Z => n12334);
   U8023 : BUF_X1 port map( A => n12340, Z => n12338);
   U8024 : BUF_X1 port map( A => n12344, Z => n12342);
   U8025 : BUF_X1 port map( A => n12348, Z => n12346);
   U8026 : BUF_X1 port map( A => n12352, Z => n12350);
   U8027 : BUF_X1 port map( A => n12356, Z => n12354);
   U8028 : BUF_X1 port map( A => n12360, Z => n12358);
   U8029 : BUF_X1 port map( A => n12364, Z => n12362);
   U8030 : BUF_X1 port map( A => n12368, Z => n12366);
   U8031 : BUF_X1 port map( A => n12372, Z => n12370);
   U8032 : BUF_X1 port map( A => n12376, Z => n12374);
   U8033 : BUF_X1 port map( A => n12380, Z => n12378);
   U8034 : BUF_X1 port map( A => n12384, Z => n12382);
   U8035 : BUF_X1 port map( A => n12264, Z => n12263);
   U8036 : BUF_X1 port map( A => n12268, Z => n12267);
   U8037 : BUF_X1 port map( A => n12272, Z => n12271);
   U8038 : BUF_X1 port map( A => n12276, Z => n12275);
   U8039 : BUF_X1 port map( A => n12280, Z => n12279);
   U8040 : BUF_X1 port map( A => n12284, Z => n12283);
   U8041 : BUF_X1 port map( A => n12288, Z => n12287);
   U8042 : BUF_X1 port map( A => n12292, Z => n12291);
   U8043 : BUF_X1 port map( A => n12296, Z => n12295);
   U8044 : BUF_X1 port map( A => n12300, Z => n12299);
   U8045 : BUF_X1 port map( A => n12304, Z => n12303);
   U8046 : BUF_X1 port map( A => n12308, Z => n12307);
   U8047 : BUF_X1 port map( A => n12312, Z => n12311);
   U8048 : BUF_X1 port map( A => n12316, Z => n12315);
   U8049 : BUF_X1 port map( A => n12320, Z => n12319);
   U8050 : BUF_X1 port map( A => n12328, Z => n12327);
   U8051 : BUF_X1 port map( A => n12332, Z => n12331);
   U8052 : BUF_X1 port map( A => n12336, Z => n12335);
   U8053 : BUF_X1 port map( A => n12340, Z => n12339);
   U8054 : BUF_X1 port map( A => n12344, Z => n12343);
   U8055 : BUF_X1 port map( A => n12348, Z => n12347);
   U8056 : BUF_X1 port map( A => n12352, Z => n12351);
   U8057 : BUF_X1 port map( A => n12356, Z => n12355);
   U8058 : BUF_X1 port map( A => n12360, Z => n12359);
   U8059 : BUF_X1 port map( A => n12364, Z => n12363);
   U8060 : BUF_X1 port map( A => n12368, Z => n12367);
   U8061 : BUF_X1 port map( A => n12372, Z => n12371);
   U8062 : BUF_X1 port map( A => n12376, Z => n12375);
   U8063 : BUF_X1 port map( A => n12380, Z => n12379);
   U8064 : BUF_X1 port map( A => n12384, Z => n12383);
   U8065 : BUF_X1 port map( A => n10525, Z => n12051);
   U8066 : BUF_X1 port map( A => n9925, Z => n12195);
   U8067 : BUF_X1 port map( A => n10518, Z => n12071);
   U8068 : BUF_X1 port map( A => n10519, Z => n12067);
   U8069 : BUF_X1 port map( A => n9918, Z => n12215);
   U8070 : BUF_X1 port map( A => n9919, Z => n12211);
   U8071 : BUF_X1 port map( A => n10513, Z => n12087);
   U8072 : BUF_X1 port map( A => n9913, Z => n12231);
   U8073 : BUF_X1 port map( A => n10509, Z => n12099);
   U8074 : BUF_X1 port map( A => n10508, Z => n12103);
   U8075 : BUF_X1 port map( A => n10507, Z => n12107);
   U8076 : BUF_X1 port map( A => n10514, Z => n12083);
   U8077 : BUF_X1 port map( A => n9909, Z => n12243);
   U8078 : BUF_X1 port map( A => n9908, Z => n12247);
   U8079 : BUF_X1 port map( A => n9907, Z => n12251);
   U8080 : BUF_X1 port map( A => n9914, Z => n12227);
   U8081 : BUF_X1 port map( A => n12059, Z => n12057);
   U8082 : BUF_X1 port map( A => n12203, Z => n12201);
   U8083 : BUF_X1 port map( A => n11868, Z => n12054);
   U8084 : BUF_X1 port map( A => n11869, Z => n12198);
   U8085 : BUF_X1 port map( A => n10520, Z => n12063);
   U8086 : BUF_X1 port map( A => n9920, Z => n12207);
   U8087 : BUF_X1 port map( A => n8781, Z => n12523);
   U8088 : BUF_X1 port map( A => n8781, Z => n12524);
   U8089 : BUF_X1 port map( A => n12059, Z => n12058);
   U8090 : BUF_X1 port map( A => n12203, Z => n12202);
   U8091 : BUF_X1 port map( A => n10504, Z => n12112);
   U8092 : BUF_X1 port map( A => n10505, Z => n12108);
   U8093 : BUF_X1 port map( A => n10510, Z => n12092);
   U8094 : BUF_X1 port map( A => n10511, Z => n12088);
   U8095 : BUF_X1 port map( A => n10515, Z => n12076);
   U8096 : BUF_X1 port map( A => n10516, Z => n12072);
   U8097 : BUF_X1 port map( A => n9904, Z => n12256);
   U8098 : BUF_X1 port map( A => n9905, Z => n12252);
   U8099 : BUF_X1 port map( A => n9910, Z => n12236);
   U8100 : BUF_X1 port map( A => n9911, Z => n12232);
   U8101 : BUF_X1 port map( A => n9915, Z => n12220);
   U8102 : BUF_X1 port map( A => n9916, Z => n12216);
   U8103 : BUF_X1 port map( A => n10539, Z => n12019);
   U8104 : BUF_X1 port map( A => n10540, Z => n12015);
   U8105 : BUF_X1 port map( A => n10538, Z => n12020);
   U8106 : BUF_X1 port map( A => n10550, Z => n11983);
   U8107 : BUF_X1 port map( A => n10551, Z => n11979);
   U8108 : BUF_X1 port map( A => n10549, Z => n11984);
   U8109 : BUF_X1 port map( A => n10545, Z => n11999);
   U8110 : BUF_X1 port map( A => n10544, Z => n12000);
   U8111 : BUF_X1 port map( A => n9939, Z => n12163);
   U8112 : BUF_X1 port map( A => n9940, Z => n12159);
   U8113 : BUF_X1 port map( A => n9938, Z => n12164);
   U8114 : BUF_X1 port map( A => n9950, Z => n12127);
   U8115 : BUF_X1 port map( A => n9951, Z => n12123);
   U8116 : BUF_X1 port map( A => n9949, Z => n12128);
   U8117 : BUF_X1 port map( A => n9945, Z => n12143);
   U8118 : BUF_X1 port map( A => n9944, Z => n12144);
   U8119 : BUF_X1 port map( A => n10534, Z => n12035);
   U8120 : BUF_X1 port map( A => n10533, Z => n12036);
   U8121 : BUF_X1 port map( A => n9934, Z => n12179);
   U8122 : BUF_X1 port map( A => n9933, Z => n12180);
   U8123 : BUF_X1 port map( A => n10536, Z => n12024);
   U8124 : BUF_X1 port map( A => n10535, Z => n12028);
   U8125 : BUF_X1 port map( A => n10547, Z => n11988);
   U8126 : BUF_X1 port map( A => n10546, Z => n11992);
   U8127 : BUF_X1 port map( A => n10531, Z => n12040);
   U8128 : BUF_X1 port map( A => n10530, Z => n12044);
   U8129 : BUF_X1 port map( A => n10542, Z => n12004);
   U8130 : BUF_X1 port map( A => n10541, Z => n12008);
   U8131 : BUF_X1 port map( A => n9936, Z => n12168);
   U8132 : BUF_X1 port map( A => n9935, Z => n12172);
   U8133 : BUF_X1 port map( A => n9947, Z => n12132);
   U8134 : BUF_X1 port map( A => n9946, Z => n12136);
   U8135 : BUF_X1 port map( A => n9931, Z => n12184);
   U8136 : BUF_X1 port map( A => n9930, Z => n12188);
   U8137 : BUF_X1 port map( A => n9942, Z => n12148);
   U8138 : BUF_X1 port map( A => n9941, Z => n12152);
   U8139 : BUF_X1 port map( A => n9854, Z => n12385);
   U8140 : BUF_X1 port map( A => n9853, Z => n12389);
   U8141 : BUF_X1 port map( A => n9852, Z => n12393);
   U8142 : BUF_X1 port map( A => n9851, Z => n12397);
   U8143 : BUF_X1 port map( A => n9850, Z => n12401);
   U8144 : BUF_X1 port map( A => n9849, Z => n12405);
   U8145 : BUF_X1 port map( A => n9848, Z => n12409);
   U8146 : BUF_X1 port map( A => n9847, Z => n12413);
   U8147 : BUF_X1 port map( A => n9846, Z => n12417);
   U8148 : BUF_X1 port map( A => n9845, Z => n12421);
   U8149 : BUF_X1 port map( A => n9844, Z => n12425);
   U8150 : BUF_X1 port map( A => n9843, Z => n12429);
   U8151 : BUF_X1 port map( A => n9842, Z => n12433);
   U8152 : BUF_X1 port map( A => n9841, Z => n12437);
   U8153 : BUF_X1 port map( A => n9840, Z => n12441);
   U8154 : BUF_X1 port map( A => n9839, Z => n12445);
   U8155 : BUF_X1 port map( A => n9838, Z => n12449);
   U8156 : BUF_X1 port map( A => n9837, Z => n12453);
   U8157 : BUF_X1 port map( A => n9836, Z => n12457);
   U8158 : BUF_X1 port map( A => n9835, Z => n12461);
   U8159 : BUF_X1 port map( A => n9834, Z => n12465);
   U8160 : BUF_X1 port map( A => n9833, Z => n12469);
   U8161 : BUF_X1 port map( A => n9832, Z => n12473);
   U8162 : BUF_X1 port map( A => n9831, Z => n12477);
   U8163 : BUF_X1 port map( A => n9830, Z => n12481);
   U8164 : BUF_X1 port map( A => n9829, Z => n12485);
   U8165 : BUF_X1 port map( A => n9828, Z => n12489);
   U8166 : BUF_X1 port map( A => n9827, Z => n12493);
   U8167 : BUF_X1 port map( A => n9826, Z => n12497);
   U8168 : BUF_X1 port map( A => n9825, Z => n12501);
   U8169 : BUF_X1 port map( A => n9824, Z => n12505);
   U8170 : BUF_X1 port map( A => n9822, Z => n12513);
   U8171 : BUF_X1 port map( A => n10552, Z => n11972);
   U8172 : BUF_X1 port map( A => n9952, Z => n12116);
   U8173 : BUF_X1 port map( A => n12323, Z => n11922);
   U8174 : BUF_X1 port map( A => n12323, Z => n11921);
   U8175 : BUF_X1 port map( A => n12511, Z => n11970);
   U8176 : BUF_X1 port map( A => n12511, Z => n11969);
   U8177 : INV_X1 port map( A => n12322, ZN => n12321);
   U8178 : INV_X1 port map( A => n12510, ZN => n12509);
   U8179 : BUF_X1 port map( A => n12323, Z => n11923);
   U8180 : BUF_X1 port map( A => n12511, Z => n11971);
   U8181 : BUF_X1 port map( A => n12263, Z => n11876);
   U8182 : BUF_X1 port map( A => n12263, Z => n11877);
   U8183 : BUF_X1 port map( A => n12267, Z => n11880);
   U8184 : BUF_X1 port map( A => n12267, Z => n11879);
   U8185 : BUF_X1 port map( A => n12271, Z => n11883);
   U8186 : BUF_X1 port map( A => n12271, Z => n11882);
   U8187 : BUF_X1 port map( A => n12275, Z => n11886);
   U8188 : BUF_X1 port map( A => n12275, Z => n11885);
   U8189 : BUF_X1 port map( A => n12279, Z => n11889);
   U8190 : BUF_X1 port map( A => n12279, Z => n11888);
   U8191 : BUF_X1 port map( A => n12283, Z => n11892);
   U8192 : BUF_X1 port map( A => n12283, Z => n11891);
   U8193 : BUF_X1 port map( A => n12287, Z => n11895);
   U8194 : BUF_X1 port map( A => n12287, Z => n11894);
   U8195 : BUF_X1 port map( A => n12291, Z => n11898);
   U8196 : BUF_X1 port map( A => n12291, Z => n11897);
   U8197 : BUF_X1 port map( A => n12295, Z => n11901);
   U8198 : BUF_X1 port map( A => n12295, Z => n11900);
   U8199 : BUF_X1 port map( A => n12299, Z => n11904);
   U8200 : BUF_X1 port map( A => n12299, Z => n11903);
   U8201 : BUF_X1 port map( A => n12303, Z => n11907);
   U8202 : BUF_X1 port map( A => n12303, Z => n11906);
   U8203 : BUF_X1 port map( A => n12307, Z => n11910);
   U8204 : BUF_X1 port map( A => n12307, Z => n11909);
   U8205 : BUF_X1 port map( A => n12311, Z => n11913);
   U8206 : BUF_X1 port map( A => n12311, Z => n11912);
   U8207 : BUF_X1 port map( A => n12315, Z => n11916);
   U8208 : BUF_X1 port map( A => n12315, Z => n11915);
   U8209 : BUF_X1 port map( A => n12319, Z => n11919);
   U8210 : BUF_X1 port map( A => n12319, Z => n11918);
   U8211 : BUF_X1 port map( A => n12327, Z => n11925);
   U8212 : BUF_X1 port map( A => n12327, Z => n11924);
   U8213 : BUF_X1 port map( A => n12331, Z => n11928);
   U8214 : BUF_X1 port map( A => n12331, Z => n11927);
   U8215 : BUF_X1 port map( A => n12335, Z => n11931);
   U8216 : BUF_X1 port map( A => n12335, Z => n11930);
   U8217 : BUF_X1 port map( A => n12339, Z => n11934);
   U8218 : BUF_X1 port map( A => n12339, Z => n11933);
   U8219 : BUF_X1 port map( A => n12343, Z => n11937);
   U8220 : BUF_X1 port map( A => n12343, Z => n11936);
   U8221 : BUF_X1 port map( A => n12347, Z => n11940);
   U8222 : BUF_X1 port map( A => n12347, Z => n11939);
   U8223 : BUF_X1 port map( A => n12351, Z => n11943);
   U8224 : BUF_X1 port map( A => n12351, Z => n11942);
   U8225 : BUF_X1 port map( A => n12355, Z => n11946);
   U8226 : BUF_X1 port map( A => n12355, Z => n11945);
   U8227 : BUF_X1 port map( A => n12359, Z => n11949);
   U8228 : BUF_X1 port map( A => n12359, Z => n11948);
   U8229 : BUF_X1 port map( A => n12363, Z => n11952);
   U8230 : BUF_X1 port map( A => n12363, Z => n11951);
   U8231 : BUF_X1 port map( A => n12367, Z => n11955);
   U8232 : BUF_X1 port map( A => n12367, Z => n11954);
   U8233 : BUF_X1 port map( A => n12371, Z => n11958);
   U8234 : BUF_X1 port map( A => n12371, Z => n11957);
   U8235 : BUF_X1 port map( A => n12375, Z => n11961);
   U8236 : BUF_X1 port map( A => n12375, Z => n11960);
   U8237 : BUF_X1 port map( A => n12379, Z => n11964);
   U8238 : BUF_X1 port map( A => n12379, Z => n11963);
   U8239 : BUF_X1 port map( A => n12383, Z => n11967);
   U8240 : BUF_X1 port map( A => n12383, Z => n11966);
   U8241 : INV_X1 port map( A => n12262, ZN => n12261);
   U8242 : INV_X1 port map( A => n12262, ZN => n12260);
   U8243 : INV_X1 port map( A => n12266, ZN => n12265);
   U8244 : INV_X1 port map( A => n12270, ZN => n12269);
   U8245 : INV_X1 port map( A => n12274, ZN => n12273);
   U8246 : INV_X1 port map( A => n12278, ZN => n12277);
   U8247 : INV_X1 port map( A => n12282, ZN => n12281);
   U8248 : INV_X1 port map( A => n12286, ZN => n12285);
   U8249 : INV_X1 port map( A => n12290, ZN => n12289);
   U8250 : INV_X1 port map( A => n12294, ZN => n12293);
   U8251 : INV_X1 port map( A => n12298, ZN => n12297);
   U8252 : INV_X1 port map( A => n12302, ZN => n12301);
   U8253 : INV_X1 port map( A => n12306, ZN => n12305);
   U8254 : INV_X1 port map( A => n12310, ZN => n12309);
   U8255 : INV_X1 port map( A => n12314, ZN => n12313);
   U8256 : INV_X1 port map( A => n12318, ZN => n12317);
   U8257 : INV_X1 port map( A => n12326, ZN => n12325);
   U8258 : INV_X1 port map( A => n12330, ZN => n12329);
   U8259 : INV_X1 port map( A => n12334, ZN => n12333);
   U8260 : INV_X1 port map( A => n12338, ZN => n12337);
   U8261 : INV_X1 port map( A => n12342, ZN => n12341);
   U8262 : INV_X1 port map( A => n12346, ZN => n12345);
   U8263 : INV_X1 port map( A => n12350, ZN => n12349);
   U8264 : INV_X1 port map( A => n12354, ZN => n12353);
   U8265 : INV_X1 port map( A => n12358, ZN => n12357);
   U8266 : INV_X1 port map( A => n12362, ZN => n12361);
   U8267 : INV_X1 port map( A => n12366, ZN => n12365);
   U8268 : INV_X1 port map( A => n12370, ZN => n12369);
   U8269 : INV_X1 port map( A => n12374, ZN => n12373);
   U8270 : INV_X1 port map( A => n12378, ZN => n12377);
   U8271 : INV_X1 port map( A => n12382, ZN => n12381);
   U8272 : BUF_X1 port map( A => n12263, Z => n11878);
   U8273 : BUF_X1 port map( A => n12267, Z => n11881);
   U8274 : BUF_X1 port map( A => n12271, Z => n11884);
   U8275 : BUF_X1 port map( A => n12275, Z => n11887);
   U8276 : BUF_X1 port map( A => n12279, Z => n11890);
   U8277 : BUF_X1 port map( A => n12283, Z => n11893);
   U8278 : BUF_X1 port map( A => n12287, Z => n11896);
   U8279 : BUF_X1 port map( A => n12291, Z => n11899);
   U8280 : BUF_X1 port map( A => n12295, Z => n11902);
   U8281 : BUF_X1 port map( A => n12299, Z => n11905);
   U8282 : BUF_X1 port map( A => n12303, Z => n11908);
   U8283 : BUF_X1 port map( A => n12307, Z => n11911);
   U8284 : BUF_X1 port map( A => n12311, Z => n11914);
   U8285 : BUF_X1 port map( A => n12315, Z => n11917);
   U8286 : BUF_X1 port map( A => n12319, Z => n11920);
   U8287 : BUF_X1 port map( A => n12327, Z => n11926);
   U8288 : BUF_X1 port map( A => n12331, Z => n11929);
   U8289 : BUF_X1 port map( A => n12335, Z => n11932);
   U8290 : BUF_X1 port map( A => n12339, Z => n11935);
   U8291 : BUF_X1 port map( A => n12343, Z => n11938);
   U8292 : BUF_X1 port map( A => n12347, Z => n11941);
   U8293 : BUF_X1 port map( A => n12351, Z => n11944);
   U8294 : BUF_X1 port map( A => n12355, Z => n11947);
   U8295 : BUF_X1 port map( A => n12359, Z => n11950);
   U8296 : BUF_X1 port map( A => n12363, Z => n11953);
   U8297 : BUF_X1 port map( A => n12367, Z => n11956);
   U8298 : BUF_X1 port map( A => n12371, Z => n11959);
   U8299 : BUF_X1 port map( A => n12375, Z => n11962);
   U8300 : BUF_X1 port map( A => n12379, Z => n11965);
   U8301 : BUF_X1 port map( A => n12383, Z => n11968);
   U8302 : INV_X1 port map( A => n9879, ZN => n12324);
   U8303 : OAI21_X1 port map( B1 => n9856, B2 => n9880, A => n12521, ZN => 
                           n9879);
   U8304 : INV_X1 port map( A => n9823, ZN => n12512);
   U8305 : OAI21_X1 port map( B1 => n9855, B2 => n9856, A => n12519, ZN => 
                           n9823);
   U8306 : BUF_X1 port map( A => n12523, Z => n12520);
   U8307 : BUF_X1 port map( A => n12523, Z => n12521);
   U8308 : BUF_X1 port map( A => n12058, Z => n11870);
   U8309 : BUF_X1 port map( A => n12202, Z => n11873);
   U8310 : BUF_X1 port map( A => n12524, Z => n12518);
   U8311 : BUF_X1 port map( A => n12524, Z => n12517);
   U8312 : BUF_X1 port map( A => n12058, Z => n11871);
   U8313 : BUF_X1 port map( A => n12202, Z => n11874);
   U8314 : BUF_X1 port map( A => n12087, Z => n12084);
   U8315 : BUF_X1 port map( A => n12071, Z => n12068);
   U8316 : BUF_X1 port map( A => n12087, Z => n12085);
   U8317 : BUF_X1 port map( A => n12071, Z => n12069);
   U8318 : BUF_X1 port map( A => n12231, Z => n12228);
   U8319 : BUF_X1 port map( A => n12215, Z => n12212);
   U8320 : BUF_X1 port map( A => n12231, Z => n12229);
   U8321 : BUF_X1 port map( A => n12215, Z => n12213);
   U8322 : BUF_X1 port map( A => n12524, Z => n12519);
   U8323 : BUF_X1 port map( A => n12051, Z => n12048);
   U8324 : BUF_X1 port map( A => n12083, Z => n12080);
   U8325 : BUF_X1 port map( A => n12067, Z => n12064);
   U8326 : BUF_X1 port map( A => n12051, Z => n12049);
   U8327 : BUF_X1 port map( A => n12083, Z => n12081);
   U8328 : BUF_X1 port map( A => n12067, Z => n12065);
   U8329 : BUF_X1 port map( A => n12195, Z => n12192);
   U8330 : BUF_X1 port map( A => n12227, Z => n12224);
   U8331 : BUF_X1 port map( A => n12211, Z => n12208);
   U8332 : BUF_X1 port map( A => n12195, Z => n12193);
   U8333 : BUF_X1 port map( A => n12227, Z => n12225);
   U8334 : BUF_X1 port map( A => n12211, Z => n12209);
   U8335 : BUF_X1 port map( A => n12112, Z => n12113);
   U8336 : BUF_X1 port map( A => n12092, Z => n12093);
   U8337 : BUF_X1 port map( A => n12076, Z => n12077);
   U8338 : BUF_X1 port map( A => n12112, Z => n12114);
   U8339 : BUF_X1 port map( A => n12092, Z => n12094);
   U8340 : BUF_X1 port map( A => n12076, Z => n12078);
   U8341 : BUF_X1 port map( A => n12256, Z => n12257);
   U8342 : BUF_X1 port map( A => n12236, Z => n12237);
   U8343 : BUF_X1 port map( A => n12220, Z => n12221);
   U8344 : BUF_X1 port map( A => n12256, Z => n12258);
   U8345 : BUF_X1 port map( A => n12236, Z => n12238);
   U8346 : BUF_X1 port map( A => n12220, Z => n12222);
   U8347 : BUF_X1 port map( A => n12063, Z => n12061);
   U8348 : BUF_X1 port map( A => n12063, Z => n12060);
   U8349 : BUF_X1 port map( A => n12207, Z => n12205);
   U8350 : BUF_X1 port map( A => n12207, Z => n12204);
   U8351 : BUF_X1 port map( A => n12024, Z => n12025);
   U8352 : BUF_X1 port map( A => n11988, Z => n11989);
   U8353 : BUF_X1 port map( A => n12040, Z => n12041);
   U8354 : BUF_X1 port map( A => n12004, Z => n12005);
   U8355 : BUF_X1 port map( A => n12024, Z => n12026);
   U8356 : BUF_X1 port map( A => n11988, Z => n11990);
   U8357 : BUF_X1 port map( A => n12040, Z => n12042);
   U8358 : BUF_X1 port map( A => n12004, Z => n12006);
   U8359 : BUF_X1 port map( A => n12168, Z => n12169);
   U8360 : BUF_X1 port map( A => n12132, Z => n12133);
   U8361 : BUF_X1 port map( A => n12184, Z => n12185);
   U8362 : BUF_X1 port map( A => n12148, Z => n12149);
   U8363 : BUF_X1 port map( A => n12168, Z => n12170);
   U8364 : BUF_X1 port map( A => n12132, Z => n12134);
   U8365 : BUF_X1 port map( A => n12184, Z => n12186);
   U8366 : BUF_X1 port map( A => n12148, Z => n12150);
   U8367 : BUF_X1 port map( A => n12020, Z => n12021);
   U8368 : BUF_X1 port map( A => n11984, Z => n11985);
   U8369 : BUF_X1 port map( A => n12020, Z => n12022);
   U8370 : BUF_X1 port map( A => n11984, Z => n11986);
   U8371 : BUF_X1 port map( A => n12164, Z => n12165);
   U8372 : BUF_X1 port map( A => n12128, Z => n12129);
   U8373 : BUF_X1 port map( A => n12164, Z => n12166);
   U8374 : BUF_X1 port map( A => n12128, Z => n12130);
   U8375 : BUF_X1 port map( A => n12036, Z => n12037);
   U8376 : BUF_X1 port map( A => n12000, Z => n12001);
   U8377 : BUF_X1 port map( A => n12036, Z => n12038);
   U8378 : BUF_X1 port map( A => n12000, Z => n12002);
   U8379 : BUF_X1 port map( A => n12180, Z => n12181);
   U8380 : BUF_X1 port map( A => n12144, Z => n12145);
   U8381 : BUF_X1 port map( A => n12180, Z => n12182);
   U8382 : BUF_X1 port map( A => n12144, Z => n12146);
   U8383 : BUF_X1 port map( A => n12108, Z => n12109);
   U8384 : BUF_X1 port map( A => n12088, Z => n12089);
   U8385 : BUF_X1 port map( A => n12072, Z => n12073);
   U8386 : BUF_X1 port map( A => n12108, Z => n12110);
   U8387 : BUF_X1 port map( A => n12088, Z => n12090);
   U8388 : BUF_X1 port map( A => n12072, Z => n12074);
   U8389 : BUF_X1 port map( A => n12252, Z => n12253);
   U8390 : BUF_X1 port map( A => n12232, Z => n12233);
   U8391 : BUF_X1 port map( A => n12216, Z => n12217);
   U8392 : BUF_X1 port map( A => n12252, Z => n12254);
   U8393 : BUF_X1 port map( A => n12232, Z => n12234);
   U8394 : BUF_X1 port map( A => n12216, Z => n12218);
   U8395 : BUF_X1 port map( A => n12028, Z => n12029);
   U8396 : BUF_X1 port map( A => n11992, Z => n11993);
   U8397 : BUF_X1 port map( A => n12044, Z => n12045);
   U8398 : BUF_X1 port map( A => n12008, Z => n12009);
   U8399 : BUF_X1 port map( A => n12028, Z => n12030);
   U8400 : BUF_X1 port map( A => n11992, Z => n11994);
   U8401 : BUF_X1 port map( A => n12044, Z => n12046);
   U8402 : BUF_X1 port map( A => n12008, Z => n12010);
   U8403 : BUF_X1 port map( A => n12172, Z => n12173);
   U8404 : BUF_X1 port map( A => n12136, Z => n12137);
   U8405 : BUF_X1 port map( A => n12188, Z => n12189);
   U8406 : BUF_X1 port map( A => n12152, Z => n12153);
   U8407 : BUF_X1 port map( A => n12172, Z => n12174);
   U8408 : BUF_X1 port map( A => n12136, Z => n12138);
   U8409 : BUF_X1 port map( A => n12188, Z => n12190);
   U8410 : BUF_X1 port map( A => n12152, Z => n12154);
   U8411 : BUF_X1 port map( A => n12099, Z => n12096);
   U8412 : BUF_X1 port map( A => n12099, Z => n12097);
   U8413 : BUF_X1 port map( A => n12243, Z => n12240);
   U8414 : BUF_X1 port map( A => n12243, Z => n12241);
   U8415 : INV_X1 port map( A => n12057, ZN => n12056);
   U8416 : INV_X1 port map( A => n12201, ZN => n12200);
   U8417 : BUF_X1 port map( A => n12019, Z => n12017);
   U8418 : BUF_X1 port map( A => n11983, Z => n11981);
   U8419 : BUF_X1 port map( A => n12019, Z => n12016);
   U8420 : BUF_X1 port map( A => n11983, Z => n11980);
   U8421 : BUF_X1 port map( A => n12163, Z => n12161);
   U8422 : BUF_X1 port map( A => n12127, Z => n12125);
   U8423 : BUF_X1 port map( A => n12163, Z => n12160);
   U8424 : BUF_X1 port map( A => n12127, Z => n12124);
   U8425 : BUF_X1 port map( A => n12103, Z => n12100);
   U8426 : BUF_X1 port map( A => n12103, Z => n12101);
   U8427 : BUF_X1 port map( A => n12247, Z => n12244);
   U8428 : BUF_X1 port map( A => n12247, Z => n12245);
   U8429 : INV_X1 port map( A => n12054, ZN => n12052);
   U8430 : INV_X1 port map( A => n12054, ZN => n12053);
   U8431 : INV_X1 port map( A => n12198, ZN => n12196);
   U8432 : INV_X1 port map( A => n12198, ZN => n12197);
   U8433 : BUF_X1 port map( A => n12107, Z => n12104);
   U8434 : BUF_X1 port map( A => n12107, Z => n12105);
   U8435 : BUF_X1 port map( A => n12251, Z => n12248);
   U8436 : BUF_X1 port map( A => n12251, Z => n12249);
   U8437 : BUF_X1 port map( A => n12035, Z => n12033);
   U8438 : BUF_X1 port map( A => n11999, Z => n11997);
   U8439 : BUF_X1 port map( A => n12035, Z => n12032);
   U8440 : BUF_X1 port map( A => n11999, Z => n11996);
   U8441 : BUF_X1 port map( A => n12179, Z => n12177);
   U8442 : BUF_X1 port map( A => n12143, Z => n12141);
   U8443 : BUF_X1 port map( A => n12179, Z => n12176);
   U8444 : BUF_X1 port map( A => n12143, Z => n12140);
   U8445 : BUF_X1 port map( A => n12015, Z => n12013);
   U8446 : BUF_X1 port map( A => n11979, Z => n11977);
   U8447 : BUF_X1 port map( A => n12015, Z => n12012);
   U8448 : BUF_X1 port map( A => n11979, Z => n11976);
   U8449 : BUF_X1 port map( A => n12159, Z => n12157);
   U8450 : BUF_X1 port map( A => n12123, Z => n12121);
   U8451 : BUF_X1 port map( A => n12159, Z => n12156);
   U8452 : BUF_X1 port map( A => n12123, Z => n12120);
   U8453 : BUF_X1 port map( A => n12087, Z => n12086);
   U8454 : BUF_X1 port map( A => n12071, Z => n12070);
   U8455 : BUF_X1 port map( A => n12231, Z => n12230);
   U8456 : BUF_X1 port map( A => n12215, Z => n12214);
   U8457 : BUF_X1 port map( A => n12051, Z => n12050);
   U8458 : BUF_X1 port map( A => n12083, Z => n12082);
   U8459 : BUF_X1 port map( A => n12067, Z => n12066);
   U8460 : BUF_X1 port map( A => n12195, Z => n12194);
   U8461 : BUF_X1 port map( A => n12227, Z => n12226);
   U8462 : BUF_X1 port map( A => n12211, Z => n12210);
   U8463 : BUF_X1 port map( A => n12112, Z => n12115);
   U8464 : BUF_X1 port map( A => n12092, Z => n12095);
   U8465 : BUF_X1 port map( A => n12076, Z => n12079);
   U8466 : BUF_X1 port map( A => n12256, Z => n12259);
   U8467 : BUF_X1 port map( A => n12236, Z => n12239);
   U8468 : BUF_X1 port map( A => n12220, Z => n12223);
   U8469 : BUF_X1 port map( A => n12063, Z => n12062);
   U8470 : BUF_X1 port map( A => n12207, Z => n12206);
   U8471 : BUF_X1 port map( A => n12024, Z => n12027);
   U8472 : BUF_X1 port map( A => n11988, Z => n11991);
   U8473 : BUF_X1 port map( A => n12040, Z => n12043);
   U8474 : BUF_X1 port map( A => n12004, Z => n12007);
   U8475 : BUF_X1 port map( A => n12168, Z => n12171);
   U8476 : BUF_X1 port map( A => n12132, Z => n12135);
   U8477 : BUF_X1 port map( A => n12184, Z => n12187);
   U8478 : BUF_X1 port map( A => n12148, Z => n12151);
   U8479 : BUF_X1 port map( A => n12020, Z => n12023);
   U8480 : BUF_X1 port map( A => n11984, Z => n11987);
   U8481 : BUF_X1 port map( A => n12164, Z => n12167);
   U8482 : BUF_X1 port map( A => n12128, Z => n12131);
   U8483 : BUF_X1 port map( A => n12036, Z => n12039);
   U8484 : BUF_X1 port map( A => n12000, Z => n12003);
   U8485 : BUF_X1 port map( A => n12180, Z => n12183);
   U8486 : BUF_X1 port map( A => n12144, Z => n12147);
   U8487 : BUF_X1 port map( A => n12108, Z => n12111);
   U8488 : BUF_X1 port map( A => n12088, Z => n12091);
   U8489 : BUF_X1 port map( A => n12072, Z => n12075);
   U8490 : BUF_X1 port map( A => n12252, Z => n12255);
   U8491 : BUF_X1 port map( A => n12232, Z => n12235);
   U8492 : BUF_X1 port map( A => n12216, Z => n12219);
   U8493 : BUF_X1 port map( A => n12028, Z => n12031);
   U8494 : BUF_X1 port map( A => n11992, Z => n11995);
   U8495 : BUF_X1 port map( A => n12044, Z => n12047);
   U8496 : BUF_X1 port map( A => n12008, Z => n12011);
   U8497 : BUF_X1 port map( A => n12172, Z => n12175);
   U8498 : BUF_X1 port map( A => n12136, Z => n12139);
   U8499 : BUF_X1 port map( A => n12188, Z => n12191);
   U8500 : BUF_X1 port map( A => n12152, Z => n12155);
   U8501 : BUF_X1 port map( A => n12099, Z => n12098);
   U8502 : BUF_X1 port map( A => n12243, Z => n12242);
   U8503 : BUF_X1 port map( A => n12019, Z => n12018);
   U8504 : BUF_X1 port map( A => n11983, Z => n11982);
   U8505 : BUF_X1 port map( A => n12163, Z => n12162);
   U8506 : BUF_X1 port map( A => n12127, Z => n12126);
   U8507 : BUF_X1 port map( A => n12103, Z => n12102);
   U8508 : BUF_X1 port map( A => n12247, Z => n12246);
   U8509 : BUF_X1 port map( A => n12107, Z => n12106);
   U8510 : BUF_X1 port map( A => n12251, Z => n12250);
   U8511 : BUF_X1 port map( A => n12035, Z => n12034);
   U8512 : BUF_X1 port map( A => n11999, Z => n11998);
   U8513 : BUF_X1 port map( A => n12179, Z => n12178);
   U8514 : BUF_X1 port map( A => n12143, Z => n12142);
   U8515 : BUF_X1 port map( A => n12015, Z => n12014);
   U8516 : BUF_X1 port map( A => n11979, Z => n11978);
   U8517 : BUF_X1 port map( A => n12159, Z => n12158);
   U8518 : BUF_X1 port map( A => n12123, Z => n12122);
   U8519 : BUF_X1 port map( A => n12058, Z => n11872);
   U8520 : BUF_X1 port map( A => n12202, Z => n11875);
   U8521 : BUF_X1 port map( A => n12523, Z => n12522);
   U8522 : OAI222_X1 port map( A1 => n9341, A2 => n12104, B1 => n9533, B2 => 
                           n12100, C1 => n9469, C2 => n12096, ZN => n11067);
   U8523 : OAI222_X1 port map( A1 => n9340, A2 => n12104, B1 => n9532, B2 => 
                           n12100, C1 => n9468, C2 => n12096, ZN => n11050);
   U8524 : OAI222_X1 port map( A1 => n9339, A2 => n12104, B1 => n9531, B2 => 
                           n12100, C1 => n9467, C2 => n12096, ZN => n11033);
   U8525 : OAI222_X1 port map( A1 => n9338, A2 => n12104, B1 => n9530, B2 => 
                           n12100, C1 => n9466, C2 => n12096, ZN => n11016);
   U8526 : OAI222_X1 port map( A1 => n9337, A2 => n12104, B1 => n9529, B2 => 
                           n12100, C1 => n9465, C2 => n12096, ZN => n10999);
   U8527 : OAI222_X1 port map( A1 => n9336, A2 => n12104, B1 => n9528, B2 => 
                           n12100, C1 => n9464, C2 => n12096, ZN => n10982);
   U8528 : OAI222_X1 port map( A1 => n9335, A2 => n12104, B1 => n9527, B2 => 
                           n12100, C1 => n9463, C2 => n12096, ZN => n10965);
   U8529 : OAI222_X1 port map( A1 => n9334, A2 => n12104, B1 => n9526, B2 => 
                           n12100, C1 => n9462, C2 => n12096, ZN => n10948);
   U8530 : OAI222_X1 port map( A1 => n9333, A2 => n12104, B1 => n9525, B2 => 
                           n12100, C1 => n9461, C2 => n12096, ZN => n10931);
   U8531 : OAI222_X1 port map( A1 => n9332, A2 => n12104, B1 => n9524, B2 => 
                           n12100, C1 => n9460, C2 => n12096, ZN => n10914);
   U8532 : OAI222_X1 port map( A1 => n9331, A2 => n12104, B1 => n9523, B2 => 
                           n12100, C1 => n9459, C2 => n12096, ZN => n10897);
   U8533 : OAI222_X1 port map( A1 => n9330, A2 => n12104, B1 => n9522, B2 => 
                           n12100, C1 => n9458, C2 => n12096, ZN => n10880);
   U8534 : OAI222_X1 port map( A1 => n9329, A2 => n12105, B1 => n9521, B2 => 
                           n12101, C1 => n9457, C2 => n12097, ZN => n10863);
   U8535 : OAI222_X1 port map( A1 => n9328, A2 => n12105, B1 => n9520, B2 => 
                           n12101, C1 => n9456, C2 => n12097, ZN => n10846);
   U8536 : OAI222_X1 port map( A1 => n9327, A2 => n12105, B1 => n9519, B2 => 
                           n12101, C1 => n9455, C2 => n12097, ZN => n10829);
   U8537 : OAI222_X1 port map( A1 => n9326, A2 => n12105, B1 => n9518, B2 => 
                           n12101, C1 => n9454, C2 => n12097, ZN => n10812);
   U8538 : OAI222_X1 port map( A1 => n9325, A2 => n12105, B1 => n9517, B2 => 
                           n12101, C1 => n9453, C2 => n12097, ZN => n10795);
   U8539 : OAI222_X1 port map( A1 => n9324, A2 => n12105, B1 => n9516, B2 => 
                           n12101, C1 => n9452, C2 => n12097, ZN => n10778);
   U8540 : OAI222_X1 port map( A1 => n9323, A2 => n12105, B1 => n9515, B2 => 
                           n12101, C1 => n9451, C2 => n12097, ZN => n10761);
   U8541 : OAI222_X1 port map( A1 => n9322, A2 => n12105, B1 => n9514, B2 => 
                           n12101, C1 => n9450, C2 => n12097, ZN => n10744);
   U8542 : OAI222_X1 port map( A1 => n9321, A2 => n12105, B1 => n9513, B2 => 
                           n12101, C1 => n9449, C2 => n12097, ZN => n10727);
   U8543 : OAI222_X1 port map( A1 => n9320, A2 => n12105, B1 => n9512, B2 => 
                           n12101, C1 => n9448, C2 => n12097, ZN => n10710);
   U8544 : OAI222_X1 port map( A1 => n9319, A2 => n12105, B1 => n9511, B2 => 
                           n12101, C1 => n9447, C2 => n12097, ZN => n10693);
   U8545 : OAI222_X1 port map( A1 => n9318, A2 => n12105, B1 => n9510, B2 => 
                           n12101, C1 => n9446, C2 => n12097, ZN => n10676);
   U8546 : OAI222_X1 port map( A1 => n9317, A2 => n12106, B1 => n9509, B2 => 
                           n12102, C1 => n9445, C2 => n12098, ZN => n10659);
   U8547 : OAI222_X1 port map( A1 => n9316, A2 => n12106, B1 => n9508, B2 => 
                           n12102, C1 => n9444, C2 => n12098, ZN => n10642);
   U8548 : OAI222_X1 port map( A1 => n9315, A2 => n12106, B1 => n9507, B2 => 
                           n12102, C1 => n9443, C2 => n12098, ZN => n10625);
   U8549 : OAI222_X1 port map( A1 => n9314, A2 => n12106, B1 => n9506, B2 => 
                           n12102, C1 => n9442, C2 => n12098, ZN => n10608);
   U8550 : OAI222_X1 port map( A1 => n9313, A2 => n12106, B1 => n9505, B2 => 
                           n12102, C1 => n9441, C2 => n12098, ZN => n10591);
   U8551 : OAI222_X1 port map( A1 => n9312, A2 => n12106, B1 => n9504, B2 => 
                           n12102, C1 => n9440, C2 => n12098, ZN => n10574);
   U8552 : OAI222_X1 port map( A1 => n9311, A2 => n12106, B1 => n9503, B2 => 
                           n12102, C1 => n9439, C2 => n12098, ZN => n10557);
   U8553 : OAI222_X1 port map( A1 => n9310, A2 => n12106, B1 => n9502, B2 => 
                           n12102, C1 => n9438, C2 => n12098, ZN => n10506);
   U8554 : OAI222_X1 port map( A1 => n9341, A2 => n12248, B1 => n9533, B2 => 
                           n12244, C1 => n9469, C2 => n12240, ZN => n10467);
   U8555 : OAI222_X1 port map( A1 => n9340, A2 => n12248, B1 => n9532, B2 => 
                           n12244, C1 => n9468, C2 => n12240, ZN => n10450);
   U8556 : OAI222_X1 port map( A1 => n9339, A2 => n12248, B1 => n9531, B2 => 
                           n12244, C1 => n9467, C2 => n12240, ZN => n10433);
   U8557 : OAI222_X1 port map( A1 => n9338, A2 => n12248, B1 => n9530, B2 => 
                           n12244, C1 => n9466, C2 => n12240, ZN => n10416);
   U8558 : OAI222_X1 port map( A1 => n9337, A2 => n12248, B1 => n9529, B2 => 
                           n12244, C1 => n9465, C2 => n12240, ZN => n10399);
   U8559 : OAI222_X1 port map( A1 => n9336, A2 => n12248, B1 => n9528, B2 => 
                           n12244, C1 => n9464, C2 => n12240, ZN => n10382);
   U8560 : OAI222_X1 port map( A1 => n9335, A2 => n12248, B1 => n9527, B2 => 
                           n12244, C1 => n9463, C2 => n12240, ZN => n10365);
   U8561 : OAI222_X1 port map( A1 => n9334, A2 => n12248, B1 => n9526, B2 => 
                           n12244, C1 => n9462, C2 => n12240, ZN => n10348);
   U8562 : OAI222_X1 port map( A1 => n9333, A2 => n12248, B1 => n9525, B2 => 
                           n12244, C1 => n9461, C2 => n12240, ZN => n10331);
   U8563 : OAI222_X1 port map( A1 => n9332, A2 => n12248, B1 => n9524, B2 => 
                           n12244, C1 => n9460, C2 => n12240, ZN => n10314);
   U8564 : OAI222_X1 port map( A1 => n9331, A2 => n12248, B1 => n9523, B2 => 
                           n12244, C1 => n9459, C2 => n12240, ZN => n10297);
   U8565 : OAI222_X1 port map( A1 => n9330, A2 => n12248, B1 => n9522, B2 => 
                           n12244, C1 => n9458, C2 => n12240, ZN => n10280);
   U8566 : OAI222_X1 port map( A1 => n9329, A2 => n12249, B1 => n9521, B2 => 
                           n12245, C1 => n9457, C2 => n12241, ZN => n10263);
   U8567 : OAI222_X1 port map( A1 => n9328, A2 => n12249, B1 => n9520, B2 => 
                           n12245, C1 => n9456, C2 => n12241, ZN => n10246);
   U8568 : OAI222_X1 port map( A1 => n9327, A2 => n12249, B1 => n9519, B2 => 
                           n12245, C1 => n9455, C2 => n12241, ZN => n10229);
   U8569 : OAI222_X1 port map( A1 => n9326, A2 => n12249, B1 => n9518, B2 => 
                           n12245, C1 => n9454, C2 => n12241, ZN => n10212);
   U8570 : OAI222_X1 port map( A1 => n9325, A2 => n12249, B1 => n9517, B2 => 
                           n12245, C1 => n9453, C2 => n12241, ZN => n10195);
   U8571 : OAI222_X1 port map( A1 => n9324, A2 => n12249, B1 => n9516, B2 => 
                           n12245, C1 => n9452, C2 => n12241, ZN => n10178);
   U8572 : OAI222_X1 port map( A1 => n9323, A2 => n12249, B1 => n9515, B2 => 
                           n12245, C1 => n9451, C2 => n12241, ZN => n10161);
   U8573 : OAI222_X1 port map( A1 => n9322, A2 => n12249, B1 => n9514, B2 => 
                           n12245, C1 => n9450, C2 => n12241, ZN => n10144);
   U8574 : OAI222_X1 port map( A1 => n9321, A2 => n12249, B1 => n9513, B2 => 
                           n12245, C1 => n9449, C2 => n12241, ZN => n10127);
   U8575 : OAI222_X1 port map( A1 => n9320, A2 => n12249, B1 => n9512, B2 => 
                           n12245, C1 => n9448, C2 => n12241, ZN => n10110);
   U8576 : OAI222_X1 port map( A1 => n9319, A2 => n12249, B1 => n9511, B2 => 
                           n12245, C1 => n9447, C2 => n12241, ZN => n10093);
   U8577 : OAI222_X1 port map( A1 => n9318, A2 => n12249, B1 => n9510, B2 => 
                           n12245, C1 => n9446, C2 => n12241, ZN => n10076);
   U8578 : OAI222_X1 port map( A1 => n9317, A2 => n12250, B1 => n9509, B2 => 
                           n12246, C1 => n9445, C2 => n12242, ZN => n10059);
   U8579 : OAI222_X1 port map( A1 => n9316, A2 => n12250, B1 => n9508, B2 => 
                           n12246, C1 => n9444, C2 => n12242, ZN => n10042);
   U8580 : OAI222_X1 port map( A1 => n9315, A2 => n12250, B1 => n9507, B2 => 
                           n12246, C1 => n9443, C2 => n12242, ZN => n10025);
   U8581 : OAI222_X1 port map( A1 => n9314, A2 => n12250, B1 => n9506, B2 => 
                           n12246, C1 => n9442, C2 => n12242, ZN => n10008);
   U8582 : OAI222_X1 port map( A1 => n9313, A2 => n12250, B1 => n9505, B2 => 
                           n12246, C1 => n9441, C2 => n12242, ZN => n9991);
   U8583 : OAI222_X1 port map( A1 => n9312, A2 => n12250, B1 => n9504, B2 => 
                           n12246, C1 => n9440, C2 => n12242, ZN => n9974);
   U8584 : OAI222_X1 port map( A1 => n9311, A2 => n12250, B1 => n9503, B2 => 
                           n12246, C1 => n9439, C2 => n12242, ZN => n9957);
   U8585 : OAI222_X1 port map( A1 => n9310, A2 => n12250, B1 => n9502, B2 => 
                           n12246, C1 => n9438, C2 => n12242, ZN => n9906);
   U8586 : OAI22_X1 port map( A1 => n9757, A2 => n12084, B1 => n9405, B2 => 
                           n12080, ZN => n11074);
   U8587 : OAI22_X1 port map( A1 => n9756, A2 => n12084, B1 => n9404, B2 => 
                           n12080, ZN => n11051);
   U8588 : OAI22_X1 port map( A1 => n9755, A2 => n12084, B1 => n9403, B2 => 
                           n12080, ZN => n11034);
   U8589 : OAI22_X1 port map( A1 => n9754, A2 => n12084, B1 => n9402, B2 => 
                           n12080, ZN => n11017);
   U8590 : OAI22_X1 port map( A1 => n9753, A2 => n12084, B1 => n9401, B2 => 
                           n12080, ZN => n11000);
   U8591 : OAI22_X1 port map( A1 => n9752, A2 => n12084, B1 => n9400, B2 => 
                           n12080, ZN => n10983);
   U8592 : OAI22_X1 port map( A1 => n9751, A2 => n12084, B1 => n9399, B2 => 
                           n12080, ZN => n10966);
   U8593 : OAI22_X1 port map( A1 => n9750, A2 => n12084, B1 => n9398, B2 => 
                           n12080, ZN => n10949);
   U8594 : OAI22_X1 port map( A1 => n9749, A2 => n12084, B1 => n9397, B2 => 
                           n12080, ZN => n10932);
   U8595 : OAI22_X1 port map( A1 => n9748, A2 => n12084, B1 => n9396, B2 => 
                           n12080, ZN => n10915);
   U8596 : OAI22_X1 port map( A1 => n9747, A2 => n12084, B1 => n9395, B2 => 
                           n12080, ZN => n10898);
   U8597 : OAI22_X1 port map( A1 => n9746, A2 => n12084, B1 => n9394, B2 => 
                           n12080, ZN => n10881);
   U8598 : OAI22_X1 port map( A1 => n9745, A2 => n12085, B1 => n9393, B2 => 
                           n12081, ZN => n10864);
   U8599 : OAI22_X1 port map( A1 => n9744, A2 => n12085, B1 => n9392, B2 => 
                           n12081, ZN => n10847);
   U8600 : OAI22_X1 port map( A1 => n9743, A2 => n12085, B1 => n9391, B2 => 
                           n12081, ZN => n10830);
   U8601 : OAI22_X1 port map( A1 => n9742, A2 => n12085, B1 => n9390, B2 => 
                           n12081, ZN => n10813);
   U8602 : OAI22_X1 port map( A1 => n9741, A2 => n12085, B1 => n9389, B2 => 
                           n12081, ZN => n10796);
   U8603 : OAI22_X1 port map( A1 => n9740, A2 => n12085, B1 => n9388, B2 => 
                           n12081, ZN => n10779);
   U8604 : OAI22_X1 port map( A1 => n9739, A2 => n12085, B1 => n9387, B2 => 
                           n12081, ZN => n10762);
   U8605 : OAI22_X1 port map( A1 => n9738, A2 => n12085, B1 => n9386, B2 => 
                           n12081, ZN => n10745);
   U8606 : OAI22_X1 port map( A1 => n9737, A2 => n12085, B1 => n9385, B2 => 
                           n12081, ZN => n10728);
   U8607 : OAI22_X1 port map( A1 => n9736, A2 => n12085, B1 => n9384, B2 => 
                           n12081, ZN => n10711);
   U8608 : OAI22_X1 port map( A1 => n9735, A2 => n12085, B1 => n9383, B2 => 
                           n12081, ZN => n10694);
   U8609 : OAI22_X1 port map( A1 => n9734, A2 => n12085, B1 => n9382, B2 => 
                           n12081, ZN => n10677);
   U8610 : OAI22_X1 port map( A1 => n9733, A2 => n12086, B1 => n9381, B2 => 
                           n12082, ZN => n10660);
   U8611 : OAI22_X1 port map( A1 => n9732, A2 => n12086, B1 => n9380, B2 => 
                           n12082, ZN => n10643);
   U8612 : OAI22_X1 port map( A1 => n9731, A2 => n12086, B1 => n9379, B2 => 
                           n12082, ZN => n10626);
   U8613 : OAI22_X1 port map( A1 => n9730, A2 => n12086, B1 => n9378, B2 => 
                           n12082, ZN => n10609);
   U8614 : OAI22_X1 port map( A1 => n9729, A2 => n12086, B1 => n9377, B2 => 
                           n12082, ZN => n10592);
   U8615 : OAI22_X1 port map( A1 => n9728, A2 => n12086, B1 => n9376, B2 => 
                           n12082, ZN => n10575);
   U8616 : OAI22_X1 port map( A1 => n9727, A2 => n12086, B1 => n9375, B2 => 
                           n12082, ZN => n10558);
   U8617 : OAI22_X1 port map( A1 => n9726, A2 => n12086, B1 => n9374, B2 => 
                           n12082, ZN => n10512);
   U8618 : OAI22_X1 port map( A1 => n9757, A2 => n12228, B1 => n9405, B2 => 
                           n12224, ZN => n10474);
   U8619 : OAI22_X1 port map( A1 => n9756, A2 => n12228, B1 => n9404, B2 => 
                           n12224, ZN => n10451);
   U8620 : OAI22_X1 port map( A1 => n9755, A2 => n12228, B1 => n9403, B2 => 
                           n12224, ZN => n10434);
   U8621 : OAI22_X1 port map( A1 => n9754, A2 => n12228, B1 => n9402, B2 => 
                           n12224, ZN => n10417);
   U8622 : OAI22_X1 port map( A1 => n9753, A2 => n12228, B1 => n9401, B2 => 
                           n12224, ZN => n10400);
   U8623 : OAI22_X1 port map( A1 => n9752, A2 => n12228, B1 => n9400, B2 => 
                           n12224, ZN => n10383);
   U8624 : OAI22_X1 port map( A1 => n9751, A2 => n12228, B1 => n9399, B2 => 
                           n12224, ZN => n10366);
   U8625 : OAI22_X1 port map( A1 => n9750, A2 => n12228, B1 => n9398, B2 => 
                           n12224, ZN => n10349);
   U8626 : OAI22_X1 port map( A1 => n9749, A2 => n12228, B1 => n9397, B2 => 
                           n12224, ZN => n10332);
   U8627 : OAI22_X1 port map( A1 => n9748, A2 => n12228, B1 => n9396, B2 => 
                           n12224, ZN => n10315);
   U8628 : OAI22_X1 port map( A1 => n9747, A2 => n12228, B1 => n9395, B2 => 
                           n12224, ZN => n10298);
   U8629 : OAI22_X1 port map( A1 => n9746, A2 => n12228, B1 => n9394, B2 => 
                           n12224, ZN => n10281);
   U8630 : OAI22_X1 port map( A1 => n9745, A2 => n12229, B1 => n9393, B2 => 
                           n12225, ZN => n10264);
   U8631 : OAI22_X1 port map( A1 => n9744, A2 => n12229, B1 => n9392, B2 => 
                           n12225, ZN => n10247);
   U8632 : OAI22_X1 port map( A1 => n9743, A2 => n12229, B1 => n9391, B2 => 
                           n12225, ZN => n10230);
   U8633 : OAI22_X1 port map( A1 => n9742, A2 => n12229, B1 => n9390, B2 => 
                           n12225, ZN => n10213);
   U8634 : OAI22_X1 port map( A1 => n9741, A2 => n12229, B1 => n9389, B2 => 
                           n12225, ZN => n10196);
   U8635 : OAI22_X1 port map( A1 => n9740, A2 => n12229, B1 => n9388, B2 => 
                           n12225, ZN => n10179);
   U8636 : OAI22_X1 port map( A1 => n9739, A2 => n12229, B1 => n9387, B2 => 
                           n12225, ZN => n10162);
   U8637 : OAI22_X1 port map( A1 => n9738, A2 => n12229, B1 => n9386, B2 => 
                           n12225, ZN => n10145);
   U8638 : OAI22_X1 port map( A1 => n9737, A2 => n12229, B1 => n9385, B2 => 
                           n12225, ZN => n10128);
   U8639 : OAI22_X1 port map( A1 => n9736, A2 => n12229, B1 => n9384, B2 => 
                           n12225, ZN => n10111);
   U8640 : OAI22_X1 port map( A1 => n9735, A2 => n12229, B1 => n9383, B2 => 
                           n12225, ZN => n10094);
   U8641 : OAI22_X1 port map( A1 => n9734, A2 => n12229, B1 => n9382, B2 => 
                           n12225, ZN => n10077);
   U8642 : OAI22_X1 port map( A1 => n9733, A2 => n12230, B1 => n9381, B2 => 
                           n12226, ZN => n10060);
   U8643 : OAI22_X1 port map( A1 => n9732, A2 => n12230, B1 => n9380, B2 => 
                           n12226, ZN => n10043);
   U8644 : OAI22_X1 port map( A1 => n9731, A2 => n12230, B1 => n9379, B2 => 
                           n12226, ZN => n10026);
   U8645 : OAI22_X1 port map( A1 => n9730, A2 => n12230, B1 => n9378, B2 => 
                           n12226, ZN => n10009);
   U8646 : OAI22_X1 port map( A1 => n9729, A2 => n12230, B1 => n9377, B2 => 
                           n12226, ZN => n9992);
   U8647 : OAI22_X1 port map( A1 => n9728, A2 => n12230, B1 => n9376, B2 => 
                           n12226, ZN => n9975);
   U8648 : OAI22_X1 port map( A1 => n9727, A2 => n12230, B1 => n9375, B2 => 
                           n12226, ZN => n9958);
   U8649 : OAI22_X1 port map( A1 => n9726, A2 => n12230, B1 => n9374, B2 => 
                           n12226, ZN => n9912);
   U8650 : OAI22_X1 port map( A1 => n9661, A2 => n12068, B1 => n9597, B2 => 
                           n12064, ZN => n11079);
   U8651 : OAI22_X1 port map( A1 => n9660, A2 => n12068, B1 => n9596, B2 => 
                           n12064, ZN => n11052);
   U8652 : OAI22_X1 port map( A1 => n9659, A2 => n12068, B1 => n9595, B2 => 
                           n12064, ZN => n11035);
   U8653 : OAI22_X1 port map( A1 => n9658, A2 => n12068, B1 => n9594, B2 => 
                           n12064, ZN => n11018);
   U8654 : OAI22_X1 port map( A1 => n9657, A2 => n12068, B1 => n9593, B2 => 
                           n12064, ZN => n11001);
   U8655 : OAI22_X1 port map( A1 => n9656, A2 => n12068, B1 => n9592, B2 => 
                           n12064, ZN => n10984);
   U8656 : OAI22_X1 port map( A1 => n9655, A2 => n12068, B1 => n9591, B2 => 
                           n12064, ZN => n10967);
   U8657 : OAI22_X1 port map( A1 => n9654, A2 => n12068, B1 => n9590, B2 => 
                           n12064, ZN => n10950);
   U8658 : OAI22_X1 port map( A1 => n9653, A2 => n12068, B1 => n9589, B2 => 
                           n12064, ZN => n10933);
   U8659 : OAI22_X1 port map( A1 => n9652, A2 => n12068, B1 => n9588, B2 => 
                           n12064, ZN => n10916);
   U8660 : OAI22_X1 port map( A1 => n9651, A2 => n12068, B1 => n9587, B2 => 
                           n12064, ZN => n10899);
   U8661 : OAI22_X1 port map( A1 => n9650, A2 => n12068, B1 => n9586, B2 => 
                           n12064, ZN => n10882);
   U8662 : OAI22_X1 port map( A1 => n9649, A2 => n12069, B1 => n9585, B2 => 
                           n12065, ZN => n10865);
   U8663 : OAI22_X1 port map( A1 => n9648, A2 => n12069, B1 => n9584, B2 => 
                           n12065, ZN => n10848);
   U8664 : OAI22_X1 port map( A1 => n9647, A2 => n12069, B1 => n9583, B2 => 
                           n12065, ZN => n10831);
   U8665 : OAI22_X1 port map( A1 => n9646, A2 => n12069, B1 => n9582, B2 => 
                           n12065, ZN => n10814);
   U8666 : OAI22_X1 port map( A1 => n9645, A2 => n12069, B1 => n9581, B2 => 
                           n12065, ZN => n10797);
   U8667 : OAI22_X1 port map( A1 => n9644, A2 => n12069, B1 => n9580, B2 => 
                           n12065, ZN => n10780);
   U8668 : OAI22_X1 port map( A1 => n9643, A2 => n12069, B1 => n9579, B2 => 
                           n12065, ZN => n10763);
   U8669 : OAI22_X1 port map( A1 => n9642, A2 => n12069, B1 => n9578, B2 => 
                           n12065, ZN => n10746);
   U8670 : OAI22_X1 port map( A1 => n9641, A2 => n12069, B1 => n9577, B2 => 
                           n12065, ZN => n10729);
   U8671 : OAI22_X1 port map( A1 => n9640, A2 => n12069, B1 => n9576, B2 => 
                           n12065, ZN => n10712);
   U8672 : OAI22_X1 port map( A1 => n9639, A2 => n12069, B1 => n9575, B2 => 
                           n12065, ZN => n10695);
   U8673 : OAI22_X1 port map( A1 => n9638, A2 => n12069, B1 => n9574, B2 => 
                           n12065, ZN => n10678);
   U8674 : OAI22_X1 port map( A1 => n9637, A2 => n12070, B1 => n9573, B2 => 
                           n12066, ZN => n10661);
   U8675 : OAI22_X1 port map( A1 => n9636, A2 => n12070, B1 => n9572, B2 => 
                           n12066, ZN => n10644);
   U8676 : OAI22_X1 port map( A1 => n9635, A2 => n12070, B1 => n9571, B2 => 
                           n12066, ZN => n10627);
   U8677 : OAI22_X1 port map( A1 => n9634, A2 => n12070, B1 => n9570, B2 => 
                           n12066, ZN => n10610);
   U8678 : OAI22_X1 port map( A1 => n9633, A2 => n12070, B1 => n9569, B2 => 
                           n12066, ZN => n10593);
   U8679 : OAI22_X1 port map( A1 => n9632, A2 => n12070, B1 => n9568, B2 => 
                           n12066, ZN => n10576);
   U8680 : OAI22_X1 port map( A1 => n9631, A2 => n12070, B1 => n9567, B2 => 
                           n12066, ZN => n10559);
   U8681 : OAI22_X1 port map( A1 => n9630, A2 => n12070, B1 => n9566, B2 => 
                           n12066, ZN => n10517);
   U8682 : OAI22_X1 port map( A1 => n9661, A2 => n12212, B1 => n9597, B2 => 
                           n12208, ZN => n10479);
   U8683 : OAI22_X1 port map( A1 => n9660, A2 => n12212, B1 => n9596, B2 => 
                           n12208, ZN => n10452);
   U8684 : OAI22_X1 port map( A1 => n9659, A2 => n12212, B1 => n9595, B2 => 
                           n12208, ZN => n10435);
   U8685 : OAI22_X1 port map( A1 => n9658, A2 => n12212, B1 => n9594, B2 => 
                           n12208, ZN => n10418);
   U8686 : OAI22_X1 port map( A1 => n9657, A2 => n12212, B1 => n9593, B2 => 
                           n12208, ZN => n10401);
   U8687 : OAI22_X1 port map( A1 => n9656, A2 => n12212, B1 => n9592, B2 => 
                           n12208, ZN => n10384);
   U8688 : OAI22_X1 port map( A1 => n9655, A2 => n12212, B1 => n9591, B2 => 
                           n12208, ZN => n10367);
   U8689 : OAI22_X1 port map( A1 => n9654, A2 => n12212, B1 => n9590, B2 => 
                           n12208, ZN => n10350);
   U8690 : OAI22_X1 port map( A1 => n9653, A2 => n12212, B1 => n9589, B2 => 
                           n12208, ZN => n10333);
   U8691 : OAI22_X1 port map( A1 => n9652, A2 => n12212, B1 => n9588, B2 => 
                           n12208, ZN => n10316);
   U8692 : OAI22_X1 port map( A1 => n9651, A2 => n12212, B1 => n9587, B2 => 
                           n12208, ZN => n10299);
   U8693 : OAI22_X1 port map( A1 => n9650, A2 => n12212, B1 => n9586, B2 => 
                           n12208, ZN => n10282);
   U8694 : OAI22_X1 port map( A1 => n9649, A2 => n12213, B1 => n9585, B2 => 
                           n12209, ZN => n10265);
   U8695 : OAI22_X1 port map( A1 => n9648, A2 => n12213, B1 => n9584, B2 => 
                           n12209, ZN => n10248);
   U8696 : OAI22_X1 port map( A1 => n9647, A2 => n12213, B1 => n9583, B2 => 
                           n12209, ZN => n10231);
   U8697 : OAI22_X1 port map( A1 => n9646, A2 => n12213, B1 => n9582, B2 => 
                           n12209, ZN => n10214);
   U8698 : OAI22_X1 port map( A1 => n9645, A2 => n12213, B1 => n9581, B2 => 
                           n12209, ZN => n10197);
   U8699 : OAI22_X1 port map( A1 => n9644, A2 => n12213, B1 => n9580, B2 => 
                           n12209, ZN => n10180);
   U8700 : OAI22_X1 port map( A1 => n9643, A2 => n12213, B1 => n9579, B2 => 
                           n12209, ZN => n10163);
   U8701 : OAI22_X1 port map( A1 => n9642, A2 => n12213, B1 => n9578, B2 => 
                           n12209, ZN => n10146);
   U8702 : OAI22_X1 port map( A1 => n9641, A2 => n12213, B1 => n9577, B2 => 
                           n12209, ZN => n10129);
   U8703 : OAI22_X1 port map( A1 => n9640, A2 => n12213, B1 => n9576, B2 => 
                           n12209, ZN => n10112);
   U8704 : OAI22_X1 port map( A1 => n9639, A2 => n12213, B1 => n9575, B2 => 
                           n12209, ZN => n10095);
   U8705 : OAI22_X1 port map( A1 => n9638, A2 => n12213, B1 => n9574, B2 => 
                           n12209, ZN => n10078);
   U8706 : OAI22_X1 port map( A1 => n9637, A2 => n12214, B1 => n9573, B2 => 
                           n12210, ZN => n10061);
   U8707 : OAI22_X1 port map( A1 => n9636, A2 => n12214, B1 => n9572, B2 => 
                           n12210, ZN => n10044);
   U8708 : OAI22_X1 port map( A1 => n9635, A2 => n12214, B1 => n9571, B2 => 
                           n12210, ZN => n10027);
   U8709 : OAI22_X1 port map( A1 => n9634, A2 => n12214, B1 => n9570, B2 => 
                           n12210, ZN => n10010);
   U8710 : OAI22_X1 port map( A1 => n9633, A2 => n12214, B1 => n9569, B2 => 
                           n12210, ZN => n9993);
   U8711 : OAI22_X1 port map( A1 => n9632, A2 => n12214, B1 => n9568, B2 => 
                           n12210, ZN => n9976);
   U8712 : OAI22_X1 port map( A1 => n9631, A2 => n12214, B1 => n9567, B2 => 
                           n12210, ZN => n9959);
   U8713 : OAI22_X1 port map( A1 => n9630, A2 => n12214, B1 => n9566, B2 => 
                           n12210, ZN => n9917);
   U8714 : OAI22_X1 port map( A1 => n11926, A2 => n12387, B1 => n12325, B2 => 
                           n9309, ZN => n2123);
   U8715 : OAI22_X1 port map( A1 => n11926, A2 => n12391, B1 => n12325, B2 => 
                           n9308, ZN => n2124);
   U8716 : OAI22_X1 port map( A1 => n11926, A2 => n12395, B1 => n12325, B2 => 
                           n9307, ZN => n2125);
   U8717 : OAI22_X1 port map( A1 => n11926, A2 => n12399, B1 => n12325, B2 => 
                           n9306, ZN => n2126);
   U8718 : OAI22_X1 port map( A1 => n11926, A2 => n12403, B1 => n12325, B2 => 
                           n9305, ZN => n2127);
   U8719 : OAI22_X1 port map( A1 => n11926, A2 => n12407, B1 => n12325, B2 => 
                           n9304, ZN => n2128);
   U8720 : OAI22_X1 port map( A1 => n11926, A2 => n12411, B1 => n12325, B2 => 
                           n9303, ZN => n2129);
   U8721 : OAI22_X1 port map( A1 => n11926, A2 => n12415, B1 => n12325, B2 => 
                           n9302, ZN => n2130);
   U8722 : OAI22_X1 port map( A1 => n11925, A2 => n12419, B1 => n12325, B2 => 
                           n9301, ZN => n2131);
   U8723 : OAI22_X1 port map( A1 => n11925, A2 => n12423, B1 => n12325, B2 => 
                           n9300, ZN => n2132);
   U8724 : OAI22_X1 port map( A1 => n11925, A2 => n12427, B1 => n12325, B2 => 
                           n9299, ZN => n2133);
   U8725 : OAI22_X1 port map( A1 => n11925, A2 => n12431, B1 => n12325, B2 => 
                           n9298, ZN => n2134);
   U8726 : OAI22_X1 port map( A1 => n11925, A2 => n12435, B1 => n9878, B2 => 
                           n9297, ZN => n2135);
   U8727 : OAI22_X1 port map( A1 => n11925, A2 => n12439, B1 => n9878, B2 => 
                           n9296, ZN => n2136);
   U8728 : OAI22_X1 port map( A1 => n11925, A2 => n12443, B1 => n9878, B2 => 
                           n9295, ZN => n2137);
   U8729 : OAI22_X1 port map( A1 => n11925, A2 => n12447, B1 => n12325, B2 => 
                           n9294, ZN => n2138);
   U8730 : OAI22_X1 port map( A1 => n11925, A2 => n12451, B1 => n12325, B2 => 
                           n9293, ZN => n2139);
   U8731 : OAI22_X1 port map( A1 => n11925, A2 => n12455, B1 => n12325, B2 => 
                           n9292, ZN => n2140);
   U8732 : OAI22_X1 port map( A1 => n11925, A2 => n12459, B1 => n12325, B2 => 
                           n9291, ZN => n2141);
   U8733 : OAI22_X1 port map( A1 => n11925, A2 => n12463, B1 => n12325, B2 => 
                           n9290, ZN => n2142);
   U8734 : OAI22_X1 port map( A1 => n11924, A2 => n12467, B1 => n12325, B2 => 
                           n9289, ZN => n2143);
   U8735 : OAI22_X1 port map( A1 => n11924, A2 => n12471, B1 => n12325, B2 => 
                           n9288, ZN => n2144);
   U8736 : OAI22_X1 port map( A1 => n11924, A2 => n12475, B1 => n12325, B2 => 
                           n9287, ZN => n2145);
   U8737 : OAI22_X1 port map( A1 => n11924, A2 => n12479, B1 => n12325, B2 => 
                           n9286, ZN => n2146);
   U8738 : OAI22_X1 port map( A1 => n11924, A2 => n12483, B1 => n9878, B2 => 
                           n9285, ZN => n2147);
   U8739 : OAI22_X1 port map( A1 => n11924, A2 => n12487, B1 => n9878, B2 => 
                           n9284, ZN => n2148);
   U8740 : OAI22_X1 port map( A1 => n11924, A2 => n12491, B1 => n9878, B2 => 
                           n9283, ZN => n2149);
   U8741 : OAI22_X1 port map( A1 => n11924, A2 => n12495, B1 => n9878, B2 => 
                           n9282, ZN => n2150);
   U8742 : OAI22_X1 port map( A1 => n11924, A2 => n12499, B1 => n9878, B2 => 
                           n9281, ZN => n2151);
   U8743 : OAI22_X1 port map( A1 => n11924, A2 => n12503, B1 => n9878, B2 => 
                           n9280, ZN => n2152);
   U8744 : OAI22_X1 port map( A1 => n11924, A2 => n12507, B1 => n9878, B2 => 
                           n9279, ZN => n2153);
   U8745 : OAI22_X1 port map( A1 => n11924, A2 => n12515, B1 => n9878, B2 => 
                           n9278, ZN => n2154);
   U8746 : OAI22_X1 port map( A1 => n11947, A2 => n12386, B1 => n12353, B2 => 
                           n9085, ZN => n2347);
   U8747 : OAI22_X1 port map( A1 => n11947, A2 => n12390, B1 => n12353, B2 => 
                           n9084, ZN => n2348);
   U8748 : OAI22_X1 port map( A1 => n11947, A2 => n12394, B1 => n12353, B2 => 
                           n9083, ZN => n2349);
   U8749 : OAI22_X1 port map( A1 => n11947, A2 => n12398, B1 => n12353, B2 => 
                           n9082, ZN => n2350);
   U8750 : OAI22_X1 port map( A1 => n11947, A2 => n12402, B1 => n12353, B2 => 
                           n9081, ZN => n2351);
   U8751 : OAI22_X1 port map( A1 => n11947, A2 => n12406, B1 => n12353, B2 => 
                           n9080, ZN => n2352);
   U8752 : OAI22_X1 port map( A1 => n11947, A2 => n12410, B1 => n12353, B2 => 
                           n9079, ZN => n2353);
   U8753 : OAI22_X1 port map( A1 => n11947, A2 => n12414, B1 => n12353, B2 => 
                           n9078, ZN => n2354);
   U8754 : OAI22_X1 port map( A1 => n11946, A2 => n12418, B1 => n12353, B2 => 
                           n9077, ZN => n2355);
   U8755 : OAI22_X1 port map( A1 => n11946, A2 => n12422, B1 => n12353, B2 => 
                           n9076, ZN => n2356);
   U8756 : OAI22_X1 port map( A1 => n11946, A2 => n12426, B1 => n12353, B2 => 
                           n9075, ZN => n2357);
   U8757 : OAI22_X1 port map( A1 => n11946, A2 => n12430, B1 => n12353, B2 => 
                           n9074, ZN => n2358);
   U8758 : OAI22_X1 port map( A1 => n11946, A2 => n12434, B1 => n9869, B2 => 
                           n9073, ZN => n2359);
   U8759 : OAI22_X1 port map( A1 => n11946, A2 => n12438, B1 => n9869, B2 => 
                           n9072, ZN => n2360);
   U8760 : OAI22_X1 port map( A1 => n11946, A2 => n12442, B1 => n9869, B2 => 
                           n9071, ZN => n2361);
   U8761 : OAI22_X1 port map( A1 => n11946, A2 => n12446, B1 => n12353, B2 => 
                           n9070, ZN => n2362);
   U8762 : OAI22_X1 port map( A1 => n11946, A2 => n12450, B1 => n12353, B2 => 
                           n9069, ZN => n2363);
   U8763 : OAI22_X1 port map( A1 => n11946, A2 => n12454, B1 => n12353, B2 => 
                           n9068, ZN => n2364);
   U8764 : OAI22_X1 port map( A1 => n11946, A2 => n12458, B1 => n12353, B2 => 
                           n9067, ZN => n2365);
   U8765 : OAI22_X1 port map( A1 => n11946, A2 => n12462, B1 => n12353, B2 => 
                           n9066, ZN => n2366);
   U8766 : OAI22_X1 port map( A1 => n11945, A2 => n12466, B1 => n12353, B2 => 
                           n9065, ZN => n2367);
   U8767 : OAI22_X1 port map( A1 => n11945, A2 => n12470, B1 => n12353, B2 => 
                           n9064, ZN => n2368);
   U8768 : OAI22_X1 port map( A1 => n11945, A2 => n12474, B1 => n12353, B2 => 
                           n9063, ZN => n2369);
   U8769 : OAI22_X1 port map( A1 => n11945, A2 => n12478, B1 => n12353, B2 => 
                           n9062, ZN => n2370);
   U8770 : OAI22_X1 port map( A1 => n11945, A2 => n12482, B1 => n9869, B2 => 
                           n9061, ZN => n2371);
   U8771 : OAI22_X1 port map( A1 => n11945, A2 => n12486, B1 => n9869, B2 => 
                           n9060, ZN => n2372);
   U8772 : OAI22_X1 port map( A1 => n11945, A2 => n12490, B1 => n9869, B2 => 
                           n9059, ZN => n2373);
   U8773 : OAI22_X1 port map( A1 => n11945, A2 => n12494, B1 => n9869, B2 => 
                           n9058, ZN => n2374);
   U8774 : OAI22_X1 port map( A1 => n11945, A2 => n12498, B1 => n9869, B2 => 
                           n9057, ZN => n2375);
   U8775 : OAI22_X1 port map( A1 => n11945, A2 => n12502, B1 => n9869, B2 => 
                           n9056, ZN => n2376);
   U8776 : OAI22_X1 port map( A1 => n11945, A2 => n12506, B1 => n9869, B2 => 
                           n9055, ZN => n2377);
   U8777 : OAI22_X1 port map( A1 => n11945, A2 => n12514, B1 => n9869, B2 => 
                           n9054, ZN => n2378);
   U8778 : OAI22_X1 port map( A1 => n11959, A2 => n12386, B1 => n12369, B2 => 
                           n8957, ZN => n2475);
   U8779 : OAI22_X1 port map( A1 => n11959, A2 => n12390, B1 => n12369, B2 => 
                           n8956, ZN => n2476);
   U8780 : OAI22_X1 port map( A1 => n11959, A2 => n12394, B1 => n12369, B2 => 
                           n8955, ZN => n2477);
   U8781 : OAI22_X1 port map( A1 => n11959, A2 => n12398, B1 => n12369, B2 => 
                           n8954, ZN => n2478);
   U8782 : OAI22_X1 port map( A1 => n11959, A2 => n12402, B1 => n12369, B2 => 
                           n8953, ZN => n2479);
   U8783 : OAI22_X1 port map( A1 => n11959, A2 => n12406, B1 => n12369, B2 => 
                           n8952, ZN => n2480);
   U8784 : OAI22_X1 port map( A1 => n11959, A2 => n12410, B1 => n12369, B2 => 
                           n8951, ZN => n2481);
   U8785 : OAI22_X1 port map( A1 => n11959, A2 => n12414, B1 => n12369, B2 => 
                           n8950, ZN => n2482);
   U8786 : OAI22_X1 port map( A1 => n11958, A2 => n12418, B1 => n12369, B2 => 
                           n8949, ZN => n2483);
   U8787 : OAI22_X1 port map( A1 => n11958, A2 => n12422, B1 => n12369, B2 => 
                           n8948, ZN => n2484);
   U8788 : OAI22_X1 port map( A1 => n11958, A2 => n12426, B1 => n12369, B2 => 
                           n8947, ZN => n2485);
   U8789 : OAI22_X1 port map( A1 => n11958, A2 => n12430, B1 => n12369, B2 => 
                           n8946, ZN => n2486);
   U8790 : OAI22_X1 port map( A1 => n11958, A2 => n12434, B1 => n9864, B2 => 
                           n8945, ZN => n2487);
   U8791 : OAI22_X1 port map( A1 => n11958, A2 => n12438, B1 => n9864, B2 => 
                           n8944, ZN => n2488);
   U8792 : OAI22_X1 port map( A1 => n11958, A2 => n12442, B1 => n9864, B2 => 
                           n8943, ZN => n2489);
   U8793 : OAI22_X1 port map( A1 => n11958, A2 => n12446, B1 => n12369, B2 => 
                           n8942, ZN => n2490);
   U8794 : OAI22_X1 port map( A1 => n11958, A2 => n12450, B1 => n12369, B2 => 
                           n8941, ZN => n2491);
   U8795 : OAI22_X1 port map( A1 => n11958, A2 => n12454, B1 => n12369, B2 => 
                           n8940, ZN => n2492);
   U8796 : OAI22_X1 port map( A1 => n11958, A2 => n12458, B1 => n12369, B2 => 
                           n8939, ZN => n2493);
   U8797 : OAI22_X1 port map( A1 => n11958, A2 => n12462, B1 => n12369, B2 => 
                           n8938, ZN => n2494);
   U8798 : OAI22_X1 port map( A1 => n11957, A2 => n12466, B1 => n12369, B2 => 
                           n8937, ZN => n2495);
   U8799 : OAI22_X1 port map( A1 => n11957, A2 => n12470, B1 => n12369, B2 => 
                           n8936, ZN => n2496);
   U8800 : OAI22_X1 port map( A1 => n11957, A2 => n12474, B1 => n12369, B2 => 
                           n8935, ZN => n2497);
   U8801 : OAI22_X1 port map( A1 => n11957, A2 => n12478, B1 => n12369, B2 => 
                           n8934, ZN => n2498);
   U8802 : OAI22_X1 port map( A1 => n11957, A2 => n12482, B1 => n9864, B2 => 
                           n8933, ZN => n2499);
   U8803 : OAI22_X1 port map( A1 => n11957, A2 => n12486, B1 => n9864, B2 => 
                           n8932, ZN => n2500);
   U8804 : OAI22_X1 port map( A1 => n11957, A2 => n12490, B1 => n9864, B2 => 
                           n8931, ZN => n2501);
   U8805 : OAI22_X1 port map( A1 => n11957, A2 => n12494, B1 => n9864, B2 => 
                           n8930, ZN => n2502);
   U8806 : OAI22_X1 port map( A1 => n11957, A2 => n12498, B1 => n9864, B2 => 
                           n8929, ZN => n2503);
   U8807 : OAI22_X1 port map( A1 => n11957, A2 => n12502, B1 => n9864, B2 => 
                           n8928, ZN => n2504);
   U8808 : OAI22_X1 port map( A1 => n11957, A2 => n12506, B1 => n9864, B2 => 
                           n8927, ZN => n2505);
   U8809 : OAI22_X1 port map( A1 => n11957, A2 => n12514, B1 => n9864, B2 => 
                           n8926, ZN => n2506);
   U8810 : OAI22_X1 port map( A1 => n11962, A2 => n12386, B1 => n12373, B2 => 
                           n8925, ZN => n2507);
   U8811 : OAI22_X1 port map( A1 => n11962, A2 => n12390, B1 => n12373, B2 => 
                           n8924, ZN => n2508);
   U8812 : OAI22_X1 port map( A1 => n11962, A2 => n12394, B1 => n12373, B2 => 
                           n8923, ZN => n2509);
   U8813 : OAI22_X1 port map( A1 => n11962, A2 => n12398, B1 => n12373, B2 => 
                           n8922, ZN => n2510);
   U8814 : OAI22_X1 port map( A1 => n11962, A2 => n12402, B1 => n12373, B2 => 
                           n8921, ZN => n2511);
   U8815 : OAI22_X1 port map( A1 => n11962, A2 => n12406, B1 => n12373, B2 => 
                           n8920, ZN => n2512);
   U8816 : OAI22_X1 port map( A1 => n11962, A2 => n12410, B1 => n12373, B2 => 
                           n8919, ZN => n2513);
   U8817 : OAI22_X1 port map( A1 => n11962, A2 => n12414, B1 => n12373, B2 => 
                           n8918, ZN => n2514);
   U8818 : OAI22_X1 port map( A1 => n11961, A2 => n12418, B1 => n12373, B2 => 
                           n8917, ZN => n2515);
   U8819 : OAI22_X1 port map( A1 => n11961, A2 => n12422, B1 => n12373, B2 => 
                           n8916, ZN => n2516);
   U8820 : OAI22_X1 port map( A1 => n11961, A2 => n12426, B1 => n12373, B2 => 
                           n8915, ZN => n2517);
   U8821 : OAI22_X1 port map( A1 => n11961, A2 => n12430, B1 => n12373, B2 => 
                           n8914, ZN => n2518);
   U8822 : OAI22_X1 port map( A1 => n11961, A2 => n12434, B1 => n9861, B2 => 
                           n8913, ZN => n2519);
   U8823 : OAI22_X1 port map( A1 => n11961, A2 => n12438, B1 => n9861, B2 => 
                           n8912, ZN => n2520);
   U8824 : OAI22_X1 port map( A1 => n11961, A2 => n12442, B1 => n9861, B2 => 
                           n8911, ZN => n2521);
   U8825 : OAI22_X1 port map( A1 => n11961, A2 => n12446, B1 => n12373, B2 => 
                           n8910, ZN => n2522);
   U8826 : OAI22_X1 port map( A1 => n11961, A2 => n12450, B1 => n12373, B2 => 
                           n8909, ZN => n2523);
   U8827 : OAI22_X1 port map( A1 => n11961, A2 => n12454, B1 => n12373, B2 => 
                           n8908, ZN => n2524);
   U8828 : OAI22_X1 port map( A1 => n11961, A2 => n12458, B1 => n12373, B2 => 
                           n8907, ZN => n2525);
   U8829 : OAI22_X1 port map( A1 => n11961, A2 => n12462, B1 => n12373, B2 => 
                           n8906, ZN => n2526);
   U8830 : OAI22_X1 port map( A1 => n11960, A2 => n12466, B1 => n12373, B2 => 
                           n8905, ZN => n2527);
   U8831 : OAI22_X1 port map( A1 => n11960, A2 => n12470, B1 => n12373, B2 => 
                           n8904, ZN => n2528);
   U8832 : OAI22_X1 port map( A1 => n11960, A2 => n12474, B1 => n12373, B2 => 
                           n8903, ZN => n2529);
   U8833 : OAI22_X1 port map( A1 => n11960, A2 => n12478, B1 => n12373, B2 => 
                           n8902, ZN => n2530);
   U8834 : OAI22_X1 port map( A1 => n11960, A2 => n12482, B1 => n9861, B2 => 
                           n8901, ZN => n2531);
   U8835 : OAI22_X1 port map( A1 => n11960, A2 => n12486, B1 => n9861, B2 => 
                           n8900, ZN => n2532);
   U8836 : OAI22_X1 port map( A1 => n11960, A2 => n12490, B1 => n9861, B2 => 
                           n8899, ZN => n2533);
   U8837 : OAI22_X1 port map( A1 => n11960, A2 => n12494, B1 => n9861, B2 => 
                           n8898, ZN => n2534);
   U8838 : OAI22_X1 port map( A1 => n11960, A2 => n12498, B1 => n9861, B2 => 
                           n8897, ZN => n2535);
   U8839 : OAI22_X1 port map( A1 => n11960, A2 => n12502, B1 => n9861, B2 => 
                           n8896, ZN => n2536);
   U8840 : OAI22_X1 port map( A1 => n11960, A2 => n12506, B1 => n9861, B2 => 
                           n8895, ZN => n2537);
   U8841 : OAI22_X1 port map( A1 => n11960, A2 => n12514, B1 => n9861, B2 => 
                           n8894, ZN => n2538);
   U8842 : OAI22_X1 port map( A1 => n11905, A2 => n12387, B1 => n12297, B2 => 
                           n9533, ZN => n1899);
   U8843 : OAI22_X1 port map( A1 => n11905, A2 => n12391, B1 => n12297, B2 => 
                           n9532, ZN => n1900);
   U8844 : OAI22_X1 port map( A1 => n11905, A2 => n12395, B1 => n12297, B2 => 
                           n9531, ZN => n1901);
   U8845 : OAI22_X1 port map( A1 => n11905, A2 => n12399, B1 => n12297, B2 => 
                           n9530, ZN => n1902);
   U8846 : OAI22_X1 port map( A1 => n11905, A2 => n12403, B1 => n12297, B2 => 
                           n9529, ZN => n1903);
   U8847 : OAI22_X1 port map( A1 => n11905, A2 => n12407, B1 => n12297, B2 => 
                           n9528, ZN => n1904);
   U8848 : OAI22_X1 port map( A1 => n11905, A2 => n12411, B1 => n12297, B2 => 
                           n9527, ZN => n1905);
   U8849 : OAI22_X1 port map( A1 => n11905, A2 => n12415, B1 => n12297, B2 => 
                           n9526, ZN => n1906);
   U8850 : OAI22_X1 port map( A1 => n11904, A2 => n12419, B1 => n12297, B2 => 
                           n9525, ZN => n1907);
   U8851 : OAI22_X1 port map( A1 => n11904, A2 => n12423, B1 => n12297, B2 => 
                           n9524, ZN => n1908);
   U8852 : OAI22_X1 port map( A1 => n11904, A2 => n12427, B1 => n12297, B2 => 
                           n9523, ZN => n1909);
   U8853 : OAI22_X1 port map( A1 => n11904, A2 => n12431, B1 => n12297, B2 => 
                           n9522, ZN => n1910);
   U8854 : OAI22_X1 port map( A1 => n11904, A2 => n12435, B1 => n9888, B2 => 
                           n9521, ZN => n1911);
   U8855 : OAI22_X1 port map( A1 => n11904, A2 => n12439, B1 => n9888, B2 => 
                           n9520, ZN => n1912);
   U8856 : OAI22_X1 port map( A1 => n11904, A2 => n12443, B1 => n9888, B2 => 
                           n9519, ZN => n1913);
   U8857 : OAI22_X1 port map( A1 => n11904, A2 => n12447, B1 => n12297, B2 => 
                           n9518, ZN => n1914);
   U8858 : OAI22_X1 port map( A1 => n11904, A2 => n12451, B1 => n12297, B2 => 
                           n9517, ZN => n1915);
   U8859 : OAI22_X1 port map( A1 => n11904, A2 => n12455, B1 => n12297, B2 => 
                           n9516, ZN => n1916);
   U8860 : OAI22_X1 port map( A1 => n11904, A2 => n12459, B1 => n12297, B2 => 
                           n9515, ZN => n1917);
   U8861 : OAI22_X1 port map( A1 => n11904, A2 => n12463, B1 => n12297, B2 => 
                           n9514, ZN => n1918);
   U8862 : OAI22_X1 port map( A1 => n11903, A2 => n12467, B1 => n12297, B2 => 
                           n9513, ZN => n1919);
   U8863 : OAI22_X1 port map( A1 => n11903, A2 => n12471, B1 => n12297, B2 => 
                           n9512, ZN => n1920);
   U8864 : OAI22_X1 port map( A1 => n11903, A2 => n12475, B1 => n12297, B2 => 
                           n9511, ZN => n1921);
   U8865 : OAI22_X1 port map( A1 => n11903, A2 => n12479, B1 => n12297, B2 => 
                           n9510, ZN => n1922);
   U8866 : OAI22_X1 port map( A1 => n11903, A2 => n12483, B1 => n9888, B2 => 
                           n9509, ZN => n1923);
   U8867 : OAI22_X1 port map( A1 => n11903, A2 => n12487, B1 => n9888, B2 => 
                           n9508, ZN => n1924);
   U8868 : OAI22_X1 port map( A1 => n11903, A2 => n12491, B1 => n9888, B2 => 
                           n9507, ZN => n1925);
   U8869 : OAI22_X1 port map( A1 => n11903, A2 => n12495, B1 => n9888, B2 => 
                           n9506, ZN => n1926);
   U8870 : OAI22_X1 port map( A1 => n11903, A2 => n12499, B1 => n9888, B2 => 
                           n9505, ZN => n1927);
   U8871 : OAI22_X1 port map( A1 => n11903, A2 => n12503, B1 => n9888, B2 => 
                           n9504, ZN => n1928);
   U8872 : OAI22_X1 port map( A1 => n11903, A2 => n12507, B1 => n9888, B2 => 
                           n9503, ZN => n1929);
   U8873 : OAI22_X1 port map( A1 => n11903, A2 => n12515, B1 => n9888, B2 => 
                           n9502, ZN => n1930);
   U8874 : OAI22_X1 port map( A1 => n11923, A2 => n12387, B1 => n12321, B2 => 
                           n9341, ZN => n2091);
   U8875 : OAI22_X1 port map( A1 => n11923, A2 => n12391, B1 => n12321, B2 => 
                           n9340, ZN => n2092);
   U8876 : OAI22_X1 port map( A1 => n11923, A2 => n12395, B1 => n12321, B2 => 
                           n9339, ZN => n2093);
   U8877 : OAI22_X1 port map( A1 => n11923, A2 => n12399, B1 => n12321, B2 => 
                           n9338, ZN => n2094);
   U8878 : OAI22_X1 port map( A1 => n11923, A2 => n12403, B1 => n12321, B2 => 
                           n9337, ZN => n2095);
   U8879 : OAI22_X1 port map( A1 => n11923, A2 => n12407, B1 => n12321, B2 => 
                           n9336, ZN => n2096);
   U8880 : OAI22_X1 port map( A1 => n11923, A2 => n12411, B1 => n12321, B2 => 
                           n9335, ZN => n2097);
   U8881 : OAI22_X1 port map( A1 => n11923, A2 => n12415, B1 => n12321, B2 => 
                           n9334, ZN => n2098);
   U8882 : OAI22_X1 port map( A1 => n11922, A2 => n12419, B1 => n12321, B2 => 
                           n9333, ZN => n2099);
   U8883 : OAI22_X1 port map( A1 => n11922, A2 => n12423, B1 => n12321, B2 => 
                           n9332, ZN => n2100);
   U8884 : OAI22_X1 port map( A1 => n11922, A2 => n12427, B1 => n12321, B2 => 
                           n9331, ZN => n2101);
   U8885 : OAI22_X1 port map( A1 => n11922, A2 => n12431, B1 => n12321, B2 => 
                           n9330, ZN => n2102);
   U8886 : OAI22_X1 port map( A1 => n11922, A2 => n12435, B1 => n9879, B2 => 
                           n9329, ZN => n2103);
   U8887 : OAI22_X1 port map( A1 => n11922, A2 => n12439, B1 => n9879, B2 => 
                           n9328, ZN => n2104);
   U8888 : OAI22_X1 port map( A1 => n11922, A2 => n12443, B1 => n9879, B2 => 
                           n9327, ZN => n2105);
   U8889 : OAI22_X1 port map( A1 => n11922, A2 => n12447, B1 => n12321, B2 => 
                           n9326, ZN => n2106);
   U8890 : OAI22_X1 port map( A1 => n11922, A2 => n12451, B1 => n12321, B2 => 
                           n9325, ZN => n2107);
   U8891 : OAI22_X1 port map( A1 => n11922, A2 => n12455, B1 => n12321, B2 => 
                           n9324, ZN => n2108);
   U8892 : OAI22_X1 port map( A1 => n11922, A2 => n12459, B1 => n12321, B2 => 
                           n9323, ZN => n2109);
   U8893 : OAI22_X1 port map( A1 => n11922, A2 => n12463, B1 => n12321, B2 => 
                           n9322, ZN => n2110);
   U8894 : OAI22_X1 port map( A1 => n11921, A2 => n12467, B1 => n12321, B2 => 
                           n9321, ZN => n2111);
   U8895 : OAI22_X1 port map( A1 => n11921, A2 => n12471, B1 => n12321, B2 => 
                           n9320, ZN => n2112);
   U8896 : OAI22_X1 port map( A1 => n11921, A2 => n12475, B1 => n12321, B2 => 
                           n9319, ZN => n2113);
   U8897 : OAI22_X1 port map( A1 => n11921, A2 => n12479, B1 => n12321, B2 => 
                           n9318, ZN => n2114);
   U8898 : OAI22_X1 port map( A1 => n11921, A2 => n12483, B1 => n9879, B2 => 
                           n9317, ZN => n2115);
   U8899 : OAI22_X1 port map( A1 => n11921, A2 => n12487, B1 => n9879, B2 => 
                           n9316, ZN => n2116);
   U8900 : OAI22_X1 port map( A1 => n11921, A2 => n12491, B1 => n9879, B2 => 
                           n9315, ZN => n2117);
   U8901 : OAI22_X1 port map( A1 => n11921, A2 => n12495, B1 => n9879, B2 => 
                           n9314, ZN => n2118);
   U8902 : OAI22_X1 port map( A1 => n11921, A2 => n12499, B1 => n9879, B2 => 
                           n9313, ZN => n2119);
   U8903 : OAI22_X1 port map( A1 => n11921, A2 => n12503, B1 => n9879, B2 => 
                           n9312, ZN => n2120);
   U8904 : OAI22_X1 port map( A1 => n11921, A2 => n12507, B1 => n9879, B2 => 
                           n9311, ZN => n2121);
   U8905 : OAI22_X1 port map( A1 => n11921, A2 => n12515, B1 => n9879, B2 => 
                           n9310, ZN => n2122);
   U8906 : OAI22_X1 port map( A1 => n11911, A2 => n12387, B1 => n12305, B2 => 
                           n9469, ZN => n1963);
   U8907 : OAI22_X1 port map( A1 => n11911, A2 => n12391, B1 => n12305, B2 => 
                           n9468, ZN => n1964);
   U8908 : OAI22_X1 port map( A1 => n11911, A2 => n12395, B1 => n12305, B2 => 
                           n9467, ZN => n1965);
   U8909 : OAI22_X1 port map( A1 => n11911, A2 => n12399, B1 => n12305, B2 => 
                           n9466, ZN => n1966);
   U8910 : OAI22_X1 port map( A1 => n11911, A2 => n12403, B1 => n12305, B2 => 
                           n9465, ZN => n1967);
   U8911 : OAI22_X1 port map( A1 => n11911, A2 => n12407, B1 => n12305, B2 => 
                           n9464, ZN => n1968);
   U8912 : OAI22_X1 port map( A1 => n11911, A2 => n12411, B1 => n12305, B2 => 
                           n9463, ZN => n1969);
   U8913 : OAI22_X1 port map( A1 => n11911, A2 => n12415, B1 => n12305, B2 => 
                           n9462, ZN => n1970);
   U8914 : OAI22_X1 port map( A1 => n11910, A2 => n12419, B1 => n12305, B2 => 
                           n9461, ZN => n1971);
   U8915 : OAI22_X1 port map( A1 => n11910, A2 => n12423, B1 => n12305, B2 => 
                           n9460, ZN => n1972);
   U8916 : OAI22_X1 port map( A1 => n11910, A2 => n12427, B1 => n12305, B2 => 
                           n9459, ZN => n1973);
   U8917 : OAI22_X1 port map( A1 => n11910, A2 => n12431, B1 => n12305, B2 => 
                           n9458, ZN => n1974);
   U8918 : OAI22_X1 port map( A1 => n11910, A2 => n12435, B1 => n9885, B2 => 
                           n9457, ZN => n1975);
   U8919 : OAI22_X1 port map( A1 => n11910, A2 => n12439, B1 => n9885, B2 => 
                           n9456, ZN => n1976);
   U8920 : OAI22_X1 port map( A1 => n11910, A2 => n12443, B1 => n9885, B2 => 
                           n9455, ZN => n1977);
   U8921 : OAI22_X1 port map( A1 => n11910, A2 => n12447, B1 => n12305, B2 => 
                           n9454, ZN => n1978);
   U8922 : OAI22_X1 port map( A1 => n11910, A2 => n12451, B1 => n12305, B2 => 
                           n9453, ZN => n1979);
   U8923 : OAI22_X1 port map( A1 => n11910, A2 => n12455, B1 => n12305, B2 => 
                           n9452, ZN => n1980);
   U8924 : OAI22_X1 port map( A1 => n11910, A2 => n12459, B1 => n12305, B2 => 
                           n9451, ZN => n1981);
   U8925 : OAI22_X1 port map( A1 => n11910, A2 => n12463, B1 => n12305, B2 => 
                           n9450, ZN => n1982);
   U8926 : OAI22_X1 port map( A1 => n11909, A2 => n12467, B1 => n12305, B2 => 
                           n9449, ZN => n1983);
   U8927 : OAI22_X1 port map( A1 => n11909, A2 => n12471, B1 => n12305, B2 => 
                           n9448, ZN => n1984);
   U8928 : OAI22_X1 port map( A1 => n11909, A2 => n12475, B1 => n12305, B2 => 
                           n9447, ZN => n1985);
   U8929 : OAI22_X1 port map( A1 => n11909, A2 => n12479, B1 => n12305, B2 => 
                           n9446, ZN => n1986);
   U8930 : OAI22_X1 port map( A1 => n11909, A2 => n12483, B1 => n9885, B2 => 
                           n9445, ZN => n1987);
   U8931 : OAI22_X1 port map( A1 => n11909, A2 => n12487, B1 => n9885, B2 => 
                           n9444, ZN => n1988);
   U8932 : OAI22_X1 port map( A1 => n11909, A2 => n12491, B1 => n9885, B2 => 
                           n9443, ZN => n1989);
   U8933 : OAI22_X1 port map( A1 => n11909, A2 => n12495, B1 => n9885, B2 => 
                           n9442, ZN => n1990);
   U8934 : OAI22_X1 port map( A1 => n11909, A2 => n12499, B1 => n9885, B2 => 
                           n9441, ZN => n1991);
   U8935 : OAI22_X1 port map( A1 => n11909, A2 => n12503, B1 => n9885, B2 => 
                           n9440, ZN => n1992);
   U8936 : OAI22_X1 port map( A1 => n11909, A2 => n12507, B1 => n9885, B2 => 
                           n9439, ZN => n1993);
   U8937 : OAI22_X1 port map( A1 => n11909, A2 => n12515, B1 => n9885, B2 => 
                           n9438, ZN => n1994);
   U8938 : OAI22_X1 port map( A1 => n11884, A2 => n12388, B1 => n12269, B2 => 
                           n9757, ZN => n1675);
   U8939 : OAI22_X1 port map( A1 => n11884, A2 => n12392, B1 => n12269, B2 => 
                           n9756, ZN => n1676);
   U8940 : OAI22_X1 port map( A1 => n11884, A2 => n12396, B1 => n12269, B2 => 
                           n9755, ZN => n1677);
   U8941 : OAI22_X1 port map( A1 => n11884, A2 => n12400, B1 => n12269, B2 => 
                           n9754, ZN => n1678);
   U8942 : OAI22_X1 port map( A1 => n11884, A2 => n12404, B1 => n12269, B2 => 
                           n9753, ZN => n1679);
   U8943 : OAI22_X1 port map( A1 => n11884, A2 => n12408, B1 => n12269, B2 => 
                           n9752, ZN => n1680);
   U8944 : OAI22_X1 port map( A1 => n11884, A2 => n12412, B1 => n12269, B2 => 
                           n9751, ZN => n1681);
   U8945 : OAI22_X1 port map( A1 => n11884, A2 => n12416, B1 => n12269, B2 => 
                           n9750, ZN => n1682);
   U8946 : OAI22_X1 port map( A1 => n11883, A2 => n12420, B1 => n12269, B2 => 
                           n9749, ZN => n1683);
   U8947 : OAI22_X1 port map( A1 => n11883, A2 => n12424, B1 => n12269, B2 => 
                           n9748, ZN => n1684);
   U8948 : OAI22_X1 port map( A1 => n11883, A2 => n12428, B1 => n12269, B2 => 
                           n9747, ZN => n1685);
   U8949 : OAI22_X1 port map( A1 => n11883, A2 => n12432, B1 => n12269, B2 => 
                           n9746, ZN => n1686);
   U8950 : OAI22_X1 port map( A1 => n11883, A2 => n12436, B1 => n9897, B2 => 
                           n9745, ZN => n1687);
   U8951 : OAI22_X1 port map( A1 => n11883, A2 => n12440, B1 => n9897, B2 => 
                           n9744, ZN => n1688);
   U8952 : OAI22_X1 port map( A1 => n11883, A2 => n12444, B1 => n9897, B2 => 
                           n9743, ZN => n1689);
   U8953 : OAI22_X1 port map( A1 => n11883, A2 => n12448, B1 => n12269, B2 => 
                           n9742, ZN => n1690);
   U8954 : OAI22_X1 port map( A1 => n11883, A2 => n12452, B1 => n12269, B2 => 
                           n9741, ZN => n1691);
   U8955 : OAI22_X1 port map( A1 => n11883, A2 => n12456, B1 => n12269, B2 => 
                           n9740, ZN => n1692);
   U8956 : OAI22_X1 port map( A1 => n11883, A2 => n12460, B1 => n12269, B2 => 
                           n9739, ZN => n1693);
   U8957 : OAI22_X1 port map( A1 => n11883, A2 => n12464, B1 => n12269, B2 => 
                           n9738, ZN => n1694);
   U8958 : OAI22_X1 port map( A1 => n11882, A2 => n12468, B1 => n12269, B2 => 
                           n9737, ZN => n1695);
   U8959 : OAI22_X1 port map( A1 => n11882, A2 => n12472, B1 => n12269, B2 => 
                           n9736, ZN => n1696);
   U8960 : OAI22_X1 port map( A1 => n11882, A2 => n12476, B1 => n12269, B2 => 
                           n9735, ZN => n1697);
   U8961 : OAI22_X1 port map( A1 => n11882, A2 => n12480, B1 => n12269, B2 => 
                           n9734, ZN => n1698);
   U8962 : OAI22_X1 port map( A1 => n11882, A2 => n12484, B1 => n9897, B2 => 
                           n9733, ZN => n1699);
   U8963 : OAI22_X1 port map( A1 => n11882, A2 => n12488, B1 => n9897, B2 => 
                           n9732, ZN => n1700);
   U8964 : OAI22_X1 port map( A1 => n11882, A2 => n12492, B1 => n9897, B2 => 
                           n9731, ZN => n1701);
   U8965 : OAI22_X1 port map( A1 => n11882, A2 => n12496, B1 => n9897, B2 => 
                           n9730, ZN => n1702);
   U8966 : OAI22_X1 port map( A1 => n11882, A2 => n12500, B1 => n9897, B2 => 
                           n9729, ZN => n1703);
   U8967 : OAI22_X1 port map( A1 => n11882, A2 => n12504, B1 => n9897, B2 => 
                           n9728, ZN => n1704);
   U8968 : OAI22_X1 port map( A1 => n11882, A2 => n12508, B1 => n9897, B2 => 
                           n9727, ZN => n1705);
   U8969 : OAI22_X1 port map( A1 => n11882, A2 => n12516, B1 => n9897, B2 => 
                           n9726, ZN => n1706);
   U8970 : OAI22_X1 port map( A1 => n11893, A2 => n12388, B1 => n12281, B2 => 
                           n9661, ZN => n1771);
   U8971 : OAI22_X1 port map( A1 => n11893, A2 => n12392, B1 => n12281, B2 => 
                           n9660, ZN => n1772);
   U8972 : OAI22_X1 port map( A1 => n11893, A2 => n12396, B1 => n12281, B2 => 
                           n9659, ZN => n1773);
   U8973 : OAI22_X1 port map( A1 => n11893, A2 => n12400, B1 => n12281, B2 => 
                           n9658, ZN => n1774);
   U8974 : OAI22_X1 port map( A1 => n11893, A2 => n12404, B1 => n12281, B2 => 
                           n9657, ZN => n1775);
   U8975 : OAI22_X1 port map( A1 => n11893, A2 => n12408, B1 => n12281, B2 => 
                           n9656, ZN => n1776);
   U8976 : OAI22_X1 port map( A1 => n11893, A2 => n12412, B1 => n12281, B2 => 
                           n9655, ZN => n1777);
   U8977 : OAI22_X1 port map( A1 => n11893, A2 => n12416, B1 => n12281, B2 => 
                           n9654, ZN => n1778);
   U8978 : OAI22_X1 port map( A1 => n11892, A2 => n12420, B1 => n12281, B2 => 
                           n9653, ZN => n1779);
   U8979 : OAI22_X1 port map( A1 => n11892, A2 => n12424, B1 => n12281, B2 => 
                           n9652, ZN => n1780);
   U8980 : OAI22_X1 port map( A1 => n11892, A2 => n12428, B1 => n12281, B2 => 
                           n9651, ZN => n1781);
   U8981 : OAI22_X1 port map( A1 => n11892, A2 => n12432, B1 => n12281, B2 => 
                           n9650, ZN => n1782);
   U8982 : OAI22_X1 port map( A1 => n11892, A2 => n12436, B1 => n9893, B2 => 
                           n9649, ZN => n1783);
   U8983 : OAI22_X1 port map( A1 => n11892, A2 => n12440, B1 => n9893, B2 => 
                           n9648, ZN => n1784);
   U8984 : OAI22_X1 port map( A1 => n11892, A2 => n12444, B1 => n9893, B2 => 
                           n9647, ZN => n1785);
   U8985 : OAI22_X1 port map( A1 => n11892, A2 => n12448, B1 => n12281, B2 => 
                           n9646, ZN => n1786);
   U8986 : OAI22_X1 port map( A1 => n11892, A2 => n12452, B1 => n12281, B2 => 
                           n9645, ZN => n1787);
   U8987 : OAI22_X1 port map( A1 => n11892, A2 => n12456, B1 => n12281, B2 => 
                           n9644, ZN => n1788);
   U8988 : OAI22_X1 port map( A1 => n11892, A2 => n12460, B1 => n12281, B2 => 
                           n9643, ZN => n1789);
   U8989 : OAI22_X1 port map( A1 => n11892, A2 => n12464, B1 => n12281, B2 => 
                           n9642, ZN => n1790);
   U8990 : OAI22_X1 port map( A1 => n11891, A2 => n12468, B1 => n12281, B2 => 
                           n9641, ZN => n1791);
   U8991 : OAI22_X1 port map( A1 => n11891, A2 => n12472, B1 => n12281, B2 => 
                           n9640, ZN => n1792);
   U8992 : OAI22_X1 port map( A1 => n11891, A2 => n12476, B1 => n12281, B2 => 
                           n9639, ZN => n1793);
   U8993 : OAI22_X1 port map( A1 => n11891, A2 => n12480, B1 => n12281, B2 => 
                           n9638, ZN => n1794);
   U8994 : OAI22_X1 port map( A1 => n11891, A2 => n12484, B1 => n9893, B2 => 
                           n9637, ZN => n1795);
   U8995 : OAI22_X1 port map( A1 => n11891, A2 => n12488, B1 => n9893, B2 => 
                           n9636, ZN => n1796);
   U8996 : OAI22_X1 port map( A1 => n11891, A2 => n12492, B1 => n9893, B2 => 
                           n9635, ZN => n1797);
   U8997 : OAI22_X1 port map( A1 => n11891, A2 => n12496, B1 => n9893, B2 => 
                           n9634, ZN => n1798);
   U8998 : OAI22_X1 port map( A1 => n11891, A2 => n12500, B1 => n9893, B2 => 
                           n9633, ZN => n1799);
   U8999 : OAI22_X1 port map( A1 => n11891, A2 => n12504, B1 => n9893, B2 => 
                           n9632, ZN => n1800);
   U9000 : OAI22_X1 port map( A1 => n11891, A2 => n12508, B1 => n9893, B2 => 
                           n9631, ZN => n1801);
   U9001 : OAI22_X1 port map( A1 => n11891, A2 => n12516, B1 => n9893, B2 => 
                           n9630, ZN => n1802);
   U9002 : OAI22_X1 port map( A1 => n11935, A2 => n12387, B1 => n12337, B2 => 
                           n9213, ZN => n2219);
   U9003 : OAI22_X1 port map( A1 => n11935, A2 => n12391, B1 => n12337, B2 => 
                           n9212, ZN => n2220);
   U9004 : OAI22_X1 port map( A1 => n11935, A2 => n12395, B1 => n12337, B2 => 
                           n9211, ZN => n2221);
   U9005 : OAI22_X1 port map( A1 => n11935, A2 => n12399, B1 => n12337, B2 => 
                           n9210, ZN => n2222);
   U9006 : OAI22_X1 port map( A1 => n11935, A2 => n12403, B1 => n12337, B2 => 
                           n9209, ZN => n2223);
   U9007 : OAI22_X1 port map( A1 => n11935, A2 => n12407, B1 => n12337, B2 => 
                           n9208, ZN => n2224);
   U9008 : OAI22_X1 port map( A1 => n11935, A2 => n12411, B1 => n12337, B2 => 
                           n9207, ZN => n2225);
   U9009 : OAI22_X1 port map( A1 => n11935, A2 => n12415, B1 => n12337, B2 => 
                           n9206, ZN => n2226);
   U9010 : OAI22_X1 port map( A1 => n11934, A2 => n12419, B1 => n12337, B2 => 
                           n9205, ZN => n2227);
   U9011 : OAI22_X1 port map( A1 => n11934, A2 => n12423, B1 => n12337, B2 => 
                           n9204, ZN => n2228);
   U9012 : OAI22_X1 port map( A1 => n11934, A2 => n12427, B1 => n12337, B2 => 
                           n9203, ZN => n2229);
   U9013 : OAI22_X1 port map( A1 => n11934, A2 => n12431, B1 => n12337, B2 => 
                           n9202, ZN => n2230);
   U9014 : OAI22_X1 port map( A1 => n11934, A2 => n12435, B1 => n9874, B2 => 
                           n9201, ZN => n2231);
   U9015 : OAI22_X1 port map( A1 => n11934, A2 => n12439, B1 => n9874, B2 => 
                           n9200, ZN => n2232);
   U9016 : OAI22_X1 port map( A1 => n11934, A2 => n12443, B1 => n9874, B2 => 
                           n9199, ZN => n2233);
   U9017 : OAI22_X1 port map( A1 => n11934, A2 => n12447, B1 => n12337, B2 => 
                           n9198, ZN => n2234);
   U9018 : OAI22_X1 port map( A1 => n11934, A2 => n12451, B1 => n12337, B2 => 
                           n9197, ZN => n2235);
   U9019 : OAI22_X1 port map( A1 => n11934, A2 => n12455, B1 => n12337, B2 => 
                           n9196, ZN => n2236);
   U9020 : OAI22_X1 port map( A1 => n11934, A2 => n12459, B1 => n12337, B2 => 
                           n9195, ZN => n2237);
   U9021 : OAI22_X1 port map( A1 => n11934, A2 => n12463, B1 => n12337, B2 => 
                           n9194, ZN => n2238);
   U9022 : OAI22_X1 port map( A1 => n11933, A2 => n12467, B1 => n12337, B2 => 
                           n9193, ZN => n2239);
   U9023 : OAI22_X1 port map( A1 => n11933, A2 => n12471, B1 => n12337, B2 => 
                           n9192, ZN => n2240);
   U9024 : OAI22_X1 port map( A1 => n11933, A2 => n12475, B1 => n12337, B2 => 
                           n9191, ZN => n2241);
   U9025 : OAI22_X1 port map( A1 => n11933, A2 => n12479, B1 => n12337, B2 => 
                           n9190, ZN => n2242);
   U9026 : OAI22_X1 port map( A1 => n11933, A2 => n12483, B1 => n9874, B2 => 
                           n9189, ZN => n2243);
   U9027 : OAI22_X1 port map( A1 => n11933, A2 => n12487, B1 => n9874, B2 => 
                           n9188, ZN => n2244);
   U9028 : OAI22_X1 port map( A1 => n11933, A2 => n12491, B1 => n9874, B2 => 
                           n9187, ZN => n2245);
   U9029 : OAI22_X1 port map( A1 => n11933, A2 => n12495, B1 => n9874, B2 => 
                           n9186, ZN => n2246);
   U9030 : OAI22_X1 port map( A1 => n11933, A2 => n12499, B1 => n9874, B2 => 
                           n9185, ZN => n2247);
   U9031 : OAI22_X1 port map( A1 => n11933, A2 => n12503, B1 => n9874, B2 => 
                           n9184, ZN => n2248);
   U9032 : OAI22_X1 port map( A1 => n11933, A2 => n12507, B1 => n9874, B2 => 
                           n9183, ZN => n2249);
   U9033 : OAI22_X1 port map( A1 => n11933, A2 => n12515, B1 => n9874, B2 => 
                           n9182, ZN => n2250);
   U9034 : OAI22_X1 port map( A1 => n11938, A2 => n12386, B1 => n12341, B2 => 
                           n9181, ZN => n2251);
   U9035 : OAI22_X1 port map( A1 => n11938, A2 => n12390, B1 => n12341, B2 => 
                           n9180, ZN => n2252);
   U9036 : OAI22_X1 port map( A1 => n11938, A2 => n12394, B1 => n12341, B2 => 
                           n9179, ZN => n2253);
   U9037 : OAI22_X1 port map( A1 => n11938, A2 => n12398, B1 => n12341, B2 => 
                           n9178, ZN => n2254);
   U9038 : OAI22_X1 port map( A1 => n11938, A2 => n12402, B1 => n12341, B2 => 
                           n9177, ZN => n2255);
   U9039 : OAI22_X1 port map( A1 => n11938, A2 => n12406, B1 => n12341, B2 => 
                           n9176, ZN => n2256);
   U9040 : OAI22_X1 port map( A1 => n11938, A2 => n12410, B1 => n12341, B2 => 
                           n9175, ZN => n2257);
   U9041 : OAI22_X1 port map( A1 => n11938, A2 => n12414, B1 => n12341, B2 => 
                           n9174, ZN => n2258);
   U9042 : OAI22_X1 port map( A1 => n11937, A2 => n12418, B1 => n12341, B2 => 
                           n9173, ZN => n2259);
   U9043 : OAI22_X1 port map( A1 => n11937, A2 => n12422, B1 => n12341, B2 => 
                           n9172, ZN => n2260);
   U9044 : OAI22_X1 port map( A1 => n11937, A2 => n12426, B1 => n12341, B2 => 
                           n9171, ZN => n2261);
   U9045 : OAI22_X1 port map( A1 => n11937, A2 => n12430, B1 => n12341, B2 => 
                           n9170, ZN => n2262);
   U9046 : OAI22_X1 port map( A1 => n11937, A2 => n12434, B1 => n9873, B2 => 
                           n9169, ZN => n2263);
   U9047 : OAI22_X1 port map( A1 => n11937, A2 => n12438, B1 => n9873, B2 => 
                           n9168, ZN => n2264);
   U9048 : OAI22_X1 port map( A1 => n11937, A2 => n12442, B1 => n9873, B2 => 
                           n9167, ZN => n2265);
   U9049 : OAI22_X1 port map( A1 => n11937, A2 => n12446, B1 => n12341, B2 => 
                           n9166, ZN => n2266);
   U9050 : OAI22_X1 port map( A1 => n11937, A2 => n12450, B1 => n12341, B2 => 
                           n9165, ZN => n2267);
   U9051 : OAI22_X1 port map( A1 => n11937, A2 => n12454, B1 => n12341, B2 => 
                           n9164, ZN => n2268);
   U9052 : OAI22_X1 port map( A1 => n11937, A2 => n12458, B1 => n12341, B2 => 
                           n9163, ZN => n2269);
   U9053 : OAI22_X1 port map( A1 => n11937, A2 => n12462, B1 => n12341, B2 => 
                           n9162, ZN => n2270);
   U9054 : OAI22_X1 port map( A1 => n11936, A2 => n12466, B1 => n12341, B2 => 
                           n9161, ZN => n2271);
   U9055 : OAI22_X1 port map( A1 => n11936, A2 => n12470, B1 => n12341, B2 => 
                           n9160, ZN => n2272);
   U9056 : OAI22_X1 port map( A1 => n11936, A2 => n12474, B1 => n12341, B2 => 
                           n9159, ZN => n2273);
   U9057 : OAI22_X1 port map( A1 => n11936, A2 => n12478, B1 => n12341, B2 => 
                           n9158, ZN => n2274);
   U9058 : OAI22_X1 port map( A1 => n11936, A2 => n12482, B1 => n9873, B2 => 
                           n9157, ZN => n2275);
   U9059 : OAI22_X1 port map( A1 => n11936, A2 => n12486, B1 => n9873, B2 => 
                           n9156, ZN => n2276);
   U9060 : OAI22_X1 port map( A1 => n11936, A2 => n12490, B1 => n9873, B2 => 
                           n9155, ZN => n2277);
   U9061 : OAI22_X1 port map( A1 => n11936, A2 => n12494, B1 => n9873, B2 => 
                           n9154, ZN => n2278);
   U9062 : OAI22_X1 port map( A1 => n11936, A2 => n12498, B1 => n9873, B2 => 
                           n9153, ZN => n2279);
   U9063 : OAI22_X1 port map( A1 => n11936, A2 => n12502, B1 => n9873, B2 => 
                           n9152, ZN => n2280);
   U9064 : OAI22_X1 port map( A1 => n11936, A2 => n12506, B1 => n9873, B2 => 
                           n9151, ZN => n2281);
   U9065 : OAI22_X1 port map( A1 => n11936, A2 => n12514, B1 => n9873, B2 => 
                           n9150, ZN => n2282);
   U9066 : OAI22_X1 port map( A1 => n11965, A2 => n12386, B1 => n12377, B2 => 
                           n8893, ZN => n2539);
   U9067 : OAI22_X1 port map( A1 => n11965, A2 => n12390, B1 => n12377, B2 => 
                           n8892, ZN => n2540);
   U9068 : OAI22_X1 port map( A1 => n11965, A2 => n12394, B1 => n12377, B2 => 
                           n8891, ZN => n2541);
   U9069 : OAI22_X1 port map( A1 => n11965, A2 => n12398, B1 => n12377, B2 => 
                           n8890, ZN => n2542);
   U9070 : OAI22_X1 port map( A1 => n11965, A2 => n12402, B1 => n12377, B2 => 
                           n8889, ZN => n2543);
   U9071 : OAI22_X1 port map( A1 => n11965, A2 => n12406, B1 => n12377, B2 => 
                           n8888, ZN => n2544);
   U9072 : OAI22_X1 port map( A1 => n11965, A2 => n12410, B1 => n12377, B2 => 
                           n8887, ZN => n2545);
   U9073 : OAI22_X1 port map( A1 => n11965, A2 => n12414, B1 => n12377, B2 => 
                           n8886, ZN => n2546);
   U9074 : OAI22_X1 port map( A1 => n11964, A2 => n12418, B1 => n12377, B2 => 
                           n8885, ZN => n2547);
   U9075 : OAI22_X1 port map( A1 => n11964, A2 => n12422, B1 => n12377, B2 => 
                           n8884, ZN => n2548);
   U9076 : OAI22_X1 port map( A1 => n11964, A2 => n12426, B1 => n12377, B2 => 
                           n8883, ZN => n2549);
   U9077 : OAI22_X1 port map( A1 => n11964, A2 => n12430, B1 => n12377, B2 => 
                           n8882, ZN => n2550);
   U9078 : OAI22_X1 port map( A1 => n11964, A2 => n12434, B1 => n9859, B2 => 
                           n8881, ZN => n2551);
   U9079 : OAI22_X1 port map( A1 => n11964, A2 => n12438, B1 => n9859, B2 => 
                           n8880, ZN => n2552);
   U9080 : OAI22_X1 port map( A1 => n11964, A2 => n12442, B1 => n9859, B2 => 
                           n8879, ZN => n2553);
   U9081 : OAI22_X1 port map( A1 => n11964, A2 => n12446, B1 => n12377, B2 => 
                           n8878, ZN => n2554);
   U9082 : OAI22_X1 port map( A1 => n11964, A2 => n12450, B1 => n12377, B2 => 
                           n8877, ZN => n2555);
   U9083 : OAI22_X1 port map( A1 => n11964, A2 => n12454, B1 => n12377, B2 => 
                           n8876, ZN => n2556);
   U9084 : OAI22_X1 port map( A1 => n11964, A2 => n12458, B1 => n12377, B2 => 
                           n8875, ZN => n2557);
   U9085 : OAI22_X1 port map( A1 => n11964, A2 => n12462, B1 => n12377, B2 => 
                           n8874, ZN => n2558);
   U9086 : OAI22_X1 port map( A1 => n11963, A2 => n12466, B1 => n12377, B2 => 
                           n8873, ZN => n2559);
   U9087 : OAI22_X1 port map( A1 => n11963, A2 => n12470, B1 => n12377, B2 => 
                           n8872, ZN => n2560);
   U9088 : OAI22_X1 port map( A1 => n11963, A2 => n12474, B1 => n12377, B2 => 
                           n8871, ZN => n2561);
   U9089 : OAI22_X1 port map( A1 => n11963, A2 => n12478, B1 => n12377, B2 => 
                           n8870, ZN => n2562);
   U9090 : OAI22_X1 port map( A1 => n11963, A2 => n12482, B1 => n9859, B2 => 
                           n8869, ZN => n2563);
   U9091 : OAI22_X1 port map( A1 => n11963, A2 => n12486, B1 => n9859, B2 => 
                           n8868, ZN => n2564);
   U9092 : OAI22_X1 port map( A1 => n11963, A2 => n12490, B1 => n9859, B2 => 
                           n8867, ZN => n2565);
   U9093 : OAI22_X1 port map( A1 => n11963, A2 => n12494, B1 => n9859, B2 => 
                           n8866, ZN => n2566);
   U9094 : OAI22_X1 port map( A1 => n11963, A2 => n12498, B1 => n9859, B2 => 
                           n8865, ZN => n2567);
   U9095 : OAI22_X1 port map( A1 => n11963, A2 => n12502, B1 => n9859, B2 => 
                           n8864, ZN => n2568);
   U9096 : OAI22_X1 port map( A1 => n11963, A2 => n12506, B1 => n9859, B2 => 
                           n8863, ZN => n2569);
   U9097 : OAI22_X1 port map( A1 => n11963, A2 => n12514, B1 => n9859, B2 => 
                           n8862, ZN => n2570);
   U9098 : OAI22_X1 port map( A1 => n11968, A2 => n12386, B1 => n12381, B2 => 
                           n8861, ZN => n2571);
   U9099 : OAI22_X1 port map( A1 => n11968, A2 => n12390, B1 => n12381, B2 => 
                           n8860, ZN => n2572);
   U9100 : OAI22_X1 port map( A1 => n11968, A2 => n12394, B1 => n12381, B2 => 
                           n8859, ZN => n2573);
   U9101 : OAI22_X1 port map( A1 => n11968, A2 => n12398, B1 => n12381, B2 => 
                           n8858, ZN => n2574);
   U9102 : OAI22_X1 port map( A1 => n11968, A2 => n12402, B1 => n12381, B2 => 
                           n8857, ZN => n2575);
   U9103 : OAI22_X1 port map( A1 => n11968, A2 => n12406, B1 => n12381, B2 => 
                           n8856, ZN => n2576);
   U9104 : OAI22_X1 port map( A1 => n11968, A2 => n12410, B1 => n12381, B2 => 
                           n8855, ZN => n2577);
   U9105 : OAI22_X1 port map( A1 => n11968, A2 => n12414, B1 => n12381, B2 => 
                           n8854, ZN => n2578);
   U9106 : OAI22_X1 port map( A1 => n11967, A2 => n12418, B1 => n12381, B2 => 
                           n8853, ZN => n2579);
   U9107 : OAI22_X1 port map( A1 => n11967, A2 => n12422, B1 => n12381, B2 => 
                           n8852, ZN => n2580);
   U9108 : OAI22_X1 port map( A1 => n11967, A2 => n12426, B1 => n12381, B2 => 
                           n8851, ZN => n2581);
   U9109 : OAI22_X1 port map( A1 => n11967, A2 => n12430, B1 => n12381, B2 => 
                           n8850, ZN => n2582);
   U9110 : OAI22_X1 port map( A1 => n11967, A2 => n12434, B1 => n9857, B2 => 
                           n8849, ZN => n2583);
   U9111 : OAI22_X1 port map( A1 => n11967, A2 => n12438, B1 => n9857, B2 => 
                           n8848, ZN => n2584);
   U9112 : OAI22_X1 port map( A1 => n11967, A2 => n12442, B1 => n9857, B2 => 
                           n8847, ZN => n2585);
   U9113 : OAI22_X1 port map( A1 => n11967, A2 => n12446, B1 => n12381, B2 => 
                           n8846, ZN => n2586);
   U9114 : OAI22_X1 port map( A1 => n11967, A2 => n12450, B1 => n12381, B2 => 
                           n8845, ZN => n2587);
   U9115 : OAI22_X1 port map( A1 => n11967, A2 => n12454, B1 => n12381, B2 => 
                           n8844, ZN => n2588);
   U9116 : OAI22_X1 port map( A1 => n11967, A2 => n12458, B1 => n12381, B2 => 
                           n8843, ZN => n2589);
   U9117 : OAI22_X1 port map( A1 => n11967, A2 => n12462, B1 => n12381, B2 => 
                           n8842, ZN => n2590);
   U9118 : OAI22_X1 port map( A1 => n11966, A2 => n12466, B1 => n12381, B2 => 
                           n8841, ZN => n2591);
   U9119 : OAI22_X1 port map( A1 => n11966, A2 => n12470, B1 => n12381, B2 => 
                           n8840, ZN => n2592);
   U9120 : OAI22_X1 port map( A1 => n11966, A2 => n12474, B1 => n12381, B2 => 
                           n8839, ZN => n2593);
   U9121 : OAI22_X1 port map( A1 => n11966, A2 => n12478, B1 => n12381, B2 => 
                           n8838, ZN => n2594);
   U9122 : OAI22_X1 port map( A1 => n11966, A2 => n12482, B1 => n9857, B2 => 
                           n8837, ZN => n2595);
   U9123 : OAI22_X1 port map( A1 => n11966, A2 => n12486, B1 => n9857, B2 => 
                           n8836, ZN => n2596);
   U9124 : OAI22_X1 port map( A1 => n11966, A2 => n12490, B1 => n9857, B2 => 
                           n8835, ZN => n2597);
   U9125 : OAI22_X1 port map( A1 => n11966, A2 => n12494, B1 => n9857, B2 => 
                           n8834, ZN => n2598);
   U9126 : OAI22_X1 port map( A1 => n11966, A2 => n12498, B1 => n9857, B2 => 
                           n8833, ZN => n2599);
   U9127 : OAI22_X1 port map( A1 => n11966, A2 => n12502, B1 => n9857, B2 => 
                           n8832, ZN => n2600);
   U9128 : OAI22_X1 port map( A1 => n11966, A2 => n12506, B1 => n9857, B2 => 
                           n8831, ZN => n2601);
   U9129 : OAI22_X1 port map( A1 => n11966, A2 => n12514, B1 => n9857, B2 => 
                           n8830, ZN => n2602);
   U9130 : OAI22_X1 port map( A1 => n11887, A2 => n12388, B1 => n12273, B2 => 
                           n9725, ZN => n1707);
   U9131 : OAI22_X1 port map( A1 => n11887, A2 => n12392, B1 => n12273, B2 => 
                           n9724, ZN => n1708);
   U9132 : OAI22_X1 port map( A1 => n11887, A2 => n12396, B1 => n12273, B2 => 
                           n9723, ZN => n1709);
   U9133 : OAI22_X1 port map( A1 => n11887, A2 => n12400, B1 => n12273, B2 => 
                           n9722, ZN => n1710);
   U9134 : OAI22_X1 port map( A1 => n11887, A2 => n12404, B1 => n12273, B2 => 
                           n9721, ZN => n1711);
   U9135 : OAI22_X1 port map( A1 => n11887, A2 => n12408, B1 => n12273, B2 => 
                           n9720, ZN => n1712);
   U9136 : OAI22_X1 port map( A1 => n11887, A2 => n12412, B1 => n12273, B2 => 
                           n9719, ZN => n1713);
   U9137 : OAI22_X1 port map( A1 => n11887, A2 => n12416, B1 => n12273, B2 => 
                           n9718, ZN => n1714);
   U9138 : OAI22_X1 port map( A1 => n11886, A2 => n12420, B1 => n12273, B2 => 
                           n9717, ZN => n1715);
   U9139 : OAI22_X1 port map( A1 => n11886, A2 => n12424, B1 => n12273, B2 => 
                           n9716, ZN => n1716);
   U9140 : OAI22_X1 port map( A1 => n11886, A2 => n12428, B1 => n12273, B2 => 
                           n9715, ZN => n1717);
   U9141 : OAI22_X1 port map( A1 => n11886, A2 => n12432, B1 => n12273, B2 => 
                           n9714, ZN => n1718);
   U9142 : OAI22_X1 port map( A1 => n11886, A2 => n12436, B1 => n9895, B2 => 
                           n9713, ZN => n1719);
   U9143 : OAI22_X1 port map( A1 => n11886, A2 => n12440, B1 => n9895, B2 => 
                           n9712, ZN => n1720);
   U9144 : OAI22_X1 port map( A1 => n11886, A2 => n12444, B1 => n9895, B2 => 
                           n9711, ZN => n1721);
   U9145 : OAI22_X1 port map( A1 => n11886, A2 => n12448, B1 => n12273, B2 => 
                           n9710, ZN => n1722);
   U9146 : OAI22_X1 port map( A1 => n11886, A2 => n12452, B1 => n12273, B2 => 
                           n9709, ZN => n1723);
   U9147 : OAI22_X1 port map( A1 => n11886, A2 => n12456, B1 => n12273, B2 => 
                           n9708, ZN => n1724);
   U9148 : OAI22_X1 port map( A1 => n11886, A2 => n12460, B1 => n12273, B2 => 
                           n9707, ZN => n1725);
   U9149 : OAI22_X1 port map( A1 => n11886, A2 => n12464, B1 => n12273, B2 => 
                           n9706, ZN => n1726);
   U9150 : OAI22_X1 port map( A1 => n11885, A2 => n12468, B1 => n12273, B2 => 
                           n9705, ZN => n1727);
   U9151 : OAI22_X1 port map( A1 => n11885, A2 => n12472, B1 => n12273, B2 => 
                           n9704, ZN => n1728);
   U9152 : OAI22_X1 port map( A1 => n11885, A2 => n12476, B1 => n12273, B2 => 
                           n9703, ZN => n1729);
   U9153 : OAI22_X1 port map( A1 => n11885, A2 => n12480, B1 => n12273, B2 => 
                           n9702, ZN => n1730);
   U9154 : OAI22_X1 port map( A1 => n11885, A2 => n12484, B1 => n9895, B2 => 
                           n9701, ZN => n1731);
   U9155 : OAI22_X1 port map( A1 => n11885, A2 => n12488, B1 => n9895, B2 => 
                           n9700, ZN => n1732);
   U9156 : OAI22_X1 port map( A1 => n11885, A2 => n12492, B1 => n9895, B2 => 
                           n9699, ZN => n1733);
   U9157 : OAI22_X1 port map( A1 => n11885, A2 => n12496, B1 => n9895, B2 => 
                           n9698, ZN => n1734);
   U9158 : OAI22_X1 port map( A1 => n11885, A2 => n12500, B1 => n9895, B2 => 
                           n9697, ZN => n1735);
   U9159 : OAI22_X1 port map( A1 => n11885, A2 => n12504, B1 => n9895, B2 => 
                           n9696, ZN => n1736);
   U9160 : OAI22_X1 port map( A1 => n11885, A2 => n12508, B1 => n9895, B2 => 
                           n9695, ZN => n1737);
   U9161 : OAI22_X1 port map( A1 => n11885, A2 => n12516, B1 => n9895, B2 => 
                           n9694, ZN => n1738);
   U9162 : OAI22_X1 port map( A1 => n11899, A2 => n12388, B1 => n12289, B2 => 
                           n9597, ZN => n1835);
   U9163 : OAI22_X1 port map( A1 => n11899, A2 => n12392, B1 => n12289, B2 => 
                           n9596, ZN => n1836);
   U9164 : OAI22_X1 port map( A1 => n11899, A2 => n12396, B1 => n12289, B2 => 
                           n9595, ZN => n1837);
   U9165 : OAI22_X1 port map( A1 => n11899, A2 => n12400, B1 => n12289, B2 => 
                           n9594, ZN => n1838);
   U9166 : OAI22_X1 port map( A1 => n11899, A2 => n12404, B1 => n12289, B2 => 
                           n9593, ZN => n1839);
   U9167 : OAI22_X1 port map( A1 => n11899, A2 => n12408, B1 => n12289, B2 => 
                           n9592, ZN => n1840);
   U9168 : OAI22_X1 port map( A1 => n11899, A2 => n12412, B1 => n12289, B2 => 
                           n9591, ZN => n1841);
   U9169 : OAI22_X1 port map( A1 => n11899, A2 => n12416, B1 => n12289, B2 => 
                           n9590, ZN => n1842);
   U9170 : OAI22_X1 port map( A1 => n11898, A2 => n12420, B1 => n12289, B2 => 
                           n9589, ZN => n1843);
   U9171 : OAI22_X1 port map( A1 => n11898, A2 => n12424, B1 => n12289, B2 => 
                           n9588, ZN => n1844);
   U9172 : OAI22_X1 port map( A1 => n11898, A2 => n12428, B1 => n12289, B2 => 
                           n9587, ZN => n1845);
   U9173 : OAI22_X1 port map( A1 => n11898, A2 => n12432, B1 => n12289, B2 => 
                           n9586, ZN => n1846);
   U9174 : OAI22_X1 port map( A1 => n11898, A2 => n12436, B1 => n9890, B2 => 
                           n9585, ZN => n1847);
   U9175 : OAI22_X1 port map( A1 => n11898, A2 => n12440, B1 => n9890, B2 => 
                           n9584, ZN => n1848);
   U9176 : OAI22_X1 port map( A1 => n11898, A2 => n12444, B1 => n9890, B2 => 
                           n9583, ZN => n1849);
   U9177 : OAI22_X1 port map( A1 => n11898, A2 => n12448, B1 => n12289, B2 => 
                           n9582, ZN => n1850);
   U9178 : OAI22_X1 port map( A1 => n11898, A2 => n12452, B1 => n12289, B2 => 
                           n9581, ZN => n1851);
   U9179 : OAI22_X1 port map( A1 => n11898, A2 => n12456, B1 => n12289, B2 => 
                           n9580, ZN => n1852);
   U9180 : OAI22_X1 port map( A1 => n11898, A2 => n12460, B1 => n12289, B2 => 
                           n9579, ZN => n1853);
   U9181 : OAI22_X1 port map( A1 => n11898, A2 => n12464, B1 => n12289, B2 => 
                           n9578, ZN => n1854);
   U9182 : OAI22_X1 port map( A1 => n11897, A2 => n12468, B1 => n12289, B2 => 
                           n9577, ZN => n1855);
   U9183 : OAI22_X1 port map( A1 => n11897, A2 => n12472, B1 => n12289, B2 => 
                           n9576, ZN => n1856);
   U9184 : OAI22_X1 port map( A1 => n11897, A2 => n12476, B1 => n12289, B2 => 
                           n9575, ZN => n1857);
   U9185 : OAI22_X1 port map( A1 => n11897, A2 => n12480, B1 => n12289, B2 => 
                           n9574, ZN => n1858);
   U9186 : OAI22_X1 port map( A1 => n11897, A2 => n12484, B1 => n9890, B2 => 
                           n9573, ZN => n1859);
   U9187 : OAI22_X1 port map( A1 => n11897, A2 => n12488, B1 => n9890, B2 => 
                           n9572, ZN => n1860);
   U9188 : OAI22_X1 port map( A1 => n11897, A2 => n12492, B1 => n9890, B2 => 
                           n9571, ZN => n1861);
   U9189 : OAI22_X1 port map( A1 => n11897, A2 => n12496, B1 => n9890, B2 => 
                           n9570, ZN => n1862);
   U9190 : OAI22_X1 port map( A1 => n11897, A2 => n12500, B1 => n9890, B2 => 
                           n9569, ZN => n1863);
   U9191 : OAI22_X1 port map( A1 => n11897, A2 => n12504, B1 => n9890, B2 => 
                           n9568, ZN => n1864);
   U9192 : OAI22_X1 port map( A1 => n11897, A2 => n12508, B1 => n9890, B2 => 
                           n9567, ZN => n1865);
   U9193 : OAI22_X1 port map( A1 => n11897, A2 => n12516, B1 => n9890, B2 => 
                           n9566, ZN => n1866);
   U9194 : OAI22_X1 port map( A1 => n11917, A2 => n12387, B1 => n12313, B2 => 
                           n9405, ZN => n2027);
   U9195 : OAI22_X1 port map( A1 => n11917, A2 => n12391, B1 => n12313, B2 => 
                           n9404, ZN => n2028);
   U9196 : OAI22_X1 port map( A1 => n11917, A2 => n12395, B1 => n12313, B2 => 
                           n9403, ZN => n2029);
   U9197 : OAI22_X1 port map( A1 => n11917, A2 => n12399, B1 => n12313, B2 => 
                           n9402, ZN => n2030);
   U9198 : OAI22_X1 port map( A1 => n11917, A2 => n12403, B1 => n12313, B2 => 
                           n9401, ZN => n2031);
   U9199 : OAI22_X1 port map( A1 => n11917, A2 => n12407, B1 => n12313, B2 => 
                           n9400, ZN => n2032);
   U9200 : OAI22_X1 port map( A1 => n11917, A2 => n12411, B1 => n12313, B2 => 
                           n9399, ZN => n2033);
   U9201 : OAI22_X1 port map( A1 => n11917, A2 => n12415, B1 => n12313, B2 => 
                           n9398, ZN => n2034);
   U9202 : OAI22_X1 port map( A1 => n11916, A2 => n12419, B1 => n12313, B2 => 
                           n9397, ZN => n2035);
   U9203 : OAI22_X1 port map( A1 => n11916, A2 => n12423, B1 => n12313, B2 => 
                           n9396, ZN => n2036);
   U9204 : OAI22_X1 port map( A1 => n11916, A2 => n12427, B1 => n12313, B2 => 
                           n9395, ZN => n2037);
   U9205 : OAI22_X1 port map( A1 => n11916, A2 => n12431, B1 => n12313, B2 => 
                           n9394, ZN => n2038);
   U9206 : OAI22_X1 port map( A1 => n11916, A2 => n12435, B1 => n9882, B2 => 
                           n9393, ZN => n2039);
   U9207 : OAI22_X1 port map( A1 => n11916, A2 => n12439, B1 => n9882, B2 => 
                           n9392, ZN => n2040);
   U9208 : OAI22_X1 port map( A1 => n11916, A2 => n12443, B1 => n9882, B2 => 
                           n9391, ZN => n2041);
   U9209 : OAI22_X1 port map( A1 => n11916, A2 => n12447, B1 => n12313, B2 => 
                           n9390, ZN => n2042);
   U9210 : OAI22_X1 port map( A1 => n11916, A2 => n12451, B1 => n12313, B2 => 
                           n9389, ZN => n2043);
   U9211 : OAI22_X1 port map( A1 => n11916, A2 => n12455, B1 => n12313, B2 => 
                           n9388, ZN => n2044);
   U9212 : OAI22_X1 port map( A1 => n11916, A2 => n12459, B1 => n12313, B2 => 
                           n9387, ZN => n2045);
   U9213 : OAI22_X1 port map( A1 => n11916, A2 => n12463, B1 => n12313, B2 => 
                           n9386, ZN => n2046);
   U9214 : OAI22_X1 port map( A1 => n11915, A2 => n12467, B1 => n12313, B2 => 
                           n9385, ZN => n2047);
   U9215 : OAI22_X1 port map( A1 => n11915, A2 => n12471, B1 => n12313, B2 => 
                           n9384, ZN => n2048);
   U9216 : OAI22_X1 port map( A1 => n11915, A2 => n12475, B1 => n12313, B2 => 
                           n9383, ZN => n2049);
   U9217 : OAI22_X1 port map( A1 => n11915, A2 => n12479, B1 => n12313, B2 => 
                           n9382, ZN => n2050);
   U9218 : OAI22_X1 port map( A1 => n11915, A2 => n12483, B1 => n9882, B2 => 
                           n9381, ZN => n2051);
   U9219 : OAI22_X1 port map( A1 => n11915, A2 => n12487, B1 => n9882, B2 => 
                           n9380, ZN => n2052);
   U9220 : OAI22_X1 port map( A1 => n11915, A2 => n12491, B1 => n9882, B2 => 
                           n9379, ZN => n2053);
   U9221 : OAI22_X1 port map( A1 => n11915, A2 => n12495, B1 => n9882, B2 => 
                           n9378, ZN => n2054);
   U9222 : OAI22_X1 port map( A1 => n11915, A2 => n12499, B1 => n9882, B2 => 
                           n9377, ZN => n2055);
   U9223 : OAI22_X1 port map( A1 => n11915, A2 => n12503, B1 => n9882, B2 => 
                           n9376, ZN => n2056);
   U9224 : OAI22_X1 port map( A1 => n11915, A2 => n12507, B1 => n9882, B2 => 
                           n9375, ZN => n2057);
   U9225 : OAI22_X1 port map( A1 => n11915, A2 => n12515, B1 => n9882, B2 => 
                           n9374, ZN => n2058);
   U9226 : NOR3_X1 port map( A1 => n8795, A2 => n8796, A3 => n8797, ZN => 
                           n11078);
   U9227 : NOR3_X1 port map( A1 => n8791, A2 => n8792, A3 => n8793, ZN => 
                           n10478);
   U9228 : NAND2_X1 port map( A1 => n8786, A2 => n8789, ZN => n9856);
   U9229 : NOR3_X1 port map( A1 => n11086, A2 => n8783, A3 => n11087, ZN => 
                           n11085);
   U9230 : NOR3_X1 port map( A1 => n10486, A2 => n8783, A3 => n10487, ZN => 
                           n10485);
   U9231 : NAND2_X1 port map( A1 => n11094, A2 => n11072, ZN => n10536);
   U9232 : NAND2_X1 port map( A1 => n11095, A2 => n11072, ZN => n10535);
   U9233 : NAND2_X1 port map( A1 => n11095, A2 => n11073, ZN => n10547);
   U9234 : NAND2_X1 port map( A1 => n11094, A2 => n11078, ZN => n10546);
   U9235 : NAND2_X1 port map( A1 => n11094, A2 => n11069, ZN => n10531);
   U9236 : NAND2_X1 port map( A1 => n11095, A2 => n11069, ZN => n10530);
   U9237 : NAND2_X1 port map( A1 => n11095, A2 => n11075, ZN => n10542);
   U9238 : NAND2_X1 port map( A1 => n11094, A2 => n11071, ZN => n10541);
   U9239 : NAND2_X1 port map( A1 => n10494, A2 => n10472, ZN => n9936);
   U9240 : NAND2_X1 port map( A1 => n10495, A2 => n10472, ZN => n9935);
   U9241 : NAND2_X1 port map( A1 => n10495, A2 => n10473, ZN => n9947);
   U9242 : NAND2_X1 port map( A1 => n10494, A2 => n10478, ZN => n9946);
   U9243 : NAND2_X1 port map( A1 => n10494, A2 => n10469, ZN => n9931);
   U9244 : NAND2_X1 port map( A1 => n10495, A2 => n10469, ZN => n9930);
   U9245 : NAND2_X1 port map( A1 => n10495, A2 => n10475, ZN => n9942);
   U9246 : NAND2_X1 port map( A1 => n10494, A2 => n10471, ZN => n9941);
   U9247 : AND3_X1 port map( A1 => n11068, A2 => n12055, A3 => n11072, ZN => 
                           n10505);
   U9248 : AND3_X1 port map( A1 => n11073, A2 => n12055, A3 => n11077, ZN => 
                           n10511);
   U9249 : AND3_X1 port map( A1 => n11072, A2 => n12055, A3 => n11077, ZN => 
                           n10516);
   U9250 : AND3_X1 port map( A1 => n10468, A2 => n12199, A3 => n10472, ZN => 
                           n9905);
   U9251 : AND3_X1 port map( A1 => n10473, A2 => n12199, A3 => n10477, ZN => 
                           n9911);
   U9252 : AND3_X1 port map( A1 => n10472, A2 => n12199, A3 => n10477, ZN => 
                           n9916);
   U9253 : AND3_X1 port map( A1 => n11068, A2 => n12055, A3 => n11073, ZN => 
                           n10504);
   U9254 : AND3_X1 port map( A1 => n11077, A2 => n12055, A3 => n11078, ZN => 
                           n10510);
   U9255 : AND3_X1 port map( A1 => n11070, A2 => n12055, A3 => n11077, ZN => 
                           n10515);
   U9256 : AND3_X1 port map( A1 => n10468, A2 => n12199, A3 => n10473, ZN => 
                           n9904);
   U9257 : AND3_X1 port map( A1 => n10477, A2 => n12199, A3 => n10478, ZN => 
                           n9910);
   U9258 : AND3_X1 port map( A1 => n10470, A2 => n12199, A3 => n10477, ZN => 
                           n9915);
   U9259 : AND2_X1 port map( A1 => n11094, A2 => n11075, ZN => n10539);
   U9260 : AND2_X1 port map( A1 => n11095, A2 => n11070, ZN => n10540);
   U9261 : AND2_X1 port map( A1 => n11094, A2 => n11070, ZN => n10538);
   U9262 : AND2_X1 port map( A1 => n11095, A2 => n11076, ZN => n10550);
   U9263 : AND2_X1 port map( A1 => n11094, A2 => n11076, ZN => n10551);
   U9264 : AND2_X1 port map( A1 => n11095, A2 => n11078, ZN => n10549);
   U9265 : AND2_X1 port map( A1 => n11095, A2 => n11071, ZN => n10545);
   U9266 : AND2_X1 port map( A1 => n11094, A2 => n11073, ZN => n10544);
   U9267 : AND2_X1 port map( A1 => n10494, A2 => n10475, ZN => n9939);
   U9268 : AND2_X1 port map( A1 => n10495, A2 => n10470, ZN => n9940);
   U9269 : AND2_X1 port map( A1 => n10494, A2 => n10470, ZN => n9938);
   U9270 : AND2_X1 port map( A1 => n10495, A2 => n10476, ZN => n9950);
   U9271 : AND2_X1 port map( A1 => n10494, A2 => n10476, ZN => n9951);
   U9272 : AND2_X1 port map( A1 => n10495, A2 => n10478, ZN => n9949);
   U9273 : AND2_X1 port map( A1 => n10495, A2 => n10471, ZN => n9945);
   U9274 : AND2_X1 port map( A1 => n10494, A2 => n10473, ZN => n9944);
   U9275 : AND2_X1 port map( A1 => n11078, A2 => n11068, ZN => n10534);
   U9276 : AND2_X1 port map( A1 => n11076, A2 => n11068, ZN => n10533);
   U9277 : AND2_X1 port map( A1 => n10478, A2 => n10468, ZN => n9934);
   U9278 : AND2_X1 port map( A1 => n10476, A2 => n10468, ZN => n9933);
   U9279 : AND4_X1 port map( A1 => n11084, A2 => n11083, A3 => n11870, A4 => 
                           n11099, ZN => n10520);
   U9280 : NOR4_X1 port map( A1 => n8783, A2 => n11087, A3 => n11086, A4 => 
                           n11088, ZN => n11099);
   U9281 : AND4_X1 port map( A1 => n10484, A2 => n10483, A3 => n11873, A4 => 
                           n10499, ZN => n9920);
   U9282 : NOR4_X1 port map( A1 => n8783, A2 => n10487, A3 => n10486, A4 => 
                           n10488, ZN => n10499);
   U9283 : BUF_X1 port map( A => n9899, Z => n12264);
   U9284 : OAI21_X1 port map( B1 => n9862, B2 => n9896, A => n12519, ZN => 
                           n9899);
   U9285 : INV_X1 port map( A => n9898, ZN => n12268);
   U9286 : OAI21_X1 port map( B1 => n9860, B2 => n9896, A => n12520, ZN => 
                           n9898);
   U9287 : INV_X1 port map( A => n9897, ZN => n12272);
   U9288 : OAI21_X1 port map( B1 => n9858, B2 => n9896, A => n12520, ZN => 
                           n9897);
   U9289 : INV_X1 port map( A => n9895, ZN => n12276);
   U9290 : OAI21_X1 port map( B1 => n9856, B2 => n9896, A => n12520, ZN => 
                           n9895);
   U9291 : INV_X1 port map( A => n9894, ZN => n12280);
   U9292 : OAI21_X1 port map( B1 => n9862, B2 => n9891, A => n12520, ZN => 
                           n9894);
   U9293 : INV_X1 port map( A => n9893, ZN => n12284);
   U9294 : OAI21_X1 port map( B1 => n9860, B2 => n9891, A => n12520, ZN => 
                           n9893);
   U9295 : INV_X1 port map( A => n9892, ZN => n12288);
   U9296 : OAI21_X1 port map( B1 => n9858, B2 => n9891, A => n12520, ZN => 
                           n9892);
   U9297 : INV_X1 port map( A => n9890, ZN => n12292);
   U9298 : OAI21_X1 port map( B1 => n9856, B2 => n9891, A => n12520, ZN => 
                           n9890);
   U9299 : INV_X1 port map( A => n9889, ZN => n12296);
   U9300 : OAI21_X1 port map( B1 => n9862, B2 => n9886, A => n12520, ZN => 
                           n9889);
   U9301 : INV_X1 port map( A => n9888, ZN => n12300);
   U9302 : OAI21_X1 port map( B1 => n9860, B2 => n9886, A => n12520, ZN => 
                           n9888);
   U9303 : INV_X1 port map( A => n9887, ZN => n12304);
   U9304 : OAI21_X1 port map( B1 => n9858, B2 => n9886, A => n12522, ZN => 
                           n9887);
   U9305 : INV_X1 port map( A => n9885, ZN => n12308);
   U9306 : OAI21_X1 port map( B1 => n9856, B2 => n9886, A => n12520, ZN => 
                           n9885);
   U9307 : INV_X1 port map( A => n9883, ZN => n12312);
   U9308 : OAI21_X1 port map( B1 => n9862, B2 => n9880, A => n12520, ZN => 
                           n9883);
   U9309 : INV_X1 port map( A => n9882, ZN => n12316);
   U9310 : OAI21_X1 port map( B1 => n9860, B2 => n9880, A => n12520, ZN => 
                           n9882);
   U9311 : INV_X1 port map( A => n9881, ZN => n12320);
   U9312 : OAI21_X1 port map( B1 => n9858, B2 => n9880, A => n12520, ZN => 
                           n9881);
   U9313 : INV_X1 port map( A => n9878, ZN => n12328);
   U9314 : OAI21_X1 port map( B1 => n9862, B2 => n9875, A => n12521, ZN => 
                           n9878);
   U9315 : INV_X1 port map( A => n9877, ZN => n12332);
   U9316 : OAI21_X1 port map( B1 => n9860, B2 => n9875, A => n12521, ZN => 
                           n9877);
   U9317 : INV_X1 port map( A => n9876, ZN => n12336);
   U9318 : OAI21_X1 port map( B1 => n9858, B2 => n9875, A => n12521, ZN => 
                           n9876);
   U9319 : INV_X1 port map( A => n9874, ZN => n12340);
   U9320 : OAI21_X1 port map( B1 => n9856, B2 => n9875, A => n12521, ZN => 
                           n9874);
   U9321 : INV_X1 port map( A => n9873, ZN => n12344);
   U9322 : OAI21_X1 port map( B1 => n9862, B2 => n9870, A => n12521, ZN => 
                           n9873);
   U9323 : INV_X1 port map( A => n9872, ZN => n12348);
   U9324 : OAI21_X1 port map( B1 => n9860, B2 => n9870, A => n12521, ZN => 
                           n9872);
   U9325 : INV_X1 port map( A => n9871, ZN => n12352);
   U9326 : OAI21_X1 port map( B1 => n9858, B2 => n9870, A => n12521, ZN => 
                           n9871);
   U9327 : INV_X1 port map( A => n9869, ZN => n12356);
   U9328 : OAI21_X1 port map( B1 => n9856, B2 => n9870, A => n12521, ZN => 
                           n9869);
   U9329 : INV_X1 port map( A => n9868, ZN => n12360);
   U9330 : OAI21_X1 port map( B1 => n9862, B2 => n9865, A => n12521, ZN => 
                           n9868);
   U9331 : INV_X1 port map( A => n9867, ZN => n12364);
   U9332 : OAI21_X1 port map( B1 => n9860, B2 => n9865, A => n12521, ZN => 
                           n9867);
   U9333 : INV_X1 port map( A => n9866, ZN => n12368);
   U9334 : OAI21_X1 port map( B1 => n9858, B2 => n9865, A => n12521, ZN => 
                           n9866);
   U9335 : INV_X1 port map( A => n9864, ZN => n12372);
   U9336 : OAI21_X1 port map( B1 => n9856, B2 => n9865, A => n12521, ZN => 
                           n9864);
   U9337 : INV_X1 port map( A => n9861, ZN => n12376);
   U9338 : OAI21_X1 port map( B1 => n9855, B2 => n9862, A => n12522, ZN => 
                           n9861);
   U9339 : INV_X1 port map( A => n9859, ZN => n12380);
   U9340 : OAI21_X1 port map( B1 => n9855, B2 => n9860, A => n12522, ZN => 
                           n9859);
   U9341 : INV_X1 port map( A => n9857, ZN => n12384);
   U9342 : OAI21_X1 port map( B1 => n9855, B2 => n9858, A => n12522, ZN => 
                           n9857);
   U9343 : BUF_X1 port map( A => n12385, Z => n12387);
   U9344 : BUF_X1 port map( A => n12389, Z => n12391);
   U9345 : BUF_X1 port map( A => n12393, Z => n12395);
   U9346 : BUF_X1 port map( A => n12397, Z => n12399);
   U9347 : BUF_X1 port map( A => n12401, Z => n12403);
   U9348 : BUF_X1 port map( A => n12405, Z => n12407);
   U9349 : BUF_X1 port map( A => n12409, Z => n12411);
   U9350 : BUF_X1 port map( A => n12413, Z => n12415);
   U9351 : BUF_X1 port map( A => n12417, Z => n12419);
   U9352 : BUF_X1 port map( A => n12421, Z => n12423);
   U9353 : BUF_X1 port map( A => n12425, Z => n12427);
   U9354 : BUF_X1 port map( A => n12429, Z => n12431);
   U9355 : BUF_X1 port map( A => n12433, Z => n12435);
   U9356 : BUF_X1 port map( A => n12437, Z => n12439);
   U9357 : BUF_X1 port map( A => n12441, Z => n12443);
   U9358 : BUF_X1 port map( A => n12445, Z => n12447);
   U9359 : BUF_X1 port map( A => n12449, Z => n12451);
   U9360 : BUF_X1 port map( A => n12453, Z => n12455);
   U9361 : BUF_X1 port map( A => n12457, Z => n12459);
   U9362 : BUF_X1 port map( A => n12461, Z => n12463);
   U9363 : BUF_X1 port map( A => n12465, Z => n12467);
   U9364 : BUF_X1 port map( A => n12469, Z => n12471);
   U9365 : BUF_X1 port map( A => n12473, Z => n12475);
   U9366 : BUF_X1 port map( A => n12477, Z => n12479);
   U9367 : BUF_X1 port map( A => n12481, Z => n12483);
   U9368 : BUF_X1 port map( A => n12485, Z => n12487);
   U9369 : BUF_X1 port map( A => n12489, Z => n12491);
   U9370 : BUF_X1 port map( A => n12493, Z => n12495);
   U9371 : BUF_X1 port map( A => n12497, Z => n12499);
   U9372 : BUF_X1 port map( A => n12501, Z => n12503);
   U9373 : BUF_X1 port map( A => n12505, Z => n12507);
   U9374 : BUF_X1 port map( A => n12513, Z => n12515);
   U9375 : BUF_X1 port map( A => n12385, Z => n12386);
   U9376 : BUF_X1 port map( A => n12389, Z => n12390);
   U9377 : BUF_X1 port map( A => n12393, Z => n12394);
   U9378 : BUF_X1 port map( A => n12397, Z => n12398);
   U9379 : BUF_X1 port map( A => n12401, Z => n12402);
   U9380 : BUF_X1 port map( A => n12405, Z => n12406);
   U9381 : BUF_X1 port map( A => n12409, Z => n12410);
   U9382 : BUF_X1 port map( A => n12413, Z => n12414);
   U9383 : BUF_X1 port map( A => n12417, Z => n12418);
   U9384 : BUF_X1 port map( A => n12421, Z => n12422);
   U9385 : BUF_X1 port map( A => n12425, Z => n12426);
   U9386 : BUF_X1 port map( A => n12429, Z => n12430);
   U9387 : BUF_X1 port map( A => n12433, Z => n12434);
   U9388 : BUF_X1 port map( A => n12437, Z => n12438);
   U9389 : BUF_X1 port map( A => n12441, Z => n12442);
   U9390 : BUF_X1 port map( A => n12445, Z => n12446);
   U9391 : BUF_X1 port map( A => n12449, Z => n12450);
   U9392 : BUF_X1 port map( A => n12453, Z => n12454);
   U9393 : BUF_X1 port map( A => n12457, Z => n12458);
   U9394 : BUF_X1 port map( A => n12461, Z => n12462);
   U9395 : BUF_X1 port map( A => n12465, Z => n12466);
   U9396 : BUF_X1 port map( A => n12469, Z => n12470);
   U9397 : BUF_X1 port map( A => n12473, Z => n12474);
   U9398 : BUF_X1 port map( A => n12477, Z => n12478);
   U9399 : BUF_X1 port map( A => n12481, Z => n12482);
   U9400 : BUF_X1 port map( A => n12485, Z => n12486);
   U9401 : BUF_X1 port map( A => n12489, Z => n12490);
   U9402 : BUF_X1 port map( A => n12493, Z => n12494);
   U9403 : BUF_X1 port map( A => n12497, Z => n12498);
   U9404 : BUF_X1 port map( A => n12501, Z => n12502);
   U9405 : BUF_X1 port map( A => n12505, Z => n12506);
   U9406 : BUF_X1 port map( A => n12513, Z => n12514);
   U9407 : BUF_X1 port map( A => n11972, Z => n11973);
   U9408 : BUF_X1 port map( A => n11972, Z => n11974);
   U9409 : BUF_X1 port map( A => n12116, Z => n12117);
   U9410 : BUF_X1 port map( A => n12116, Z => n12118);
   U9411 : BUF_X1 port map( A => n11868, Z => n12055);
   U9412 : BUF_X1 port map( A => n11869, Z => n12199);
   U9413 : BUF_X1 port map( A => n12385, Z => n12388);
   U9414 : BUF_X1 port map( A => n12389, Z => n12392);
   U9415 : BUF_X1 port map( A => n12393, Z => n12396);
   U9416 : BUF_X1 port map( A => n12397, Z => n12400);
   U9417 : BUF_X1 port map( A => n12401, Z => n12404);
   U9418 : BUF_X1 port map( A => n12405, Z => n12408);
   U9419 : BUF_X1 port map( A => n12409, Z => n12412);
   U9420 : BUF_X1 port map( A => n12413, Z => n12416);
   U9421 : BUF_X1 port map( A => n12417, Z => n12420);
   U9422 : BUF_X1 port map( A => n12421, Z => n12424);
   U9423 : BUF_X1 port map( A => n12425, Z => n12428);
   U9424 : BUF_X1 port map( A => n12429, Z => n12432);
   U9425 : BUF_X1 port map( A => n12433, Z => n12436);
   U9426 : BUF_X1 port map( A => n12437, Z => n12440);
   U9427 : BUF_X1 port map( A => n12441, Z => n12444);
   U9428 : BUF_X1 port map( A => n12445, Z => n12448);
   U9429 : BUF_X1 port map( A => n12449, Z => n12452);
   U9430 : BUF_X1 port map( A => n12453, Z => n12456);
   U9431 : BUF_X1 port map( A => n12457, Z => n12460);
   U9432 : BUF_X1 port map( A => n12461, Z => n12464);
   U9433 : BUF_X1 port map( A => n12465, Z => n12468);
   U9434 : BUF_X1 port map( A => n12469, Z => n12472);
   U9435 : BUF_X1 port map( A => n12473, Z => n12476);
   U9436 : BUF_X1 port map( A => n12477, Z => n12480);
   U9437 : BUF_X1 port map( A => n12481, Z => n12484);
   U9438 : BUF_X1 port map( A => n12485, Z => n12488);
   U9439 : BUF_X1 port map( A => n12489, Z => n12492);
   U9440 : BUF_X1 port map( A => n12493, Z => n12496);
   U9441 : BUF_X1 port map( A => n12497, Z => n12500);
   U9442 : BUF_X1 port map( A => n12501, Z => n12504);
   U9443 : BUF_X1 port map( A => n12505, Z => n12508);
   U9444 : BUF_X1 port map( A => n12513, Z => n12516);
   U9445 : BUF_X1 port map( A => n11972, Z => n11975);
   U9446 : BUF_X1 port map( A => n12116, Z => n12119);
   U9447 : OAI221_X1 port map( B1 => n8925, B2 => n12029, C1 => n9181, C2 => 
                           n12025, A => n11096, ZN => n11091);
   U9448 : AOI222_X1 port map( A1 => n12021, A2 => n11613, B1 => n12018, B2 => 
                           n11677, C1 => n12014, C2 => n11741, ZN => n11096);
   U9449 : OAI221_X1 port map( B1 => n8924, B2 => n12029, C1 => n9180, C2 => 
                           n12025, A => n11060, ZN => n11057);
   U9450 : AOI222_X1 port map( A1 => n12021, A2 => n11614, B1 => n12018, B2 => 
                           n11678, C1 => n12014, C2 => n11742, ZN => n11060);
   U9451 : OAI221_X1 port map( B1 => n8923, B2 => n12029, C1 => n9179, C2 => 
                           n12025, A => n11043, ZN => n11040);
   U9452 : AOI222_X1 port map( A1 => n12021, A2 => n11615, B1 => n12018, B2 => 
                           n11679, C1 => n12014, C2 => n11743, ZN => n11043);
   U9453 : OAI221_X1 port map( B1 => n8922, B2 => n12029, C1 => n9178, C2 => 
                           n12025, A => n11026, ZN => n11023);
   U9454 : AOI222_X1 port map( A1 => n12021, A2 => n11616, B1 => n12018, B2 => 
                           n11680, C1 => n12014, C2 => n11744, ZN => n11026);
   U9455 : OAI221_X1 port map( B1 => n8921, B2 => n12029, C1 => n9177, C2 => 
                           n12025, A => n11009, ZN => n11006);
   U9456 : AOI222_X1 port map( A1 => n12021, A2 => n11617, B1 => n12018, B2 => 
                           n11681, C1 => n12014, C2 => n11745, ZN => n11009);
   U9457 : OAI221_X1 port map( B1 => n8920, B2 => n12029, C1 => n9176, C2 => 
                           n12025, A => n10992, ZN => n10989);
   U9458 : AOI222_X1 port map( A1 => n12021, A2 => n11618, B1 => n12018, B2 => 
                           n11682, C1 => n12014, C2 => n11746, ZN => n10992);
   U9459 : OAI221_X1 port map( B1 => n8919, B2 => n12029, C1 => n9175, C2 => 
                           n12025, A => n10975, ZN => n10972);
   U9460 : AOI222_X1 port map( A1 => n12021, A2 => n11619, B1 => n12018, B2 => 
                           n11683, C1 => n12014, C2 => n11747, ZN => n10975);
   U9461 : OAI221_X1 port map( B1 => n8918, B2 => n12029, C1 => n9174, C2 => 
                           n12025, A => n10958, ZN => n10955);
   U9462 : AOI222_X1 port map( A1 => n12021, A2 => n11620, B1 => n12018, B2 => 
                           n11684, C1 => n12014, C2 => n11748, ZN => n10958);
   U9463 : OAI221_X1 port map( B1 => n8917, B2 => n12029, C1 => n9173, C2 => 
                           n12025, A => n10941, ZN => n10938);
   U9464 : AOI222_X1 port map( A1 => n12021, A2 => n11621, B1 => n12017, B2 => 
                           n11685, C1 => n12013, C2 => n11749, ZN => n10941);
   U9465 : OAI221_X1 port map( B1 => n8916, B2 => n12029, C1 => n9172, C2 => 
                           n12025, A => n10924, ZN => n10921);
   U9466 : AOI222_X1 port map( A1 => n12021, A2 => n11622, B1 => n12017, B2 => 
                           n11686, C1 => n12013, C2 => n11750, ZN => n10924);
   U9467 : OAI221_X1 port map( B1 => n8915, B2 => n12029, C1 => n9171, C2 => 
                           n12025, A => n10907, ZN => n10904);
   U9468 : AOI222_X1 port map( A1 => n12021, A2 => n11623, B1 => n12017, B2 => 
                           n11687, C1 => n12013, C2 => n11751, ZN => n10907);
   U9469 : OAI221_X1 port map( B1 => n8914, B2 => n12029, C1 => n9170, C2 => 
                           n12025, A => n10890, ZN => n10887);
   U9470 : AOI222_X1 port map( A1 => n12021, A2 => n11624, B1 => n12017, B2 => 
                           n11688, C1 => n12013, C2 => n11752, ZN => n10890);
   U9471 : OAI221_X1 port map( B1 => n8913, B2 => n12030, C1 => n9169, C2 => 
                           n12026, A => n10873, ZN => n10870);
   U9472 : AOI222_X1 port map( A1 => n12022, A2 => n11625, B1 => n12017, B2 => 
                           n11689, C1 => n12013, C2 => n11753, ZN => n10873);
   U9473 : OAI221_X1 port map( B1 => n8912, B2 => n12030, C1 => n9168, C2 => 
                           n12026, A => n10856, ZN => n10853);
   U9474 : AOI222_X1 port map( A1 => n12022, A2 => n11626, B1 => n12017, B2 => 
                           n11690, C1 => n12013, C2 => n11754, ZN => n10856);
   U9475 : OAI221_X1 port map( B1 => n8911, B2 => n12030, C1 => n9167, C2 => 
                           n12026, A => n10839, ZN => n10836);
   U9476 : AOI222_X1 port map( A1 => n12022, A2 => n11627, B1 => n12017, B2 => 
                           n11691, C1 => n12013, C2 => n11755, ZN => n10839);
   U9477 : OAI221_X1 port map( B1 => n8910, B2 => n12030, C1 => n9166, C2 => 
                           n12026, A => n10822, ZN => n10819);
   U9478 : AOI222_X1 port map( A1 => n12022, A2 => n11628, B1 => n12017, B2 => 
                           n11692, C1 => n12013, C2 => n11756, ZN => n10822);
   U9479 : OAI221_X1 port map( B1 => n8909, B2 => n12030, C1 => n9165, C2 => 
                           n12026, A => n10805, ZN => n10802);
   U9480 : AOI222_X1 port map( A1 => n12022, A2 => n11629, B1 => n12017, B2 => 
                           n11693, C1 => n12013, C2 => n11757, ZN => n10805);
   U9481 : OAI221_X1 port map( B1 => n8908, B2 => n12030, C1 => n9164, C2 => 
                           n12026, A => n10788, ZN => n10785);
   U9482 : AOI222_X1 port map( A1 => n12022, A2 => n11630, B1 => n12017, B2 => 
                           n11694, C1 => n12013, C2 => n11758, ZN => n10788);
   U9483 : OAI221_X1 port map( B1 => n8907, B2 => n12030, C1 => n9163, C2 => 
                           n12026, A => n10771, ZN => n10768);
   U9484 : AOI222_X1 port map( A1 => n12022, A2 => n11631, B1 => n12017, B2 => 
                           n11695, C1 => n12013, C2 => n11759, ZN => n10771);
   U9485 : OAI221_X1 port map( B1 => n8906, B2 => n12030, C1 => n9162, C2 => 
                           n12026, A => n10754, ZN => n10751);
   U9486 : AOI222_X1 port map( A1 => n12022, A2 => n11632, B1 => n12017, B2 => 
                           n11696, C1 => n12013, C2 => n11760, ZN => n10754);
   U9487 : OAI221_X1 port map( B1 => n8905, B2 => n12030, C1 => n9161, C2 => 
                           n12026, A => n10737, ZN => n10734);
   U9488 : AOI222_X1 port map( A1 => n12022, A2 => n11633, B1 => n12016, B2 => 
                           n11697, C1 => n12012, C2 => n11761, ZN => n10737);
   U9489 : OAI221_X1 port map( B1 => n8904, B2 => n12030, C1 => n9160, C2 => 
                           n12026, A => n10720, ZN => n10717);
   U9490 : AOI222_X1 port map( A1 => n12022, A2 => n11634, B1 => n12016, B2 => 
                           n11698, C1 => n12012, C2 => n11762, ZN => n10720);
   U9491 : OAI221_X1 port map( B1 => n8903, B2 => n12030, C1 => n9159, C2 => 
                           n12026, A => n10703, ZN => n10700);
   U9492 : AOI222_X1 port map( A1 => n12022, A2 => n11635, B1 => n12016, B2 => 
                           n11699, C1 => n12012, C2 => n11763, ZN => n10703);
   U9493 : OAI221_X1 port map( B1 => n8902, B2 => n12030, C1 => n9158, C2 => 
                           n12026, A => n10686, ZN => n10683);
   U9494 : AOI222_X1 port map( A1 => n12022, A2 => n11636, B1 => n12016, B2 => 
                           n11700, C1 => n12012, C2 => n11764, ZN => n10686);
   U9495 : OAI221_X1 port map( B1 => n8901, B2 => n12031, C1 => n9157, C2 => 
                           n12027, A => n10669, ZN => n10666);
   U9496 : AOI222_X1 port map( A1 => n12023, A2 => n11637, B1 => n12016, B2 => 
                           n11701, C1 => n12012, C2 => n11765, ZN => n10669);
   U9497 : OAI221_X1 port map( B1 => n8900, B2 => n12031, C1 => n9156, C2 => 
                           n12027, A => n10652, ZN => n10649);
   U9498 : AOI222_X1 port map( A1 => n12023, A2 => n11638, B1 => n12016, B2 => 
                           n11702, C1 => n12012, C2 => n11766, ZN => n10652);
   U9499 : OAI221_X1 port map( B1 => n8899, B2 => n12031, C1 => n9155, C2 => 
                           n12027, A => n10635, ZN => n10632);
   U9500 : AOI222_X1 port map( A1 => n12023, A2 => n11639, B1 => n12016, B2 => 
                           n11703, C1 => n12012, C2 => n11767, ZN => n10635);
   U9501 : OAI221_X1 port map( B1 => n8898, B2 => n12031, C1 => n9154, C2 => 
                           n12027, A => n10618, ZN => n10615);
   U9502 : AOI222_X1 port map( A1 => n12023, A2 => n11640, B1 => n12016, B2 => 
                           n11704, C1 => n12012, C2 => n11768, ZN => n10618);
   U9503 : OAI221_X1 port map( B1 => n8897, B2 => n12031, C1 => n9153, C2 => 
                           n12027, A => n10601, ZN => n10598);
   U9504 : AOI222_X1 port map( A1 => n12023, A2 => n11641, B1 => n12016, B2 => 
                           n11705, C1 => n12012, C2 => n11769, ZN => n10601);
   U9505 : OAI221_X1 port map( B1 => n8896, B2 => n12031, C1 => n9152, C2 => 
                           n12027, A => n10584, ZN => n10581);
   U9506 : AOI222_X1 port map( A1 => n12023, A2 => n11642, B1 => n12016, B2 => 
                           n11706, C1 => n12012, C2 => n11770, ZN => n10584);
   U9507 : OAI221_X1 port map( B1 => n8895, B2 => n12031, C1 => n9151, C2 => 
                           n12027, A => n10567, ZN => n10564);
   U9508 : AOI222_X1 port map( A1 => n12023, A2 => n11643, B1 => n12016, B2 => 
                           n11707, C1 => n12012, C2 => n11771, ZN => n10567);
   U9509 : OAI221_X1 port map( B1 => n8894, B2 => n12031, C1 => n9150, C2 => 
                           n12027, A => n10537, ZN => n10528);
   U9510 : AOI222_X1 port map( A1 => n12023, A2 => n11644, B1 => n12016, B2 => 
                           n11708, C1 => n12012, C2 => n11772, ZN => n10537);
   U9511 : OAI221_X1 port map( B1 => n8925, B2 => n12173, C1 => n9181, C2 => 
                           n12169, A => n10496, ZN => n10491);
   U9512 : AOI222_X1 port map( A1 => n12165, A2 => n11613, B1 => n12162, B2 => 
                           n11677, C1 => n12158, C2 => n11741, ZN => n10496);
   U9513 : OAI221_X1 port map( B1 => n8924, B2 => n12173, C1 => n9180, C2 => 
                           n12169, A => n10460, ZN => n10457);
   U9514 : AOI222_X1 port map( A1 => n12165, A2 => n11614, B1 => n12162, B2 => 
                           n11678, C1 => n12158, C2 => n11742, ZN => n10460);
   U9515 : OAI221_X1 port map( B1 => n8923, B2 => n12173, C1 => n9179, C2 => 
                           n12169, A => n10443, ZN => n10440);
   U9516 : AOI222_X1 port map( A1 => n12165, A2 => n11615, B1 => n12162, B2 => 
                           n11679, C1 => n12158, C2 => n11743, ZN => n10443);
   U9517 : OAI221_X1 port map( B1 => n8922, B2 => n12173, C1 => n9178, C2 => 
                           n12169, A => n10426, ZN => n10423);
   U9518 : AOI222_X1 port map( A1 => n12165, A2 => n11616, B1 => n12162, B2 => 
                           n11680, C1 => n12158, C2 => n11744, ZN => n10426);
   U9519 : OAI221_X1 port map( B1 => n8921, B2 => n12173, C1 => n9177, C2 => 
                           n12169, A => n10409, ZN => n10406);
   U9520 : AOI222_X1 port map( A1 => n12165, A2 => n11617, B1 => n12162, B2 => 
                           n11681, C1 => n12158, C2 => n11745, ZN => n10409);
   U9521 : OAI221_X1 port map( B1 => n8920, B2 => n12173, C1 => n9176, C2 => 
                           n12169, A => n10392, ZN => n10389);
   U9522 : AOI222_X1 port map( A1 => n12165, A2 => n11618, B1 => n12162, B2 => 
                           n11682, C1 => n12158, C2 => n11746, ZN => n10392);
   U9523 : OAI221_X1 port map( B1 => n8919, B2 => n12173, C1 => n9175, C2 => 
                           n12169, A => n10375, ZN => n10372);
   U9524 : AOI222_X1 port map( A1 => n12165, A2 => n11619, B1 => n12162, B2 => 
                           n11683, C1 => n12158, C2 => n11747, ZN => n10375);
   U9525 : OAI221_X1 port map( B1 => n8918, B2 => n12173, C1 => n9174, C2 => 
                           n12169, A => n10358, ZN => n10355);
   U9526 : AOI222_X1 port map( A1 => n12165, A2 => n11620, B1 => n12162, B2 => 
                           n11684, C1 => n12158, C2 => n11748, ZN => n10358);
   U9527 : OAI221_X1 port map( B1 => n8917, B2 => n12173, C1 => n9173, C2 => 
                           n12169, A => n10341, ZN => n10338);
   U9528 : AOI222_X1 port map( A1 => n12165, A2 => n11621, B1 => n12161, B2 => 
                           n11685, C1 => n12157, C2 => n11749, ZN => n10341);
   U9529 : OAI221_X1 port map( B1 => n8916, B2 => n12173, C1 => n9172, C2 => 
                           n12169, A => n10324, ZN => n10321);
   U9530 : AOI222_X1 port map( A1 => n12165, A2 => n11622, B1 => n12161, B2 => 
                           n11686, C1 => n12157, C2 => n11750, ZN => n10324);
   U9531 : OAI221_X1 port map( B1 => n8915, B2 => n12173, C1 => n9171, C2 => 
                           n12169, A => n10307, ZN => n10304);
   U9532 : AOI222_X1 port map( A1 => n12165, A2 => n11623, B1 => n12161, B2 => 
                           n11687, C1 => n12157, C2 => n11751, ZN => n10307);
   U9533 : OAI221_X1 port map( B1 => n8914, B2 => n12173, C1 => n9170, C2 => 
                           n12169, A => n10290, ZN => n10287);
   U9534 : AOI222_X1 port map( A1 => n12165, A2 => n11624, B1 => n12161, B2 => 
                           n11688, C1 => n12157, C2 => n11752, ZN => n10290);
   U9535 : OAI221_X1 port map( B1 => n8913, B2 => n12174, C1 => n9169, C2 => 
                           n12170, A => n10273, ZN => n10270);
   U9536 : AOI222_X1 port map( A1 => n12166, A2 => n11625, B1 => n12161, B2 => 
                           n11689, C1 => n12157, C2 => n11753, ZN => n10273);
   U9537 : OAI221_X1 port map( B1 => n8912, B2 => n12174, C1 => n9168, C2 => 
                           n12170, A => n10256, ZN => n10253);
   U9538 : AOI222_X1 port map( A1 => n12166, A2 => n11626, B1 => n12161, B2 => 
                           n11690, C1 => n12157, C2 => n11754, ZN => n10256);
   U9539 : OAI221_X1 port map( B1 => n8911, B2 => n12174, C1 => n9167, C2 => 
                           n12170, A => n10239, ZN => n10236);
   U9540 : AOI222_X1 port map( A1 => n12166, A2 => n11627, B1 => n12161, B2 => 
                           n11691, C1 => n12157, C2 => n11755, ZN => n10239);
   U9541 : OAI221_X1 port map( B1 => n8910, B2 => n12174, C1 => n9166, C2 => 
                           n12170, A => n10222, ZN => n10219);
   U9542 : AOI222_X1 port map( A1 => n12166, A2 => n11628, B1 => n12161, B2 => 
                           n11692, C1 => n12157, C2 => n11756, ZN => n10222);
   U9543 : OAI221_X1 port map( B1 => n8909, B2 => n12174, C1 => n9165, C2 => 
                           n12170, A => n10205, ZN => n10202);
   U9544 : AOI222_X1 port map( A1 => n12166, A2 => n11629, B1 => n12161, B2 => 
                           n11693, C1 => n12157, C2 => n11757, ZN => n10205);
   U9545 : OAI221_X1 port map( B1 => n8908, B2 => n12174, C1 => n9164, C2 => 
                           n12170, A => n10188, ZN => n10185);
   U9546 : AOI222_X1 port map( A1 => n12166, A2 => n11630, B1 => n12161, B2 => 
                           n11694, C1 => n12157, C2 => n11758, ZN => n10188);
   U9547 : OAI221_X1 port map( B1 => n8907, B2 => n12174, C1 => n9163, C2 => 
                           n12170, A => n10171, ZN => n10168);
   U9548 : AOI222_X1 port map( A1 => n12166, A2 => n11631, B1 => n12161, B2 => 
                           n11695, C1 => n12157, C2 => n11759, ZN => n10171);
   U9549 : OAI221_X1 port map( B1 => n8906, B2 => n12174, C1 => n9162, C2 => 
                           n12170, A => n10154, ZN => n10151);
   U9550 : AOI222_X1 port map( A1 => n12166, A2 => n11632, B1 => n12161, B2 => 
                           n11696, C1 => n12157, C2 => n11760, ZN => n10154);
   U9551 : OAI221_X1 port map( B1 => n8905, B2 => n12174, C1 => n9161, C2 => 
                           n12170, A => n10137, ZN => n10134);
   U9552 : AOI222_X1 port map( A1 => n12166, A2 => n11633, B1 => n12160, B2 => 
                           n11697, C1 => n12156, C2 => n11761, ZN => n10137);
   U9553 : OAI221_X1 port map( B1 => n8904, B2 => n12174, C1 => n9160, C2 => 
                           n12170, A => n10120, ZN => n10117);
   U9554 : AOI222_X1 port map( A1 => n12166, A2 => n11634, B1 => n12160, B2 => 
                           n11698, C1 => n12156, C2 => n11762, ZN => n10120);
   U9555 : OAI221_X1 port map( B1 => n8903, B2 => n12174, C1 => n9159, C2 => 
                           n12170, A => n10103, ZN => n10100);
   U9556 : AOI222_X1 port map( A1 => n12166, A2 => n11635, B1 => n12160, B2 => 
                           n11699, C1 => n12156, C2 => n11763, ZN => n10103);
   U9557 : OAI221_X1 port map( B1 => n8902, B2 => n12174, C1 => n9158, C2 => 
                           n12170, A => n10086, ZN => n10083);
   U9558 : AOI222_X1 port map( A1 => n12166, A2 => n11636, B1 => n12160, B2 => 
                           n11700, C1 => n12156, C2 => n11764, ZN => n10086);
   U9559 : OAI221_X1 port map( B1 => n8901, B2 => n12175, C1 => n9157, C2 => 
                           n12171, A => n10069, ZN => n10066);
   U9560 : AOI222_X1 port map( A1 => n12167, A2 => n11637, B1 => n12160, B2 => 
                           n11701, C1 => n12156, C2 => n11765, ZN => n10069);
   U9561 : OAI221_X1 port map( B1 => n8900, B2 => n12175, C1 => n9156, C2 => 
                           n12171, A => n10052, ZN => n10049);
   U9562 : AOI222_X1 port map( A1 => n12167, A2 => n11638, B1 => n12160, B2 => 
                           n11702, C1 => n12156, C2 => n11766, ZN => n10052);
   U9563 : OAI221_X1 port map( B1 => n8899, B2 => n12175, C1 => n9155, C2 => 
                           n12171, A => n10035, ZN => n10032);
   U9564 : AOI222_X1 port map( A1 => n12167, A2 => n11639, B1 => n12160, B2 => 
                           n11703, C1 => n12156, C2 => n11767, ZN => n10035);
   U9565 : OAI221_X1 port map( B1 => n8898, B2 => n12175, C1 => n9154, C2 => 
                           n12171, A => n10018, ZN => n10015);
   U9566 : AOI222_X1 port map( A1 => n12167, A2 => n11640, B1 => n12160, B2 => 
                           n11704, C1 => n12156, C2 => n11768, ZN => n10018);
   U9567 : OAI221_X1 port map( B1 => n8897, B2 => n12175, C1 => n9153, C2 => 
                           n12171, A => n10001, ZN => n9998);
   U9568 : AOI222_X1 port map( A1 => n12167, A2 => n11641, B1 => n12160, B2 => 
                           n11705, C1 => n12156, C2 => n11769, ZN => n10001);
   U9569 : OAI221_X1 port map( B1 => n8896, B2 => n12175, C1 => n9152, C2 => 
                           n12171, A => n9984, ZN => n9981);
   U9570 : AOI222_X1 port map( A1 => n12167, A2 => n11642, B1 => n12160, B2 => 
                           n11706, C1 => n12156, C2 => n11770, ZN => n9984);
   U9571 : OAI221_X1 port map( B1 => n8895, B2 => n12175, C1 => n9151, C2 => 
                           n12171, A => n9967, ZN => n9964);
   U9572 : AOI222_X1 port map( A1 => n12167, A2 => n11643, B1 => n12160, B2 => 
                           n11707, C1 => n12156, C2 => n11771, ZN => n9967);
   U9573 : OAI221_X1 port map( B1 => n8894, B2 => n12175, C1 => n9150, C2 => 
                           n12171, A => n9937, ZN => n9928);
   U9574 : AOI222_X1 port map( A1 => n12167, A2 => n11644, B1 => n12160, B2 => 
                           n11708, C1 => n12156, C2 => n11772, ZN => n9937);
   U9575 : AOI221_X1 port map( B1 => n12062, B2 => DATAIN(0), C1 => n11100, C2 
                           => n10521, A => n11080, ZN => n11063);
   U9576 : OAI22_X1 port map( A1 => n11081, A2 => n12052, B1 => n9725, B2 => 
                           n12048, ZN => n11080);
   U9577 : NOR4_X1 port map( A1 => n11089, A2 => n11090, A3 => n11091, A4 => 
                           n11092, ZN => n11081);
   U9578 : OAI221_X1 port map( B1 => n9085, B2 => n12009, C1 => n8893, C2 => 
                           n12005, A => n11097, ZN => n11090);
   U9579 : AOI221_X1 port map( B1 => n12062, B2 => DATAIN(1), C1 => n11101, C2 
                           => n10521, A => n11053, ZN => n11046);
   U9580 : OAI22_X1 port map( A1 => n11054, A2 => n12052, B1 => n9724, B2 => 
                           n12048, ZN => n11053);
   U9581 : NOR4_X1 port map( A1 => n11055, A2 => n11056, A3 => n11057, A4 => 
                           n11058, ZN => n11054);
   U9582 : OAI221_X1 port map( B1 => n9084, B2 => n12009, C1 => n8892, C2 => 
                           n12005, A => n11061, ZN => n11056);
   U9583 : AOI221_X1 port map( B1 => n12062, B2 => DATAIN(2), C1 => n11102, C2 
                           => n10521, A => n11036, ZN => n11029);
   U9584 : OAI22_X1 port map( A1 => n11037, A2 => n12052, B1 => n9723, B2 => 
                           n12048, ZN => n11036);
   U9585 : NOR4_X1 port map( A1 => n11038, A2 => n11039, A3 => n11040, A4 => 
                           n11041, ZN => n11037);
   U9586 : OAI221_X1 port map( B1 => n9083, B2 => n12009, C1 => n8891, C2 => 
                           n12005, A => n11044, ZN => n11039);
   U9587 : AOI221_X1 port map( B1 => n12062, B2 => DATAIN(3), C1 => n11103, C2 
                           => n10521, A => n11019, ZN => n11012);
   U9588 : OAI22_X1 port map( A1 => n11020, A2 => n12052, B1 => n9722, B2 => 
                           n12048, ZN => n11019);
   U9589 : NOR4_X1 port map( A1 => n11021, A2 => n11022, A3 => n11023, A4 => 
                           n11024, ZN => n11020);
   U9590 : OAI221_X1 port map( B1 => n9082, B2 => n12009, C1 => n8890, C2 => 
                           n12005, A => n11027, ZN => n11022);
   U9591 : AOI221_X1 port map( B1 => n12062, B2 => DATAIN(4), C1 => n11104, C2 
                           => n10521, A => n11002, ZN => n10995);
   U9592 : OAI22_X1 port map( A1 => n11003, A2 => n12052, B1 => n9721, B2 => 
                           n12048, ZN => n11002);
   U9593 : NOR4_X1 port map( A1 => n11004, A2 => n11005, A3 => n11006, A4 => 
                           n11007, ZN => n11003);
   U9594 : OAI221_X1 port map( B1 => n9081, B2 => n12009, C1 => n8889, C2 => 
                           n12005, A => n11010, ZN => n11005);
   U9595 : AOI221_X1 port map( B1 => n12062, B2 => DATAIN(5), C1 => n11105, C2 
                           => n10521, A => n10985, ZN => n10978);
   U9596 : OAI22_X1 port map( A1 => n10986, A2 => n12052, B1 => n9720, B2 => 
                           n12048, ZN => n10985);
   U9597 : NOR4_X1 port map( A1 => n10987, A2 => n10988, A3 => n10989, A4 => 
                           n10990, ZN => n10986);
   U9598 : OAI221_X1 port map( B1 => n9080, B2 => n12009, C1 => n8888, C2 => 
                           n12005, A => n10993, ZN => n10988);
   U9599 : AOI221_X1 port map( B1 => n12062, B2 => DATAIN(6), C1 => n11106, C2 
                           => n10521, A => n10968, ZN => n10961);
   U9600 : OAI22_X1 port map( A1 => n10969, A2 => n12052, B1 => n9719, B2 => 
                           n12048, ZN => n10968);
   U9601 : NOR4_X1 port map( A1 => n10970, A2 => n10971, A3 => n10972, A4 => 
                           n10973, ZN => n10969);
   U9602 : OAI221_X1 port map( B1 => n9079, B2 => n12009, C1 => n8887, C2 => 
                           n12005, A => n10976, ZN => n10971);
   U9603 : AOI221_X1 port map( B1 => n12062, B2 => DATAIN(7), C1 => n11107, C2 
                           => n10521, A => n10951, ZN => n10944);
   U9604 : OAI22_X1 port map( A1 => n10952, A2 => n12052, B1 => n9718, B2 => 
                           n12048, ZN => n10951);
   U9605 : NOR4_X1 port map( A1 => n10953, A2 => n10954, A3 => n10955, A4 => 
                           n10956, ZN => n10952);
   U9606 : OAI221_X1 port map( B1 => n9078, B2 => n12009, C1 => n8886, C2 => 
                           n12005, A => n10959, ZN => n10954);
   U9607 : AOI221_X1 port map( B1 => n12061, B2 => DATAIN(8), C1 => n11108, C2 
                           => n12056, A => n10934, ZN => n10927);
   U9608 : OAI22_X1 port map( A1 => n10935, A2 => n12052, B1 => n9717, B2 => 
                           n12048, ZN => n10934);
   U9609 : NOR4_X1 port map( A1 => n10936, A2 => n10937, A3 => n10938, A4 => 
                           n10939, ZN => n10935);
   U9610 : OAI221_X1 port map( B1 => n9077, B2 => n12009, C1 => n8885, C2 => 
                           n12005, A => n10942, ZN => n10937);
   U9611 : AOI221_X1 port map( B1 => n12061, B2 => DATAIN(9), C1 => n11109, C2 
                           => n12056, A => n10917, ZN => n10910);
   U9612 : OAI22_X1 port map( A1 => n10918, A2 => n12052, B1 => n9716, B2 => 
                           n12048, ZN => n10917);
   U9613 : NOR4_X1 port map( A1 => n10919, A2 => n10920, A3 => n10921, A4 => 
                           n10922, ZN => n10918);
   U9614 : OAI221_X1 port map( B1 => n9076, B2 => n12009, C1 => n8884, C2 => 
                           n12005, A => n10925, ZN => n10920);
   U9615 : AOI221_X1 port map( B1 => n12061, B2 => DATAIN(10), C1 => n11110, C2
                           => n12056, A => n10900, ZN => n10893);
   U9616 : OAI22_X1 port map( A1 => n10901, A2 => n12052, B1 => n9715, B2 => 
                           n12048, ZN => n10900);
   U9617 : NOR4_X1 port map( A1 => n10902, A2 => n10903, A3 => n10904, A4 => 
                           n10905, ZN => n10901);
   U9618 : OAI221_X1 port map( B1 => n9075, B2 => n12009, C1 => n8883, C2 => 
                           n12005, A => n10908, ZN => n10903);
   U9619 : AOI221_X1 port map( B1 => n12061, B2 => DATAIN(11), C1 => n11111, C2
                           => n12056, A => n10883, ZN => n10876);
   U9620 : OAI22_X1 port map( A1 => n10884, A2 => n12052, B1 => n9714, B2 => 
                           n12048, ZN => n10883);
   U9621 : NOR4_X1 port map( A1 => n10885, A2 => n10886, A3 => n10887, A4 => 
                           n10888, ZN => n10884);
   U9622 : OAI221_X1 port map( B1 => n9074, B2 => n12009, C1 => n8882, C2 => 
                           n12005, A => n10891, ZN => n10886);
   U9623 : AOI221_X1 port map( B1 => n12061, B2 => DATAIN(12), C1 => n11112, C2
                           => n12056, A => n10866, ZN => n10859);
   U9624 : OAI22_X1 port map( A1 => n10867, A2 => n12053, B1 => n9713, B2 => 
                           n12049, ZN => n10866);
   U9625 : NOR4_X1 port map( A1 => n10868, A2 => n10869, A3 => n10870, A4 => 
                           n10871, ZN => n10867);
   U9626 : OAI221_X1 port map( B1 => n9073, B2 => n12010, C1 => n8881, C2 => 
                           n12006, A => n10874, ZN => n10869);
   U9627 : AOI221_X1 port map( B1 => n12061, B2 => DATAIN(13), C1 => n11113, C2
                           => n12056, A => n10849, ZN => n10842);
   U9628 : OAI22_X1 port map( A1 => n10850, A2 => n12053, B1 => n9712, B2 => 
                           n12049, ZN => n10849);
   U9629 : NOR4_X1 port map( A1 => n10851, A2 => n10852, A3 => n10853, A4 => 
                           n10854, ZN => n10850);
   U9630 : OAI221_X1 port map( B1 => n9072, B2 => n12010, C1 => n8880, C2 => 
                           n12006, A => n10857, ZN => n10852);
   U9631 : AOI221_X1 port map( B1 => n12061, B2 => DATAIN(14), C1 => n11114, C2
                           => n12056, A => n10832, ZN => n10825);
   U9632 : OAI22_X1 port map( A1 => n10833, A2 => n12053, B1 => n9711, B2 => 
                           n12049, ZN => n10832);
   U9633 : NOR4_X1 port map( A1 => n10834, A2 => n10835, A3 => n10836, A4 => 
                           n10837, ZN => n10833);
   U9634 : OAI221_X1 port map( B1 => n9071, B2 => n12010, C1 => n8879, C2 => 
                           n12006, A => n10840, ZN => n10835);
   U9635 : AOI221_X1 port map( B1 => n12061, B2 => DATAIN(15), C1 => n11115, C2
                           => n12056, A => n10815, ZN => n10808);
   U9636 : OAI22_X1 port map( A1 => n10816, A2 => n12053, B1 => n9710, B2 => 
                           n12049, ZN => n10815);
   U9637 : NOR4_X1 port map( A1 => n10817, A2 => n10818, A3 => n10819, A4 => 
                           n10820, ZN => n10816);
   U9638 : OAI221_X1 port map( B1 => n9070, B2 => n12010, C1 => n8878, C2 => 
                           n12006, A => n10823, ZN => n10818);
   U9639 : AOI221_X1 port map( B1 => n12061, B2 => DATAIN(16), C1 => n11116, C2
                           => n12056, A => n10798, ZN => n10791);
   U9640 : OAI22_X1 port map( A1 => n10799, A2 => n12053, B1 => n9709, B2 => 
                           n12049, ZN => n10798);
   U9641 : NOR4_X1 port map( A1 => n10800, A2 => n10801, A3 => n10802, A4 => 
                           n10803, ZN => n10799);
   U9642 : OAI221_X1 port map( B1 => n9069, B2 => n12010, C1 => n8877, C2 => 
                           n12006, A => n10806, ZN => n10801);
   U9643 : AOI221_X1 port map( B1 => n12061, B2 => DATAIN(17), C1 => n11117, C2
                           => n12056, A => n10781, ZN => n10774);
   U9644 : OAI22_X1 port map( A1 => n10782, A2 => n12053, B1 => n9708, B2 => 
                           n12049, ZN => n10781);
   U9645 : NOR4_X1 port map( A1 => n10783, A2 => n10784, A3 => n10785, A4 => 
                           n10786, ZN => n10782);
   U9646 : OAI221_X1 port map( B1 => n9068, B2 => n12010, C1 => n8876, C2 => 
                           n12006, A => n10789, ZN => n10784);
   U9647 : AOI221_X1 port map( B1 => n12061, B2 => DATAIN(18), C1 => n11118, C2
                           => n12056, A => n10764, ZN => n10757);
   U9648 : OAI22_X1 port map( A1 => n10765, A2 => n12053, B1 => n9707, B2 => 
                           n12049, ZN => n10764);
   U9649 : NOR4_X1 port map( A1 => n10766, A2 => n10767, A3 => n10768, A4 => 
                           n10769, ZN => n10765);
   U9650 : OAI221_X1 port map( B1 => n9067, B2 => n12010, C1 => n8875, C2 => 
                           n12006, A => n10772, ZN => n10767);
   U9651 : AOI221_X1 port map( B1 => n12061, B2 => DATAIN(19), C1 => n11119, C2
                           => n12056, A => n10747, ZN => n10740);
   U9652 : OAI22_X1 port map( A1 => n10748, A2 => n12053, B1 => n9706, B2 => 
                           n12049, ZN => n10747);
   U9653 : NOR4_X1 port map( A1 => n10749, A2 => n10750, A3 => n10751, A4 => 
                           n10752, ZN => n10748);
   U9654 : OAI221_X1 port map( B1 => n9066, B2 => n12010, C1 => n8874, C2 => 
                           n12006, A => n10755, ZN => n10750);
   U9655 : AOI221_X1 port map( B1 => n12060, B2 => DATAIN(20), C1 => n11120, C2
                           => n10521, A => n10730, ZN => n10723);
   U9656 : OAI22_X1 port map( A1 => n10731, A2 => n12053, B1 => n9705, B2 => 
                           n12049, ZN => n10730);
   U9657 : NOR4_X1 port map( A1 => n10732, A2 => n10733, A3 => n10734, A4 => 
                           n10735, ZN => n10731);
   U9658 : OAI221_X1 port map( B1 => n9065, B2 => n12010, C1 => n8873, C2 => 
                           n12006, A => n10738, ZN => n10733);
   U9659 : AOI221_X1 port map( B1 => n12060, B2 => DATAIN(21), C1 => n11121, C2
                           => n10521, A => n10713, ZN => n10706);
   U9660 : OAI22_X1 port map( A1 => n10714, A2 => n12053, B1 => n9704, B2 => 
                           n12049, ZN => n10713);
   U9661 : NOR4_X1 port map( A1 => n10715, A2 => n10716, A3 => n10717, A4 => 
                           n10718, ZN => n10714);
   U9662 : OAI221_X1 port map( B1 => n9064, B2 => n12010, C1 => n8872, C2 => 
                           n12006, A => n10721, ZN => n10716);
   U9663 : AOI221_X1 port map( B1 => n12060, B2 => DATAIN(22), C1 => n11122, C2
                           => n12056, A => n10696, ZN => n10689);
   U9664 : OAI22_X1 port map( A1 => n10697, A2 => n12053, B1 => n9703, B2 => 
                           n12049, ZN => n10696);
   U9665 : NOR4_X1 port map( A1 => n10698, A2 => n10699, A3 => n10700, A4 => 
                           n10701, ZN => n10697);
   U9666 : OAI221_X1 port map( B1 => n9063, B2 => n12010, C1 => n8871, C2 => 
                           n12006, A => n10704, ZN => n10699);
   U9667 : AOI221_X1 port map( B1 => n12060, B2 => DATAIN(23), C1 => n11123, C2
                           => n12056, A => n10679, ZN => n10672);
   U9668 : OAI22_X1 port map( A1 => n10680, A2 => n12053, B1 => n9702, B2 => 
                           n12049, ZN => n10679);
   U9669 : NOR4_X1 port map( A1 => n10681, A2 => n10682, A3 => n10683, A4 => 
                           n10684, ZN => n10680);
   U9670 : OAI221_X1 port map( B1 => n9062, B2 => n12010, C1 => n8870, C2 => 
                           n12006, A => n10687, ZN => n10682);
   U9671 : AOI221_X1 port map( B1 => n12060, B2 => DATAIN(24), C1 => n11124, C2
                           => n12056, A => n10662, ZN => n10655);
   U9672 : OAI22_X1 port map( A1 => n10663, A2 => n12052, B1 => n9701, B2 => 
                           n12050, ZN => n10662);
   U9673 : NOR4_X1 port map( A1 => n10664, A2 => n10665, A3 => n10666, A4 => 
                           n10667, ZN => n10663);
   U9674 : OAI221_X1 port map( B1 => n9061, B2 => n12011, C1 => n8869, C2 => 
                           n12007, A => n10670, ZN => n10665);
   U9675 : AOI221_X1 port map( B1 => n12060, B2 => DATAIN(25), C1 => n11125, C2
                           => n12056, A => n10645, ZN => n10638);
   U9676 : OAI22_X1 port map( A1 => n10646, A2 => n12053, B1 => n9700, B2 => 
                           n12050, ZN => n10645);
   U9677 : NOR4_X1 port map( A1 => n10647, A2 => n10648, A3 => n10649, A4 => 
                           n10650, ZN => n10646);
   U9678 : OAI221_X1 port map( B1 => n9060, B2 => n12011, C1 => n8868, C2 => 
                           n12007, A => n10653, ZN => n10648);
   U9679 : AOI221_X1 port map( B1 => n12060, B2 => DATAIN(26), C1 => n11126, C2
                           => n12056, A => n10628, ZN => n10621);
   U9680 : OAI22_X1 port map( A1 => n10629, A2 => n12052, B1 => n9699, B2 => 
                           n12050, ZN => n10628);
   U9681 : NOR4_X1 port map( A1 => n10630, A2 => n10631, A3 => n10632, A4 => 
                           n10633, ZN => n10629);
   U9682 : OAI221_X1 port map( B1 => n9059, B2 => n12011, C1 => n8867, C2 => 
                           n12007, A => n10636, ZN => n10631);
   U9683 : AOI221_X1 port map( B1 => n12060, B2 => DATAIN(27), C1 => n11127, C2
                           => n12056, A => n10611, ZN => n10604);
   U9684 : OAI22_X1 port map( A1 => n10612, A2 => n12053, B1 => n9698, B2 => 
                           n12050, ZN => n10611);
   U9685 : NOR4_X1 port map( A1 => n10613, A2 => n10614, A3 => n10615, A4 => 
                           n10616, ZN => n10612);
   U9686 : OAI221_X1 port map( B1 => n9058, B2 => n12011, C1 => n8866, C2 => 
                           n12007, A => n10619, ZN => n10614);
   U9687 : AOI221_X1 port map( B1 => n12060, B2 => DATAIN(28), C1 => n11128, C2
                           => n12056, A => n10594, ZN => n10587);
   U9688 : OAI22_X1 port map( A1 => n10595, A2 => n12052, B1 => n9697, B2 => 
                           n12050, ZN => n10594);
   U9689 : NOR4_X1 port map( A1 => n10596, A2 => n10597, A3 => n10598, A4 => 
                           n10599, ZN => n10595);
   U9690 : OAI221_X1 port map( B1 => n9057, B2 => n12011, C1 => n8865, C2 => 
                           n12007, A => n10602, ZN => n10597);
   U9691 : AOI221_X1 port map( B1 => n12060, B2 => DATAIN(29), C1 => n11129, C2
                           => n12056, A => n10577, ZN => n10570);
   U9692 : OAI22_X1 port map( A1 => n10578, A2 => n12053, B1 => n9696, B2 => 
                           n12050, ZN => n10577);
   U9693 : NOR4_X1 port map( A1 => n10579, A2 => n10580, A3 => n10581, A4 => 
                           n10582, ZN => n10578);
   U9694 : OAI221_X1 port map( B1 => n9056, B2 => n12011, C1 => n8864, C2 => 
                           n12007, A => n10585, ZN => n10580);
   U9695 : AOI221_X1 port map( B1 => n12060, B2 => DATAIN(30), C1 => n11130, C2
                           => n12056, A => n10560, ZN => n10553);
   U9696 : OAI22_X1 port map( A1 => n10561, A2 => n12052, B1 => n9695, B2 => 
                           n12050, ZN => n10560);
   U9697 : NOR4_X1 port map( A1 => n10562, A2 => n10563, A3 => n10564, A4 => 
                           n10565, ZN => n10561);
   U9698 : OAI221_X1 port map( B1 => n9055, B2 => n12011, C1 => n8863, C2 => 
                           n12007, A => n10568, ZN => n10563);
   U9699 : AOI221_X1 port map( B1 => n12060, B2 => DATAIN(31), C1 => n11131, C2
                           => n12056, A => n10522, ZN => n10500);
   U9700 : OAI22_X1 port map( A1 => n10523, A2 => n12053, B1 => n9694, B2 => 
                           n12050, ZN => n10522);
   U9701 : NOR4_X1 port map( A1 => n10526, A2 => n10527, A3 => n10528, A4 => 
                           n10529, ZN => n10523);
   U9702 : OAI221_X1 port map( B1 => n9054, B2 => n12011, C1 => n8862, C2 => 
                           n12007, A => n10543, ZN => n10527);
   U9703 : AOI221_X1 port map( B1 => n12206, B2 => DATAIN(0), C1 => n11132, C2 
                           => n9921, A => n10480, ZN => n10463);
   U9704 : OAI22_X1 port map( A1 => n10481, A2 => n12196, B1 => n9725, B2 => 
                           n12192, ZN => n10480);
   U9705 : NOR4_X1 port map( A1 => n10489, A2 => n10490, A3 => n10491, A4 => 
                           n10492, ZN => n10481);
   U9706 : OAI221_X1 port map( B1 => n9085, B2 => n12153, C1 => n8893, C2 => 
                           n12149, A => n10497, ZN => n10490);
   U9707 : AOI221_X1 port map( B1 => n12206, B2 => DATAIN(1), C1 => n11133, C2 
                           => n9921, A => n10453, ZN => n10446);
   U9708 : OAI22_X1 port map( A1 => n10454, A2 => n12196, B1 => n9724, B2 => 
                           n12192, ZN => n10453);
   U9709 : NOR4_X1 port map( A1 => n10455, A2 => n10456, A3 => n10457, A4 => 
                           n10458, ZN => n10454);
   U9710 : OAI221_X1 port map( B1 => n9084, B2 => n12153, C1 => n8892, C2 => 
                           n12149, A => n10461, ZN => n10456);
   U9711 : AOI221_X1 port map( B1 => n12206, B2 => DATAIN(2), C1 => n11134, C2 
                           => n9921, A => n10436, ZN => n10429);
   U9712 : OAI22_X1 port map( A1 => n10437, A2 => n12196, B1 => n9723, B2 => 
                           n12192, ZN => n10436);
   U9713 : NOR4_X1 port map( A1 => n10438, A2 => n10439, A3 => n10440, A4 => 
                           n10441, ZN => n10437);
   U9714 : OAI221_X1 port map( B1 => n9083, B2 => n12153, C1 => n8891, C2 => 
                           n12149, A => n10444, ZN => n10439);
   U9715 : AOI221_X1 port map( B1 => n12206, B2 => DATAIN(3), C1 => n11135, C2 
                           => n9921, A => n10419, ZN => n10412);
   U9716 : OAI22_X1 port map( A1 => n10420, A2 => n12196, B1 => n9722, B2 => 
                           n12192, ZN => n10419);
   U9717 : NOR4_X1 port map( A1 => n10421, A2 => n10422, A3 => n10423, A4 => 
                           n10424, ZN => n10420);
   U9718 : OAI221_X1 port map( B1 => n9082, B2 => n12153, C1 => n8890, C2 => 
                           n12149, A => n10427, ZN => n10422);
   U9719 : AOI221_X1 port map( B1 => n12206, B2 => DATAIN(4), C1 => n11136, C2 
                           => n9921, A => n10402, ZN => n10395);
   U9720 : OAI22_X1 port map( A1 => n10403, A2 => n12196, B1 => n9721, B2 => 
                           n12192, ZN => n10402);
   U9721 : NOR4_X1 port map( A1 => n10404, A2 => n10405, A3 => n10406, A4 => 
                           n10407, ZN => n10403);
   U9722 : OAI221_X1 port map( B1 => n9081, B2 => n12153, C1 => n8889, C2 => 
                           n12149, A => n10410, ZN => n10405);
   U9723 : AOI221_X1 port map( B1 => n12206, B2 => DATAIN(5), C1 => n11137, C2 
                           => n9921, A => n10385, ZN => n10378);
   U9724 : OAI22_X1 port map( A1 => n10386, A2 => n12196, B1 => n9720, B2 => 
                           n12192, ZN => n10385);
   U9725 : NOR4_X1 port map( A1 => n10387, A2 => n10388, A3 => n10389, A4 => 
                           n10390, ZN => n10386);
   U9726 : OAI221_X1 port map( B1 => n9080, B2 => n12153, C1 => n8888, C2 => 
                           n12149, A => n10393, ZN => n10388);
   U9727 : AOI221_X1 port map( B1 => n12206, B2 => DATAIN(6), C1 => n11138, C2 
                           => n9921, A => n10368, ZN => n10361);
   U9728 : OAI22_X1 port map( A1 => n10369, A2 => n12196, B1 => n9719, B2 => 
                           n12192, ZN => n10368);
   U9729 : NOR4_X1 port map( A1 => n10370, A2 => n10371, A3 => n10372, A4 => 
                           n10373, ZN => n10369);
   U9730 : OAI221_X1 port map( B1 => n9079, B2 => n12153, C1 => n8887, C2 => 
                           n12149, A => n10376, ZN => n10371);
   U9731 : AOI221_X1 port map( B1 => n12206, B2 => DATAIN(7), C1 => n11139, C2 
                           => n9921, A => n10351, ZN => n10344);
   U9732 : OAI22_X1 port map( A1 => n10352, A2 => n12196, B1 => n9718, B2 => 
                           n12192, ZN => n10351);
   U9733 : NOR4_X1 port map( A1 => n10353, A2 => n10354, A3 => n10355, A4 => 
                           n10356, ZN => n10352);
   U9734 : OAI221_X1 port map( B1 => n9078, B2 => n12153, C1 => n8886, C2 => 
                           n12149, A => n10359, ZN => n10354);
   U9735 : AOI221_X1 port map( B1 => n12205, B2 => DATAIN(8), C1 => n11140, C2 
                           => n12200, A => n10334, ZN => n10327);
   U9736 : OAI22_X1 port map( A1 => n10335, A2 => n12196, B1 => n9717, B2 => 
                           n12192, ZN => n10334);
   U9737 : NOR4_X1 port map( A1 => n10336, A2 => n10337, A3 => n10338, A4 => 
                           n10339, ZN => n10335);
   U9738 : OAI221_X1 port map( B1 => n9077, B2 => n12153, C1 => n8885, C2 => 
                           n12149, A => n10342, ZN => n10337);
   U9739 : AOI221_X1 port map( B1 => n12205, B2 => DATAIN(9), C1 => n11141, C2 
                           => n12200, A => n10317, ZN => n10310);
   U9740 : OAI22_X1 port map( A1 => n10318, A2 => n12196, B1 => n9716, B2 => 
                           n12192, ZN => n10317);
   U9741 : NOR4_X1 port map( A1 => n10319, A2 => n10320, A3 => n10321, A4 => 
                           n10322, ZN => n10318);
   U9742 : OAI221_X1 port map( B1 => n9076, B2 => n12153, C1 => n8884, C2 => 
                           n12149, A => n10325, ZN => n10320);
   U9743 : AOI221_X1 port map( B1 => n12205, B2 => DATAIN(10), C1 => n11142, C2
                           => n12200, A => n10300, ZN => n10293);
   U9744 : OAI22_X1 port map( A1 => n10301, A2 => n12196, B1 => n9715, B2 => 
                           n12192, ZN => n10300);
   U9745 : NOR4_X1 port map( A1 => n10302, A2 => n10303, A3 => n10304, A4 => 
                           n10305, ZN => n10301);
   U9746 : OAI221_X1 port map( B1 => n9075, B2 => n12153, C1 => n8883, C2 => 
                           n12149, A => n10308, ZN => n10303);
   U9747 : AOI221_X1 port map( B1 => n12205, B2 => DATAIN(11), C1 => n11143, C2
                           => n12200, A => n10283, ZN => n10276);
   U9748 : OAI22_X1 port map( A1 => n10284, A2 => n12196, B1 => n9714, B2 => 
                           n12192, ZN => n10283);
   U9749 : NOR4_X1 port map( A1 => n10285, A2 => n10286, A3 => n10287, A4 => 
                           n10288, ZN => n10284);
   U9750 : OAI221_X1 port map( B1 => n9074, B2 => n12153, C1 => n8882, C2 => 
                           n12149, A => n10291, ZN => n10286);
   U9751 : AOI221_X1 port map( B1 => n12205, B2 => DATAIN(12), C1 => n11144, C2
                           => n12200, A => n10266, ZN => n10259);
   U9752 : OAI22_X1 port map( A1 => n10267, A2 => n12197, B1 => n9713, B2 => 
                           n12193, ZN => n10266);
   U9753 : NOR4_X1 port map( A1 => n10268, A2 => n10269, A3 => n10270, A4 => 
                           n10271, ZN => n10267);
   U9754 : OAI221_X1 port map( B1 => n9073, B2 => n12154, C1 => n8881, C2 => 
                           n12150, A => n10274, ZN => n10269);
   U9755 : AOI221_X1 port map( B1 => n12205, B2 => DATAIN(13), C1 => n11145, C2
                           => n12200, A => n10249, ZN => n10242);
   U9756 : OAI22_X1 port map( A1 => n10250, A2 => n12197, B1 => n9712, B2 => 
                           n12193, ZN => n10249);
   U9757 : NOR4_X1 port map( A1 => n10251, A2 => n10252, A3 => n10253, A4 => 
                           n10254, ZN => n10250);
   U9758 : OAI221_X1 port map( B1 => n9072, B2 => n12154, C1 => n8880, C2 => 
                           n12150, A => n10257, ZN => n10252);
   U9759 : AOI221_X1 port map( B1 => n12205, B2 => DATAIN(14), C1 => n11146, C2
                           => n12200, A => n10232, ZN => n10225);
   U9760 : OAI22_X1 port map( A1 => n10233, A2 => n12197, B1 => n9711, B2 => 
                           n12193, ZN => n10232);
   U9761 : NOR4_X1 port map( A1 => n10234, A2 => n10235, A3 => n10236, A4 => 
                           n10237, ZN => n10233);
   U9762 : OAI221_X1 port map( B1 => n9071, B2 => n12154, C1 => n8879, C2 => 
                           n12150, A => n10240, ZN => n10235);
   U9763 : AOI221_X1 port map( B1 => n12205, B2 => DATAIN(15), C1 => n11147, C2
                           => n12200, A => n10215, ZN => n10208);
   U9764 : OAI22_X1 port map( A1 => n10216, A2 => n12197, B1 => n9710, B2 => 
                           n12193, ZN => n10215);
   U9765 : NOR4_X1 port map( A1 => n10217, A2 => n10218, A3 => n10219, A4 => 
                           n10220, ZN => n10216);
   U9766 : OAI221_X1 port map( B1 => n9070, B2 => n12154, C1 => n8878, C2 => 
                           n12150, A => n10223, ZN => n10218);
   U9767 : AOI221_X1 port map( B1 => n12205, B2 => DATAIN(16), C1 => n11148, C2
                           => n12200, A => n10198, ZN => n10191);
   U9768 : OAI22_X1 port map( A1 => n10199, A2 => n12197, B1 => n9709, B2 => 
                           n12193, ZN => n10198);
   U9769 : NOR4_X1 port map( A1 => n10200, A2 => n10201, A3 => n10202, A4 => 
                           n10203, ZN => n10199);
   U9770 : OAI221_X1 port map( B1 => n9069, B2 => n12154, C1 => n8877, C2 => 
                           n12150, A => n10206, ZN => n10201);
   U9771 : AOI221_X1 port map( B1 => n12205, B2 => DATAIN(17), C1 => n11149, C2
                           => n12200, A => n10181, ZN => n10174);
   U9772 : OAI22_X1 port map( A1 => n10182, A2 => n12197, B1 => n9708, B2 => 
                           n12193, ZN => n10181);
   U9773 : NOR4_X1 port map( A1 => n10183, A2 => n10184, A3 => n10185, A4 => 
                           n10186, ZN => n10182);
   U9774 : OAI221_X1 port map( B1 => n9068, B2 => n12154, C1 => n8876, C2 => 
                           n12150, A => n10189, ZN => n10184);
   U9775 : AOI221_X1 port map( B1 => n12205, B2 => DATAIN(18), C1 => n11150, C2
                           => n12200, A => n10164, ZN => n10157);
   U9776 : OAI22_X1 port map( A1 => n10165, A2 => n12197, B1 => n9707, B2 => 
                           n12193, ZN => n10164);
   U9777 : NOR4_X1 port map( A1 => n10166, A2 => n10167, A3 => n10168, A4 => 
                           n10169, ZN => n10165);
   U9778 : OAI221_X1 port map( B1 => n9067, B2 => n12154, C1 => n8875, C2 => 
                           n12150, A => n10172, ZN => n10167);
   U9779 : AOI221_X1 port map( B1 => n12205, B2 => DATAIN(19), C1 => n11151, C2
                           => n12200, A => n10147, ZN => n10140);
   U9780 : OAI22_X1 port map( A1 => n10148, A2 => n12197, B1 => n9706, B2 => 
                           n12193, ZN => n10147);
   U9781 : NOR4_X1 port map( A1 => n10149, A2 => n10150, A3 => n10151, A4 => 
                           n10152, ZN => n10148);
   U9782 : OAI221_X1 port map( B1 => n9066, B2 => n12154, C1 => n8874, C2 => 
                           n12150, A => n10155, ZN => n10150);
   U9783 : AOI221_X1 port map( B1 => n12204, B2 => DATAIN(20), C1 => n11152, C2
                           => n9921, A => n10130, ZN => n10123);
   U9784 : OAI22_X1 port map( A1 => n10131, A2 => n12197, B1 => n9705, B2 => 
                           n12193, ZN => n10130);
   U9785 : NOR4_X1 port map( A1 => n10132, A2 => n10133, A3 => n10134, A4 => 
                           n10135, ZN => n10131);
   U9786 : OAI221_X1 port map( B1 => n9065, B2 => n12154, C1 => n8873, C2 => 
                           n12150, A => n10138, ZN => n10133);
   U9787 : AOI221_X1 port map( B1 => n12204, B2 => DATAIN(21), C1 => n11153, C2
                           => n9921, A => n10113, ZN => n10106);
   U9788 : OAI22_X1 port map( A1 => n10114, A2 => n12197, B1 => n9704, B2 => 
                           n12193, ZN => n10113);
   U9789 : NOR4_X1 port map( A1 => n10115, A2 => n10116, A3 => n10117, A4 => 
                           n10118, ZN => n10114);
   U9790 : OAI221_X1 port map( B1 => n9064, B2 => n12154, C1 => n8872, C2 => 
                           n12150, A => n10121, ZN => n10116);
   U9791 : AOI221_X1 port map( B1 => n12204, B2 => DATAIN(22), C1 => n11154, C2
                           => n12200, A => n10096, ZN => n10089);
   U9792 : OAI22_X1 port map( A1 => n10097, A2 => n12197, B1 => n9703, B2 => 
                           n12193, ZN => n10096);
   U9793 : NOR4_X1 port map( A1 => n10098, A2 => n10099, A3 => n10100, A4 => 
                           n10101, ZN => n10097);
   U9794 : OAI221_X1 port map( B1 => n9063, B2 => n12154, C1 => n8871, C2 => 
                           n12150, A => n10104, ZN => n10099);
   U9795 : AOI221_X1 port map( B1 => n12204, B2 => DATAIN(23), C1 => n11155, C2
                           => n12200, A => n10079, ZN => n10072);
   U9796 : OAI22_X1 port map( A1 => n10080, A2 => n12197, B1 => n9702, B2 => 
                           n12193, ZN => n10079);
   U9797 : NOR4_X1 port map( A1 => n10081, A2 => n10082, A3 => n10083, A4 => 
                           n10084, ZN => n10080);
   U9798 : OAI221_X1 port map( B1 => n9062, B2 => n12154, C1 => n8870, C2 => 
                           n12150, A => n10087, ZN => n10082);
   U9799 : AOI221_X1 port map( B1 => n12204, B2 => DATAIN(24), C1 => n11156, C2
                           => n12200, A => n10062, ZN => n10055);
   U9800 : OAI22_X1 port map( A1 => n10063, A2 => n12196, B1 => n9701, B2 => 
                           n12194, ZN => n10062);
   U9801 : NOR4_X1 port map( A1 => n10064, A2 => n10065, A3 => n10066, A4 => 
                           n10067, ZN => n10063);
   U9802 : OAI221_X1 port map( B1 => n9061, B2 => n12155, C1 => n8869, C2 => 
                           n12151, A => n10070, ZN => n10065);
   U9803 : AOI221_X1 port map( B1 => n12204, B2 => DATAIN(25), C1 => n11157, C2
                           => n12200, A => n10045, ZN => n10038);
   U9804 : OAI22_X1 port map( A1 => n10046, A2 => n12197, B1 => n9700, B2 => 
                           n12194, ZN => n10045);
   U9805 : NOR4_X1 port map( A1 => n10047, A2 => n10048, A3 => n10049, A4 => 
                           n10050, ZN => n10046);
   U9806 : OAI221_X1 port map( B1 => n9060, B2 => n12155, C1 => n8868, C2 => 
                           n12151, A => n10053, ZN => n10048);
   U9807 : AOI221_X1 port map( B1 => n12204, B2 => DATAIN(26), C1 => n11158, C2
                           => n12200, A => n10028, ZN => n10021);
   U9808 : OAI22_X1 port map( A1 => n10029, A2 => n12196, B1 => n9699, B2 => 
                           n12194, ZN => n10028);
   U9809 : NOR4_X1 port map( A1 => n10030, A2 => n10031, A3 => n10032, A4 => 
                           n10033, ZN => n10029);
   U9810 : OAI221_X1 port map( B1 => n9059, B2 => n12155, C1 => n8867, C2 => 
                           n12151, A => n10036, ZN => n10031);
   U9811 : AOI221_X1 port map( B1 => n12204, B2 => DATAIN(27), C1 => n11159, C2
                           => n12200, A => n10011, ZN => n10004);
   U9812 : OAI22_X1 port map( A1 => n10012, A2 => n12197, B1 => n9698, B2 => 
                           n12194, ZN => n10011);
   U9813 : NOR4_X1 port map( A1 => n10013, A2 => n10014, A3 => n10015, A4 => 
                           n10016, ZN => n10012);
   U9814 : OAI221_X1 port map( B1 => n9058, B2 => n12155, C1 => n8866, C2 => 
                           n12151, A => n10019, ZN => n10014);
   U9815 : AOI221_X1 port map( B1 => n12204, B2 => DATAIN(28), C1 => n11160, C2
                           => n12200, A => n9994, ZN => n9987);
   U9816 : OAI22_X1 port map( A1 => n9995, A2 => n12196, B1 => n9697, B2 => 
                           n12194, ZN => n9994);
   U9817 : NOR4_X1 port map( A1 => n9996, A2 => n9997, A3 => n9998, A4 => n9999
                           , ZN => n9995);
   U9818 : OAI221_X1 port map( B1 => n9057, B2 => n12155, C1 => n8865, C2 => 
                           n12151, A => n10002, ZN => n9997);
   U9819 : AOI221_X1 port map( B1 => n12204, B2 => DATAIN(29), C1 => n11161, C2
                           => n12200, A => n9977, ZN => n9970);
   U9820 : OAI22_X1 port map( A1 => n9978, A2 => n12197, B1 => n9696, B2 => 
                           n12194, ZN => n9977);
   U9821 : NOR4_X1 port map( A1 => n9979, A2 => n9980, A3 => n9981, A4 => n9982
                           , ZN => n9978);
   U9822 : OAI221_X1 port map( B1 => n9056, B2 => n12155, C1 => n8864, C2 => 
                           n12151, A => n9985, ZN => n9980);
   U9823 : AOI221_X1 port map( B1 => n12204, B2 => DATAIN(30), C1 => n11162, C2
                           => n12200, A => n9960, ZN => n9953);
   U9824 : OAI22_X1 port map( A1 => n9961, A2 => n12196, B1 => n9695, B2 => 
                           n12194, ZN => n9960);
   U9825 : NOR4_X1 port map( A1 => n9962, A2 => n9963, A3 => n9964, A4 => n9965
                           , ZN => n9961);
   U9826 : OAI221_X1 port map( B1 => n9055, B2 => n12155, C1 => n8863, C2 => 
                           n12151, A => n9968, ZN => n9963);
   U9827 : AOI221_X1 port map( B1 => n12204, B2 => DATAIN(31), C1 => n11163, C2
                           => n12200, A => n9922, ZN => n9900);
   U9828 : OAI22_X1 port map( A1 => n9923, A2 => n12197, B1 => n9694, B2 => 
                           n12194, ZN => n9922);
   U9829 : NOR4_X1 port map( A1 => n9926, A2 => n9927, A3 => n9928, A4 => n9929
                           , ZN => n9923);
   U9830 : OAI221_X1 port map( B1 => n9054, B2 => n12155, C1 => n8862, C2 => 
                           n12151, A => n9943, ZN => n9927);
   U9831 : NAND4_X1 port map( A1 => n11063, A2 => n11064, A3 => n11065, A4 => 
                           n11066, ZN => n1484);
   U9832 : AOI221_X1 port map( B1 => n12077, B2 => n8007, C1 => n12073, C2 => 
                           n11517, A => n11079, ZN => n11064);
   U9833 : AOI221_X1 port map( B1 => n12093, B2 => n11516, C1 => n12089, C2 => 
                           n11196, A => n11074, ZN => n11065);
   U9834 : AOI221_X1 port map( B1 => n12113, B2 => n11549, C1 => n12109, C2 => 
                           n11228, A => n11067, ZN => n11066);
   U9835 : NAND4_X1 port map( A1 => n11046, A2 => n11047, A3 => n11048, A4 => 
                           n11049, ZN => n1486);
   U9836 : AOI221_X1 port map( B1 => n12077, B2 => n8008, C1 => n12073, C2 => 
                           n11518, A => n11052, ZN => n11047);
   U9837 : AOI221_X1 port map( B1 => n12093, B2 => n11837, C1 => n12089, C2 => 
                           n11197, A => n11051, ZN => n11048);
   U9838 : AOI221_X1 port map( B1 => n12113, B2 => n11550, C1 => n12109, C2 => 
                           n11229, A => n11050, ZN => n11049);
   U9839 : NAND4_X1 port map( A1 => n11029, A2 => n11030, A3 => n11031, A4 => 
                           n11032, ZN => n1488);
   U9840 : AOI221_X1 port map( B1 => n12077, B2 => n8009, C1 => n12073, C2 => 
                           n11519, A => n11035, ZN => n11030);
   U9841 : AOI221_X1 port map( B1 => n12093, B2 => n11838, C1 => n12089, C2 => 
                           n11198, A => n11034, ZN => n11031);
   U9842 : AOI221_X1 port map( B1 => n12113, B2 => n11551, C1 => n12109, C2 => 
                           n11230, A => n11033, ZN => n11032);
   U9843 : NAND4_X1 port map( A1 => n11012, A2 => n11013, A3 => n11014, A4 => 
                           n11015, ZN => n1490);
   U9844 : AOI221_X1 port map( B1 => n12077, B2 => n8010, C1 => n12073, C2 => 
                           n11520, A => n11018, ZN => n11013);
   U9845 : AOI221_X1 port map( B1 => n12093, B2 => n11839, C1 => n12089, C2 => 
                           n11199, A => n11017, ZN => n11014);
   U9846 : AOI221_X1 port map( B1 => n12113, B2 => n11552, C1 => n12109, C2 => 
                           n11231, A => n11016, ZN => n11015);
   U9847 : NAND4_X1 port map( A1 => n10995, A2 => n10996, A3 => n10997, A4 => 
                           n10998, ZN => n1492);
   U9848 : AOI221_X1 port map( B1 => n12077, B2 => n8011, C1 => n12073, C2 => 
                           n11521, A => n11001, ZN => n10996);
   U9849 : AOI221_X1 port map( B1 => n12093, B2 => n11840, C1 => n12089, C2 => 
                           n11200, A => n11000, ZN => n10997);
   U9850 : AOI221_X1 port map( B1 => n12113, B2 => n11553, C1 => n12109, C2 => 
                           n11232, A => n10999, ZN => n10998);
   U9851 : NAND4_X1 port map( A1 => n10978, A2 => n10979, A3 => n10980, A4 => 
                           n10981, ZN => n1494);
   U9852 : AOI221_X1 port map( B1 => n12077, B2 => n8012, C1 => n12073, C2 => 
                           n11522, A => n10984, ZN => n10979);
   U9853 : AOI221_X1 port map( B1 => n12093, B2 => n11841, C1 => n12089, C2 => 
                           n11201, A => n10983, ZN => n10980);
   U9854 : AOI221_X1 port map( B1 => n12113, B2 => n11554, C1 => n12109, C2 => 
                           n11233, A => n10982, ZN => n10981);
   U9855 : NAND4_X1 port map( A1 => n10961, A2 => n10962, A3 => n10963, A4 => 
                           n10964, ZN => n1496);
   U9856 : AOI221_X1 port map( B1 => n12077, B2 => n8013, C1 => n12073, C2 => 
                           n11523, A => n10967, ZN => n10962);
   U9857 : AOI221_X1 port map( B1 => n12093, B2 => n11842, C1 => n12089, C2 => 
                           n11202, A => n10966, ZN => n10963);
   U9858 : AOI221_X1 port map( B1 => n12113, B2 => n11555, C1 => n12109, C2 => 
                           n11234, A => n10965, ZN => n10964);
   U9859 : NAND4_X1 port map( A1 => n10944, A2 => n10945, A3 => n10946, A4 => 
                           n10947, ZN => n1498);
   U9860 : AOI221_X1 port map( B1 => n12077, B2 => n8014, C1 => n12073, C2 => 
                           n11524, A => n10950, ZN => n10945);
   U9861 : AOI221_X1 port map( B1 => n12093, B2 => n11843, C1 => n12089, C2 => 
                           n11203, A => n10949, ZN => n10946);
   U9862 : AOI221_X1 port map( B1 => n12113, B2 => n11556, C1 => n12109, C2 => 
                           n11235, A => n10948, ZN => n10947);
   U9863 : NAND4_X1 port map( A1 => n10927, A2 => n10928, A3 => n10929, A4 => 
                           n10930, ZN => n1500);
   U9864 : AOI221_X1 port map( B1 => n12077, B2 => n8015, C1 => n12073, C2 => 
                           n11525, A => n10933, ZN => n10928);
   U9865 : AOI221_X1 port map( B1 => n12093, B2 => n11844, C1 => n12089, C2 => 
                           n11204, A => n10932, ZN => n10929);
   U9866 : AOI221_X1 port map( B1 => n12113, B2 => n11557, C1 => n12109, C2 => 
                           n11236, A => n10931, ZN => n10930);
   U9867 : NAND4_X1 port map( A1 => n10910, A2 => n10911, A3 => n10912, A4 => 
                           n10913, ZN => n1502);
   U9868 : AOI221_X1 port map( B1 => n12077, B2 => n8016, C1 => n12073, C2 => 
                           n11526, A => n10916, ZN => n10911);
   U9869 : AOI221_X1 port map( B1 => n12093, B2 => n11845, C1 => n12089, C2 => 
                           n11205, A => n10915, ZN => n10912);
   U9870 : AOI221_X1 port map( B1 => n12113, B2 => n11558, C1 => n12109, C2 => 
                           n11237, A => n10914, ZN => n10913);
   U9871 : NAND4_X1 port map( A1 => n10893, A2 => n10894, A3 => n10895, A4 => 
                           n10896, ZN => n1504);
   U9872 : AOI221_X1 port map( B1 => n12077, B2 => n8017, C1 => n12073, C2 => 
                           n11527, A => n10899, ZN => n10894);
   U9873 : AOI221_X1 port map( B1 => n12093, B2 => n11846, C1 => n12089, C2 => 
                           n11206, A => n10898, ZN => n10895);
   U9874 : AOI221_X1 port map( B1 => n12113, B2 => n11559, C1 => n12109, C2 => 
                           n11238, A => n10897, ZN => n10896);
   U9875 : NAND4_X1 port map( A1 => n10876, A2 => n10877, A3 => n10878, A4 => 
                           n10879, ZN => n1506);
   U9876 : AOI221_X1 port map( B1 => n12077, B2 => n8018, C1 => n12073, C2 => 
                           n11528, A => n10882, ZN => n10877);
   U9877 : AOI221_X1 port map( B1 => n12093, B2 => n11847, C1 => n12089, C2 => 
                           n11207, A => n10881, ZN => n10878);
   U9878 : AOI221_X1 port map( B1 => n12113, B2 => n11560, C1 => n12109, C2 => 
                           n11239, A => n10880, ZN => n10879);
   U9879 : NAND4_X1 port map( A1 => n10859, A2 => n10860, A3 => n10861, A4 => 
                           n10862, ZN => n1508);
   U9880 : AOI221_X1 port map( B1 => n12078, B2 => n8019, C1 => n12074, C2 => 
                           n11529, A => n10865, ZN => n10860);
   U9881 : AOI221_X1 port map( B1 => n12094, B2 => n11848, C1 => n12090, C2 => 
                           n11208, A => n10864, ZN => n10861);
   U9882 : AOI221_X1 port map( B1 => n12114, B2 => n11561, C1 => n12110, C2 => 
                           n11240, A => n10863, ZN => n10862);
   U9883 : NAND4_X1 port map( A1 => n10842, A2 => n10843, A3 => n10844, A4 => 
                           n10845, ZN => n1510);
   U9884 : AOI221_X1 port map( B1 => n12078, B2 => n8020, C1 => n12074, C2 => 
                           n11530, A => n10848, ZN => n10843);
   U9885 : AOI221_X1 port map( B1 => n12094, B2 => n11849, C1 => n12090, C2 => 
                           n11209, A => n10847, ZN => n10844);
   U9886 : AOI221_X1 port map( B1 => n12114, B2 => n11562, C1 => n12110, C2 => 
                           n11241, A => n10846, ZN => n10845);
   U9887 : NAND4_X1 port map( A1 => n10825, A2 => n10826, A3 => n10827, A4 => 
                           n10828, ZN => n1512);
   U9888 : AOI221_X1 port map( B1 => n12078, B2 => n8021, C1 => n12074, C2 => 
                           n11531, A => n10831, ZN => n10826);
   U9889 : AOI221_X1 port map( B1 => n12094, B2 => n11850, C1 => n12090, C2 => 
                           n11210, A => n10830, ZN => n10827);
   U9890 : AOI221_X1 port map( B1 => n12114, B2 => n11563, C1 => n12110, C2 => 
                           n11242, A => n10829, ZN => n10828);
   U9891 : NAND4_X1 port map( A1 => n10808, A2 => n10809, A3 => n10810, A4 => 
                           n10811, ZN => n1514);
   U9892 : AOI221_X1 port map( B1 => n12078, B2 => n8022, C1 => n12074, C2 => 
                           n11532, A => n10814, ZN => n10809);
   U9893 : AOI221_X1 port map( B1 => n12094, B2 => n11851, C1 => n12090, C2 => 
                           n11211, A => n10813, ZN => n10810);
   U9894 : AOI221_X1 port map( B1 => n12114, B2 => n11564, C1 => n12110, C2 => 
                           n11243, A => n10812, ZN => n10811);
   U9895 : NAND4_X1 port map( A1 => n10791, A2 => n10792, A3 => n10793, A4 => 
                           n10794, ZN => n1516);
   U9896 : AOI221_X1 port map( B1 => n12078, B2 => n8023, C1 => n12074, C2 => 
                           n11533, A => n10797, ZN => n10792);
   U9897 : AOI221_X1 port map( B1 => n12094, B2 => n11852, C1 => n12090, C2 => 
                           n11212, A => n10796, ZN => n10793);
   U9898 : AOI221_X1 port map( B1 => n12114, B2 => n11565, C1 => n12110, C2 => 
                           n11244, A => n10795, ZN => n10794);
   U9899 : NAND4_X1 port map( A1 => n10774, A2 => n10775, A3 => n10776, A4 => 
                           n10777, ZN => n1518);
   U9900 : AOI221_X1 port map( B1 => n12078, B2 => n8024, C1 => n12074, C2 => 
                           n11534, A => n10780, ZN => n10775);
   U9901 : AOI221_X1 port map( B1 => n12094, B2 => n11853, C1 => n12090, C2 => 
                           n11213, A => n10779, ZN => n10776);
   U9902 : AOI221_X1 port map( B1 => n12114, B2 => n11566, C1 => n12110, C2 => 
                           n11245, A => n10778, ZN => n10777);
   U9903 : NAND4_X1 port map( A1 => n10757, A2 => n10758, A3 => n10759, A4 => 
                           n10760, ZN => n1520);
   U9904 : AOI221_X1 port map( B1 => n12078, B2 => n8025, C1 => n12074, C2 => 
                           n11535, A => n10763, ZN => n10758);
   U9905 : AOI221_X1 port map( B1 => n12094, B2 => n11854, C1 => n12090, C2 => 
                           n11214, A => n10762, ZN => n10759);
   U9906 : AOI221_X1 port map( B1 => n12114, B2 => n11567, C1 => n12110, C2 => 
                           n11246, A => n10761, ZN => n10760);
   U9907 : NAND4_X1 port map( A1 => n10740, A2 => n10741, A3 => n10742, A4 => 
                           n10743, ZN => n1522);
   U9908 : AOI221_X1 port map( B1 => n12078, B2 => n8026, C1 => n12074, C2 => 
                           n11536, A => n10746, ZN => n10741);
   U9909 : AOI221_X1 port map( B1 => n12094, B2 => n11855, C1 => n12090, C2 => 
                           n11215, A => n10745, ZN => n10742);
   U9910 : AOI221_X1 port map( B1 => n12114, B2 => n11568, C1 => n12110, C2 => 
                           n11247, A => n10744, ZN => n10743);
   U9911 : NAND4_X1 port map( A1 => n10723, A2 => n10724, A3 => n10725, A4 => 
                           n10726, ZN => n1524);
   U9912 : AOI221_X1 port map( B1 => n12078, B2 => n8027, C1 => n12074, C2 => 
                           n11537, A => n10729, ZN => n10724);
   U9913 : AOI221_X1 port map( B1 => n12094, B2 => n11856, C1 => n12090, C2 => 
                           n11216, A => n10728, ZN => n10725);
   U9914 : AOI221_X1 port map( B1 => n12114, B2 => n11569, C1 => n12110, C2 => 
                           n11248, A => n10727, ZN => n10726);
   U9915 : NAND4_X1 port map( A1 => n10706, A2 => n10707, A3 => n10708, A4 => 
                           n10709, ZN => n1526);
   U9916 : AOI221_X1 port map( B1 => n12078, B2 => n8028, C1 => n12074, C2 => 
                           n11538, A => n10712, ZN => n10707);
   U9917 : AOI221_X1 port map( B1 => n12094, B2 => n11857, C1 => n12090, C2 => 
                           n11217, A => n10711, ZN => n10708);
   U9918 : AOI221_X1 port map( B1 => n12114, B2 => n11570, C1 => n12110, C2 => 
                           n11249, A => n10710, ZN => n10709);
   U9919 : NAND4_X1 port map( A1 => n10689, A2 => n10690, A3 => n10691, A4 => 
                           n10692, ZN => n1528);
   U9920 : AOI221_X1 port map( B1 => n12078, B2 => n8029, C1 => n12074, C2 => 
                           n11539, A => n10695, ZN => n10690);
   U9921 : AOI221_X1 port map( B1 => n12094, B2 => n11858, C1 => n12090, C2 => 
                           n11218, A => n10694, ZN => n10691);
   U9922 : AOI221_X1 port map( B1 => n12114, B2 => n11571, C1 => n12110, C2 => 
                           n11250, A => n10693, ZN => n10692);
   U9923 : NAND4_X1 port map( A1 => n10672, A2 => n10673, A3 => n10674, A4 => 
                           n10675, ZN => n1530);
   U9924 : AOI221_X1 port map( B1 => n12078, B2 => n8030, C1 => n12074, C2 => 
                           n11540, A => n10678, ZN => n10673);
   U9925 : AOI221_X1 port map( B1 => n12094, B2 => n11859, C1 => n12090, C2 => 
                           n11219, A => n10677, ZN => n10674);
   U9926 : AOI221_X1 port map( B1 => n12114, B2 => n11572, C1 => n12110, C2 => 
                           n11251, A => n10676, ZN => n10675);
   U9927 : NAND4_X1 port map( A1 => n10655, A2 => n10656, A3 => n10657, A4 => 
                           n10658, ZN => n1532);
   U9928 : AOI221_X1 port map( B1 => n12079, B2 => n8031, C1 => n12075, C2 => 
                           n11541, A => n10661, ZN => n10656);
   U9929 : AOI221_X1 port map( B1 => n12095, B2 => n11860, C1 => n12091, C2 => 
                           n11220, A => n10660, ZN => n10657);
   U9930 : AOI221_X1 port map( B1 => n12115, B2 => n11573, C1 => n12111, C2 => 
                           n11252, A => n10659, ZN => n10658);
   U9931 : NAND4_X1 port map( A1 => n10638, A2 => n10639, A3 => n10640, A4 => 
                           n10641, ZN => n1534);
   U9932 : AOI221_X1 port map( B1 => n12079, B2 => n8032, C1 => n12075, C2 => 
                           n11542, A => n10644, ZN => n10639);
   U9933 : AOI221_X1 port map( B1 => n12095, B2 => n11861, C1 => n12091, C2 => 
                           n11221, A => n10643, ZN => n10640);
   U9934 : AOI221_X1 port map( B1 => n12115, B2 => n11574, C1 => n12111, C2 => 
                           n11253, A => n10642, ZN => n10641);
   U9935 : NAND4_X1 port map( A1 => n10621, A2 => n10622, A3 => n10623, A4 => 
                           n10624, ZN => n1536);
   U9936 : AOI221_X1 port map( B1 => n12079, B2 => n8033, C1 => n12075, C2 => 
                           n11543, A => n10627, ZN => n10622);
   U9937 : AOI221_X1 port map( B1 => n12095, B2 => n11862, C1 => n12091, C2 => 
                           n11222, A => n10626, ZN => n10623);
   U9938 : AOI221_X1 port map( B1 => n12115, B2 => n11575, C1 => n12111, C2 => 
                           n11254, A => n10625, ZN => n10624);
   U9939 : NAND4_X1 port map( A1 => n10604, A2 => n10605, A3 => n10606, A4 => 
                           n10607, ZN => n1538);
   U9940 : AOI221_X1 port map( B1 => n12079, B2 => n8034, C1 => n12075, C2 => 
                           n11544, A => n10610, ZN => n10605);
   U9941 : AOI221_X1 port map( B1 => n12095, B2 => n11863, C1 => n12091, C2 => 
                           n11223, A => n10609, ZN => n10606);
   U9942 : AOI221_X1 port map( B1 => n12115, B2 => n11576, C1 => n12111, C2 => 
                           n11255, A => n10608, ZN => n10607);
   U9943 : NAND4_X1 port map( A1 => n10587, A2 => n10588, A3 => n10589, A4 => 
                           n10590, ZN => n1540);
   U9944 : AOI221_X1 port map( B1 => n12079, B2 => n8035, C1 => n12075, C2 => 
                           n11545, A => n10593, ZN => n10588);
   U9945 : AOI221_X1 port map( B1 => n12095, B2 => n11864, C1 => n12091, C2 => 
                           n11224, A => n10592, ZN => n10589);
   U9946 : AOI221_X1 port map( B1 => n12115, B2 => n11577, C1 => n12111, C2 => 
                           n11256, A => n10591, ZN => n10590);
   U9947 : NAND4_X1 port map( A1 => n10570, A2 => n10571, A3 => n10572, A4 => 
                           n10573, ZN => n1542);
   U9948 : AOI221_X1 port map( B1 => n12079, B2 => n8036, C1 => n12075, C2 => 
                           n11546, A => n10576, ZN => n10571);
   U9949 : AOI221_X1 port map( B1 => n12095, B2 => n11865, C1 => n12091, C2 => 
                           n11225, A => n10575, ZN => n10572);
   U9950 : AOI221_X1 port map( B1 => n12115, B2 => n11578, C1 => n12111, C2 => 
                           n11257, A => n10574, ZN => n10573);
   U9951 : NAND4_X1 port map( A1 => n10553, A2 => n10554, A3 => n10555, A4 => 
                           n10556, ZN => n1544);
   U9952 : AOI221_X1 port map( B1 => n12079, B2 => n8037, C1 => n12075, C2 => 
                           n11547, A => n10559, ZN => n10554);
   U9953 : AOI221_X1 port map( B1 => n12095, B2 => n11866, C1 => n12091, C2 => 
                           n11226, A => n10558, ZN => n10555);
   U9954 : AOI221_X1 port map( B1 => n12115, B2 => n11579, C1 => n12111, C2 => 
                           n11258, A => n10557, ZN => n10556);
   U9955 : NAND4_X1 port map( A1 => n10500, A2 => n10501, A3 => n10502, A4 => 
                           n10503, ZN => n1546);
   U9956 : AOI221_X1 port map( B1 => n12079, B2 => n8038, C1 => n12075, C2 => 
                           n11548, A => n10517, ZN => n10501);
   U9957 : AOI221_X1 port map( B1 => n12095, B2 => n11867, C1 => n12091, C2 => 
                           n11227, A => n10512, ZN => n10502);
   U9958 : AOI221_X1 port map( B1 => n12115, B2 => n11580, C1 => n12111, C2 => 
                           n11259, A => n10506, ZN => n10503);
   U9959 : NAND4_X1 port map( A1 => n10463, A2 => n10464, A3 => n10465, A4 => 
                           n10466, ZN => n1548);
   U9960 : AOI221_X1 port map( B1 => n12221, B2 => n8007, C1 => n12217, C2 => 
                           n11517, A => n10479, ZN => n10464);
   U9961 : AOI221_X1 port map( B1 => n12237, B2 => n11516, C1 => n12233, C2 => 
                           n11196, A => n10474, ZN => n10465);
   U9962 : AOI221_X1 port map( B1 => n12257, B2 => n11549, C1 => n12253, C2 => 
                           n11228, A => n10467, ZN => n10466);
   U9963 : NAND4_X1 port map( A1 => n10446, A2 => n10447, A3 => n10448, A4 => 
                           n10449, ZN => n1550);
   U9964 : AOI221_X1 port map( B1 => n12221, B2 => n8008, C1 => n12217, C2 => 
                           n11518, A => n10452, ZN => n10447);
   U9965 : AOI221_X1 port map( B1 => n12237, B2 => n11837, C1 => n12233, C2 => 
                           n11197, A => n10451, ZN => n10448);
   U9966 : AOI221_X1 port map( B1 => n12257, B2 => n11550, C1 => n12253, C2 => 
                           n11229, A => n10450, ZN => n10449);
   U9967 : NAND4_X1 port map( A1 => n10429, A2 => n10430, A3 => n10431, A4 => 
                           n10432, ZN => n1552);
   U9968 : AOI221_X1 port map( B1 => n12221, B2 => n8009, C1 => n12217, C2 => 
                           n11519, A => n10435, ZN => n10430);
   U9969 : AOI221_X1 port map( B1 => n12237, B2 => n11838, C1 => n12233, C2 => 
                           n11198, A => n10434, ZN => n10431);
   U9970 : AOI221_X1 port map( B1 => n12257, B2 => n11551, C1 => n12253, C2 => 
                           n11230, A => n10433, ZN => n10432);
   U9971 : NAND4_X1 port map( A1 => n10412, A2 => n10413, A3 => n10414, A4 => 
                           n10415, ZN => n1554);
   U9972 : AOI221_X1 port map( B1 => n12221, B2 => n8010, C1 => n12217, C2 => 
                           n11520, A => n10418, ZN => n10413);
   U9973 : AOI221_X1 port map( B1 => n12237, B2 => n11839, C1 => n12233, C2 => 
                           n11199, A => n10417, ZN => n10414);
   U9974 : AOI221_X1 port map( B1 => n12257, B2 => n11552, C1 => n12253, C2 => 
                           n11231, A => n10416, ZN => n10415);
   U9975 : NAND4_X1 port map( A1 => n10395, A2 => n10396, A3 => n10397, A4 => 
                           n10398, ZN => n1556);
   U9976 : AOI221_X1 port map( B1 => n12221, B2 => n8011, C1 => n12217, C2 => 
                           n11521, A => n10401, ZN => n10396);
   U9977 : AOI221_X1 port map( B1 => n12237, B2 => n11840, C1 => n12233, C2 => 
                           n11200, A => n10400, ZN => n10397);
   U9978 : AOI221_X1 port map( B1 => n12257, B2 => n11553, C1 => n12253, C2 => 
                           n11232, A => n10399, ZN => n10398);
   U9979 : NAND4_X1 port map( A1 => n10378, A2 => n10379, A3 => n10380, A4 => 
                           n10381, ZN => n1558);
   U9980 : AOI221_X1 port map( B1 => n12221, B2 => n8012, C1 => n12217, C2 => 
                           n11522, A => n10384, ZN => n10379);
   U9981 : AOI221_X1 port map( B1 => n12237, B2 => n11841, C1 => n12233, C2 => 
                           n11201, A => n10383, ZN => n10380);
   U9982 : AOI221_X1 port map( B1 => n12257, B2 => n11554, C1 => n12253, C2 => 
                           n11233, A => n10382, ZN => n10381);
   U9983 : NAND4_X1 port map( A1 => n10361, A2 => n10362, A3 => n10363, A4 => 
                           n10364, ZN => n1560);
   U9984 : AOI221_X1 port map( B1 => n12221, B2 => n8013, C1 => n12217, C2 => 
                           n11523, A => n10367, ZN => n10362);
   U9985 : AOI221_X1 port map( B1 => n12237, B2 => n11842, C1 => n12233, C2 => 
                           n11202, A => n10366, ZN => n10363);
   U9986 : AOI221_X1 port map( B1 => n12257, B2 => n11555, C1 => n12253, C2 => 
                           n11234, A => n10365, ZN => n10364);
   U9987 : NAND4_X1 port map( A1 => n10344, A2 => n10345, A3 => n10346, A4 => 
                           n10347, ZN => n1562);
   U9988 : AOI221_X1 port map( B1 => n12221, B2 => n8014, C1 => n12217, C2 => 
                           n11524, A => n10350, ZN => n10345);
   U9989 : AOI221_X1 port map( B1 => n12237, B2 => n11843, C1 => n12233, C2 => 
                           n11203, A => n10349, ZN => n10346);
   U9990 : AOI221_X1 port map( B1 => n12257, B2 => n11556, C1 => n12253, C2 => 
                           n11235, A => n10348, ZN => n10347);
   U9991 : NAND4_X1 port map( A1 => n10327, A2 => n10328, A3 => n10329, A4 => 
                           n10330, ZN => n1564);
   U9992 : AOI221_X1 port map( B1 => n12221, B2 => n8015, C1 => n12217, C2 => 
                           n11525, A => n10333, ZN => n10328);
   U9993 : AOI221_X1 port map( B1 => n12237, B2 => n11844, C1 => n12233, C2 => 
                           n11204, A => n10332, ZN => n10329);
   U9994 : AOI221_X1 port map( B1 => n12257, B2 => n11557, C1 => n12253, C2 => 
                           n11236, A => n10331, ZN => n10330);
   U9995 : NAND4_X1 port map( A1 => n10310, A2 => n10311, A3 => n10312, A4 => 
                           n10313, ZN => n1566);
   U9996 : AOI221_X1 port map( B1 => n12221, B2 => n8016, C1 => n12217, C2 => 
                           n11526, A => n10316, ZN => n10311);
   U9997 : AOI221_X1 port map( B1 => n12237, B2 => n11845, C1 => n12233, C2 => 
                           n11205, A => n10315, ZN => n10312);
   U9998 : AOI221_X1 port map( B1 => n12257, B2 => n11558, C1 => n12253, C2 => 
                           n11237, A => n10314, ZN => n10313);
   U9999 : NAND4_X1 port map( A1 => n10293, A2 => n10294, A3 => n10295, A4 => 
                           n10296, ZN => n1568);
   U10000 : AOI221_X1 port map( B1 => n12221, B2 => n8017, C1 => n12217, C2 => 
                           n11527, A => n10299, ZN => n10294);
   U10001 : AOI221_X1 port map( B1 => n12237, B2 => n11846, C1 => n12233, C2 =>
                           n11206, A => n10298, ZN => n10295);
   U10002 : AOI221_X1 port map( B1 => n12257, B2 => n11559, C1 => n12253, C2 =>
                           n11238, A => n10297, ZN => n10296);
   U10003 : NAND4_X1 port map( A1 => n10276, A2 => n10277, A3 => n10278, A4 => 
                           n10279, ZN => n1570);
   U10004 : AOI221_X1 port map( B1 => n12221, B2 => n8018, C1 => n12217, C2 => 
                           n11528, A => n10282, ZN => n10277);
   U10005 : AOI221_X1 port map( B1 => n12237, B2 => n11847, C1 => n12233, C2 =>
                           n11207, A => n10281, ZN => n10278);
   U10006 : AOI221_X1 port map( B1 => n12257, B2 => n11560, C1 => n12253, C2 =>
                           n11239, A => n10280, ZN => n10279);
   U10007 : NAND4_X1 port map( A1 => n10259, A2 => n10260, A3 => n10261, A4 => 
                           n10262, ZN => n1572);
   U10008 : AOI221_X1 port map( B1 => n12222, B2 => n8019, C1 => n12218, C2 => 
                           n11529, A => n10265, ZN => n10260);
   U10009 : AOI221_X1 port map( B1 => n12238, B2 => n11848, C1 => n12234, C2 =>
                           n11208, A => n10264, ZN => n10261);
   U10010 : AOI221_X1 port map( B1 => n12258, B2 => n11561, C1 => n12254, C2 =>
                           n11240, A => n10263, ZN => n10262);
   U10011 : NAND4_X1 port map( A1 => n10242, A2 => n10243, A3 => n10244, A4 => 
                           n10245, ZN => n1574);
   U10012 : AOI221_X1 port map( B1 => n12222, B2 => n8020, C1 => n12218, C2 => 
                           n11530, A => n10248, ZN => n10243);
   U10013 : AOI221_X1 port map( B1 => n12238, B2 => n11849, C1 => n12234, C2 =>
                           n11209, A => n10247, ZN => n10244);
   U10014 : AOI221_X1 port map( B1 => n12258, B2 => n11562, C1 => n12254, C2 =>
                           n11241, A => n10246, ZN => n10245);
   U10015 : NAND4_X1 port map( A1 => n10225, A2 => n10226, A3 => n10227, A4 => 
                           n10228, ZN => n1576);
   U10016 : AOI221_X1 port map( B1 => n12222, B2 => n8021, C1 => n12218, C2 => 
                           n11531, A => n10231, ZN => n10226);
   U10017 : AOI221_X1 port map( B1 => n12238, B2 => n11850, C1 => n12234, C2 =>
                           n11210, A => n10230, ZN => n10227);
   U10018 : AOI221_X1 port map( B1 => n12258, B2 => n11563, C1 => n12254, C2 =>
                           n11242, A => n10229, ZN => n10228);
   U10019 : NAND4_X1 port map( A1 => n10208, A2 => n10209, A3 => n10210, A4 => 
                           n10211, ZN => n1578);
   U10020 : AOI221_X1 port map( B1 => n12222, B2 => n8022, C1 => n12218, C2 => 
                           n11532, A => n10214, ZN => n10209);
   U10021 : AOI221_X1 port map( B1 => n12238, B2 => n11851, C1 => n12234, C2 =>
                           n11211, A => n10213, ZN => n10210);
   U10022 : AOI221_X1 port map( B1 => n12258, B2 => n11564, C1 => n12254, C2 =>
                           n11243, A => n10212, ZN => n10211);
   U10023 : NAND4_X1 port map( A1 => n10191, A2 => n10192, A3 => n10193, A4 => 
                           n10194, ZN => n1580);
   U10024 : AOI221_X1 port map( B1 => n12222, B2 => n8023, C1 => n12218, C2 => 
                           n11533, A => n10197, ZN => n10192);
   U10025 : AOI221_X1 port map( B1 => n12238, B2 => n11852, C1 => n12234, C2 =>
                           n11212, A => n10196, ZN => n10193);
   U10026 : AOI221_X1 port map( B1 => n12258, B2 => n11565, C1 => n12254, C2 =>
                           n11244, A => n10195, ZN => n10194);
   U10027 : NAND4_X1 port map( A1 => n10174, A2 => n10175, A3 => n10176, A4 => 
                           n10177, ZN => n1582);
   U10028 : AOI221_X1 port map( B1 => n12222, B2 => n8024, C1 => n12218, C2 => 
                           n11534, A => n10180, ZN => n10175);
   U10029 : AOI221_X1 port map( B1 => n12238, B2 => n11853, C1 => n12234, C2 =>
                           n11213, A => n10179, ZN => n10176);
   U10030 : AOI221_X1 port map( B1 => n12258, B2 => n11566, C1 => n12254, C2 =>
                           n11245, A => n10178, ZN => n10177);
   U10031 : NAND4_X1 port map( A1 => n10157, A2 => n10158, A3 => n10159, A4 => 
                           n10160, ZN => n1584);
   U10032 : AOI221_X1 port map( B1 => n12222, B2 => n8025, C1 => n12218, C2 => 
                           n11535, A => n10163, ZN => n10158);
   U10033 : AOI221_X1 port map( B1 => n12238, B2 => n11854, C1 => n12234, C2 =>
                           n11214, A => n10162, ZN => n10159);
   U10034 : AOI221_X1 port map( B1 => n12258, B2 => n11567, C1 => n12254, C2 =>
                           n11246, A => n10161, ZN => n10160);
   U10035 : NAND4_X1 port map( A1 => n10140, A2 => n10141, A3 => n10142, A4 => 
                           n10143, ZN => n1586);
   U10036 : AOI221_X1 port map( B1 => n12222, B2 => n8026, C1 => n12218, C2 => 
                           n11536, A => n10146, ZN => n10141);
   U10037 : AOI221_X1 port map( B1 => n12238, B2 => n11855, C1 => n12234, C2 =>
                           n11215, A => n10145, ZN => n10142);
   U10038 : AOI221_X1 port map( B1 => n12258, B2 => n11568, C1 => n12254, C2 =>
                           n11247, A => n10144, ZN => n10143);
   U10039 : NAND4_X1 port map( A1 => n10123, A2 => n10124, A3 => n10125, A4 => 
                           n10126, ZN => n1588);
   U10040 : AOI221_X1 port map( B1 => n12222, B2 => n8027, C1 => n12218, C2 => 
                           n11537, A => n10129, ZN => n10124);
   U10041 : AOI221_X1 port map( B1 => n12238, B2 => n11856, C1 => n12234, C2 =>
                           n11216, A => n10128, ZN => n10125);
   U10042 : AOI221_X1 port map( B1 => n12258, B2 => n11569, C1 => n12254, C2 =>
                           n11248, A => n10127, ZN => n10126);
   U10043 : NAND4_X1 port map( A1 => n10106, A2 => n10107, A3 => n10108, A4 => 
                           n10109, ZN => n1590);
   U10044 : AOI221_X1 port map( B1 => n12222, B2 => n8028, C1 => n12218, C2 => 
                           n11538, A => n10112, ZN => n10107);
   U10045 : AOI221_X1 port map( B1 => n12238, B2 => n11857, C1 => n12234, C2 =>
                           n11217, A => n10111, ZN => n10108);
   U10046 : AOI221_X1 port map( B1 => n12258, B2 => n11570, C1 => n12254, C2 =>
                           n11249, A => n10110, ZN => n10109);
   U10047 : NAND4_X1 port map( A1 => n10089, A2 => n10090, A3 => n10091, A4 => 
                           n10092, ZN => n1592);
   U10048 : AOI221_X1 port map( B1 => n12222, B2 => n8029, C1 => n12218, C2 => 
                           n11539, A => n10095, ZN => n10090);
   U10049 : AOI221_X1 port map( B1 => n12238, B2 => n11858, C1 => n12234, C2 =>
                           n11218, A => n10094, ZN => n10091);
   U10050 : AOI221_X1 port map( B1 => n12258, B2 => n11571, C1 => n12254, C2 =>
                           n11250, A => n10093, ZN => n10092);
   U10051 : NAND4_X1 port map( A1 => n10072, A2 => n10073, A3 => n10074, A4 => 
                           n10075, ZN => n1594);
   U10052 : AOI221_X1 port map( B1 => n12222, B2 => n8030, C1 => n12218, C2 => 
                           n11540, A => n10078, ZN => n10073);
   U10053 : AOI221_X1 port map( B1 => n12238, B2 => n11859, C1 => n12234, C2 =>
                           n11219, A => n10077, ZN => n10074);
   U10054 : AOI221_X1 port map( B1 => n12258, B2 => n11572, C1 => n12254, C2 =>
                           n11251, A => n10076, ZN => n10075);
   U10055 : NAND4_X1 port map( A1 => n10055, A2 => n10056, A3 => n10057, A4 => 
                           n10058, ZN => n1596);
   U10056 : AOI221_X1 port map( B1 => n12223, B2 => n8031, C1 => n12219, C2 => 
                           n11541, A => n10061, ZN => n10056);
   U10057 : AOI221_X1 port map( B1 => n12239, B2 => n11860, C1 => n12235, C2 =>
                           n11220, A => n10060, ZN => n10057);
   U10058 : AOI221_X1 port map( B1 => n12259, B2 => n11573, C1 => n12255, C2 =>
                           n11252, A => n10059, ZN => n10058);
   U10059 : NAND4_X1 port map( A1 => n10038, A2 => n10039, A3 => n10040, A4 => 
                           n10041, ZN => n1598);
   U10060 : AOI221_X1 port map( B1 => n12223, B2 => n8032, C1 => n12219, C2 => 
                           n11542, A => n10044, ZN => n10039);
   U10061 : AOI221_X1 port map( B1 => n12239, B2 => n11861, C1 => n12235, C2 =>
                           n11221, A => n10043, ZN => n10040);
   U10062 : AOI221_X1 port map( B1 => n12259, B2 => n11574, C1 => n12255, C2 =>
                           n11253, A => n10042, ZN => n10041);
   U10063 : NAND4_X1 port map( A1 => n10021, A2 => n10022, A3 => n10023, A4 => 
                           n10024, ZN => n1600);
   U10064 : AOI221_X1 port map( B1 => n12223, B2 => n8033, C1 => n12219, C2 => 
                           n11543, A => n10027, ZN => n10022);
   U10065 : AOI221_X1 port map( B1 => n12239, B2 => n11862, C1 => n12235, C2 =>
                           n11222, A => n10026, ZN => n10023);
   U10066 : AOI221_X1 port map( B1 => n12259, B2 => n11575, C1 => n12255, C2 =>
                           n11254, A => n10025, ZN => n10024);
   U10067 : NAND4_X1 port map( A1 => n10004, A2 => n10005, A3 => n10006, A4 => 
                           n10007, ZN => n1602);
   U10068 : AOI221_X1 port map( B1 => n12223, B2 => n8034, C1 => n12219, C2 => 
                           n11544, A => n10010, ZN => n10005);
   U10069 : AOI221_X1 port map( B1 => n12239, B2 => n11863, C1 => n12235, C2 =>
                           n11223, A => n10009, ZN => n10006);
   U10070 : AOI221_X1 port map( B1 => n12259, B2 => n11576, C1 => n12255, C2 =>
                           n11255, A => n10008, ZN => n10007);
   U10071 : NAND4_X1 port map( A1 => n9987, A2 => n9988, A3 => n9989, A4 => 
                           n9990, ZN => n1604);
   U10072 : AOI221_X1 port map( B1 => n12223, B2 => n8035, C1 => n12219, C2 => 
                           n11545, A => n9993, ZN => n9988);
   U10073 : AOI221_X1 port map( B1 => n12239, B2 => n11864, C1 => n12235, C2 =>
                           n11224, A => n9992, ZN => n9989);
   U10074 : AOI221_X1 port map( B1 => n12259, B2 => n11577, C1 => n12255, C2 =>
                           n11256, A => n9991, ZN => n9990);
   U10075 : NAND4_X1 port map( A1 => n9970, A2 => n9971, A3 => n9972, A4 => 
                           n9973, ZN => n1606);
   U10076 : AOI221_X1 port map( B1 => n12223, B2 => n8036, C1 => n12219, C2 => 
                           n11546, A => n9976, ZN => n9971);
   U10077 : AOI221_X1 port map( B1 => n12239, B2 => n11865, C1 => n12235, C2 =>
                           n11225, A => n9975, ZN => n9972);
   U10078 : AOI221_X1 port map( B1 => n12259, B2 => n11578, C1 => n12255, C2 =>
                           n11257, A => n9974, ZN => n9973);
   U10079 : NAND4_X1 port map( A1 => n9953, A2 => n9954, A3 => n9955, A4 => 
                           n9956, ZN => n1608);
   U10080 : AOI221_X1 port map( B1 => n12223, B2 => n8037, C1 => n12219, C2 => 
                           n11547, A => n9959, ZN => n9954);
   U10081 : AOI221_X1 port map( B1 => n12239, B2 => n11866, C1 => n12235, C2 =>
                           n11226, A => n9958, ZN => n9955);
   U10082 : AOI221_X1 port map( B1 => n12259, B2 => n11579, C1 => n12255, C2 =>
                           n11258, A => n9957, ZN => n9956);
   U10083 : NAND4_X1 port map( A1 => n9900, A2 => n9901, A3 => n9902, A4 => 
                           n9903, ZN => n1610);
   U10084 : AOI221_X1 port map( B1 => n12223, B2 => n8038, C1 => n12219, C2 => 
                           n11548, A => n9917, ZN => n9901);
   U10085 : AOI221_X1 port map( B1 => n12239, B2 => n11867, C1 => n12235, C2 =>
                           n11227, A => n9912, ZN => n9902);
   U10086 : AOI221_X1 port map( B1 => n12259, B2 => n11580, C1 => n12255, C2 =>
                           n11259, A => n9906, ZN => n9903);
   U10087 : OAI221_X1 port map( B1 => n9309, B2 => n11993, C1 => n8861, C2 => 
                           n11989, A => n11098, ZN => n11089);
   U10088 : AOI222_X1 port map( A1 => n11985, A2 => n11709, B1 => n11982, B2 =>
                           n11388, C1 => n11978, C2 => n11260, ZN => n11098);
   U10089 : OAI221_X1 port map( B1 => n9308, B2 => n11993, C1 => n8860, C2 => 
                           n11989, A => n11062, ZN => n11055);
   U10090 : AOI222_X1 port map( A1 => n11985, A2 => n11710, B1 => n11982, B2 =>
                           n11389, C1 => n11978, C2 => n11261, ZN => n11062);
   U10091 : OAI221_X1 port map( B1 => n9307, B2 => n11993, C1 => n8859, C2 => 
                           n11989, A => n11045, ZN => n11038);
   U10092 : AOI222_X1 port map( A1 => n11985, A2 => n11711, B1 => n11982, B2 =>
                           n11390, C1 => n11978, C2 => n11262, ZN => n11045);
   U10093 : OAI221_X1 port map( B1 => n9306, B2 => n11993, C1 => n8858, C2 => 
                           n11989, A => n11028, ZN => n11021);
   U10094 : AOI222_X1 port map( A1 => n11985, A2 => n11712, B1 => n11982, B2 =>
                           n11391, C1 => n11978, C2 => n11263, ZN => n11028);
   U10095 : OAI221_X1 port map( B1 => n9305, B2 => n11993, C1 => n8857, C2 => 
                           n11989, A => n11011, ZN => n11004);
   U10096 : AOI222_X1 port map( A1 => n11985, A2 => n11713, B1 => n11982, B2 =>
                           n11392, C1 => n11978, C2 => n11264, ZN => n11011);
   U10097 : OAI221_X1 port map( B1 => n9304, B2 => n11993, C1 => n8856, C2 => 
                           n11989, A => n10994, ZN => n10987);
   U10098 : AOI222_X1 port map( A1 => n11985, A2 => n11714, B1 => n11982, B2 =>
                           n11393, C1 => n11978, C2 => n11265, ZN => n10994);
   U10099 : OAI221_X1 port map( B1 => n9303, B2 => n11993, C1 => n8855, C2 => 
                           n11989, A => n10977, ZN => n10970);
   U10100 : AOI222_X1 port map( A1 => n11985, A2 => n11715, B1 => n11982, B2 =>
                           n11394, C1 => n11978, C2 => n11266, ZN => n10977);
   U10101 : OAI221_X1 port map( B1 => n9302, B2 => n11993, C1 => n8854, C2 => 
                           n11989, A => n10960, ZN => n10953);
   U10102 : AOI222_X1 port map( A1 => n11985, A2 => n11716, B1 => n11982, B2 =>
                           n11395, C1 => n11978, C2 => n11267, ZN => n10960);
   U10103 : OAI221_X1 port map( B1 => n9301, B2 => n11993, C1 => n8853, C2 => 
                           n11989, A => n10943, ZN => n10936);
   U10104 : AOI222_X1 port map( A1 => n11985, A2 => n11717, B1 => n11981, B2 =>
                           n11396, C1 => n11977, C2 => n11268, ZN => n10943);
   U10105 : OAI221_X1 port map( B1 => n9300, B2 => n11993, C1 => n8852, C2 => 
                           n11989, A => n10926, ZN => n10919);
   U10106 : AOI222_X1 port map( A1 => n11985, A2 => n11718, B1 => n11981, B2 =>
                           n11397, C1 => n11977, C2 => n11269, ZN => n10926);
   U10107 : OAI221_X1 port map( B1 => n9299, B2 => n11993, C1 => n8851, C2 => 
                           n11989, A => n10909, ZN => n10902);
   U10108 : AOI222_X1 port map( A1 => n11985, A2 => n11719, B1 => n11981, B2 =>
                           n11398, C1 => n11977, C2 => n11270, ZN => n10909);
   U10109 : OAI221_X1 port map( B1 => n9298, B2 => n11993, C1 => n8850, C2 => 
                           n11989, A => n10892, ZN => n10885);
   U10110 : AOI222_X1 port map( A1 => n11985, A2 => n11720, B1 => n11981, B2 =>
                           n11399, C1 => n11977, C2 => n11271, ZN => n10892);
   U10111 : OAI221_X1 port map( B1 => n9297, B2 => n11994, C1 => n8849, C2 => 
                           n11990, A => n10875, ZN => n10868);
   U10112 : AOI222_X1 port map( A1 => n11986, A2 => n11721, B1 => n11981, B2 =>
                           n11400, C1 => n11977, C2 => n11272, ZN => n10875);
   U10113 : OAI221_X1 port map( B1 => n9296, B2 => n11994, C1 => n8848, C2 => 
                           n11990, A => n10858, ZN => n10851);
   U10114 : AOI222_X1 port map( A1 => n11986, A2 => n11722, B1 => n11981, B2 =>
                           n11401, C1 => n11977, C2 => n11273, ZN => n10858);
   U10115 : OAI221_X1 port map( B1 => n9295, B2 => n11994, C1 => n8847, C2 => 
                           n11990, A => n10841, ZN => n10834);
   U10116 : AOI222_X1 port map( A1 => n11986, A2 => n11723, B1 => n11981, B2 =>
                           n11402, C1 => n11977, C2 => n11274, ZN => n10841);
   U10117 : OAI221_X1 port map( B1 => n9294, B2 => n11994, C1 => n8846, C2 => 
                           n11990, A => n10824, ZN => n10817);
   U10118 : AOI222_X1 port map( A1 => n11986, A2 => n11724, B1 => n11981, B2 =>
                           n11403, C1 => n11977, C2 => n11275, ZN => n10824);
   U10119 : OAI221_X1 port map( B1 => n9293, B2 => n11994, C1 => n8845, C2 => 
                           n11990, A => n10807, ZN => n10800);
   U10120 : AOI222_X1 port map( A1 => n11986, A2 => n11725, B1 => n11981, B2 =>
                           n11404, C1 => n11977, C2 => n11276, ZN => n10807);
   U10121 : OAI221_X1 port map( B1 => n9292, B2 => n11994, C1 => n8844, C2 => 
                           n11990, A => n10790, ZN => n10783);
   U10122 : AOI222_X1 port map( A1 => n11986, A2 => n11726, B1 => n11981, B2 =>
                           n11405, C1 => n11977, C2 => n11277, ZN => n10790);
   U10123 : OAI221_X1 port map( B1 => n9291, B2 => n11994, C1 => n8843, C2 => 
                           n11990, A => n10773, ZN => n10766);
   U10124 : AOI222_X1 port map( A1 => n11986, A2 => n11727, B1 => n11981, B2 =>
                           n11406, C1 => n11977, C2 => n11278, ZN => n10773);
   U10125 : OAI221_X1 port map( B1 => n9290, B2 => n11994, C1 => n8842, C2 => 
                           n11990, A => n10756, ZN => n10749);
   U10126 : AOI222_X1 port map( A1 => n11986, A2 => n11728, B1 => n11981, B2 =>
                           n11407, C1 => n11977, C2 => n11279, ZN => n10756);
   U10127 : OAI221_X1 port map( B1 => n9289, B2 => n11994, C1 => n8841, C2 => 
                           n11990, A => n10739, ZN => n10732);
   U10128 : AOI222_X1 port map( A1 => n11986, A2 => n11729, B1 => n11980, B2 =>
                           n11408, C1 => n11976, C2 => n11280, ZN => n10739);
   U10129 : OAI221_X1 port map( B1 => n9288, B2 => n11994, C1 => n8840, C2 => 
                           n11990, A => n10722, ZN => n10715);
   U10130 : AOI222_X1 port map( A1 => n11986, A2 => n11730, B1 => n11980, B2 =>
                           n11409, C1 => n11976, C2 => n11281, ZN => n10722);
   U10131 : OAI221_X1 port map( B1 => n9287, B2 => n11994, C1 => n8839, C2 => 
                           n11990, A => n10705, ZN => n10698);
   U10132 : AOI222_X1 port map( A1 => n11986, A2 => n11731, B1 => n11980, B2 =>
                           n11410, C1 => n11976, C2 => n11282, ZN => n10705);
   U10133 : OAI221_X1 port map( B1 => n9286, B2 => n11994, C1 => n8838, C2 => 
                           n11990, A => n10688, ZN => n10681);
   U10134 : AOI222_X1 port map( A1 => n11986, A2 => n11732, B1 => n11980, B2 =>
                           n11411, C1 => n11976, C2 => n11283, ZN => n10688);
   U10135 : OAI221_X1 port map( B1 => n9285, B2 => n11995, C1 => n8837, C2 => 
                           n11991, A => n10671, ZN => n10664);
   U10136 : AOI222_X1 port map( A1 => n11987, A2 => n11733, B1 => n11980, B2 =>
                           n11412, C1 => n11976, C2 => n11284, ZN => n10671);
   U10137 : OAI221_X1 port map( B1 => n9284, B2 => n11995, C1 => n8836, C2 => 
                           n11991, A => n10654, ZN => n10647);
   U10138 : AOI222_X1 port map( A1 => n11987, A2 => n11734, B1 => n11980, B2 =>
                           n11413, C1 => n11976, C2 => n11285, ZN => n10654);
   U10139 : OAI221_X1 port map( B1 => n9283, B2 => n11995, C1 => n8835, C2 => 
                           n11991, A => n10637, ZN => n10630);
   U10140 : AOI222_X1 port map( A1 => n11987, A2 => n11735, B1 => n11980, B2 =>
                           n11414, C1 => n11976, C2 => n11286, ZN => n10637);
   U10141 : OAI221_X1 port map( B1 => n9282, B2 => n11995, C1 => n8834, C2 => 
                           n11991, A => n10620, ZN => n10613);
   U10142 : AOI222_X1 port map( A1 => n11987, A2 => n11736, B1 => n11980, B2 =>
                           n11415, C1 => n11976, C2 => n11287, ZN => n10620);
   U10143 : OAI221_X1 port map( B1 => n9281, B2 => n11995, C1 => n8833, C2 => 
                           n11991, A => n10603, ZN => n10596);
   U10144 : AOI222_X1 port map( A1 => n11987, A2 => n11737, B1 => n11980, B2 =>
                           n11416, C1 => n11976, C2 => n11288, ZN => n10603);
   U10145 : OAI221_X1 port map( B1 => n9280, B2 => n11995, C1 => n8832, C2 => 
                           n11991, A => n10586, ZN => n10579);
   U10146 : AOI222_X1 port map( A1 => n11987, A2 => n11738, B1 => n11980, B2 =>
                           n11417, C1 => n11976, C2 => n11289, ZN => n10586);
   U10147 : OAI221_X1 port map( B1 => n9279, B2 => n11995, C1 => n8831, C2 => 
                           n11991, A => n10569, ZN => n10562);
   U10148 : AOI222_X1 port map( A1 => n11987, A2 => n11739, B1 => n11980, B2 =>
                           n11418, C1 => n11976, C2 => n11290, ZN => n10569);
   U10149 : OAI221_X1 port map( B1 => n9278, B2 => n11995, C1 => n8830, C2 => 
                           n11991, A => n10548, ZN => n10526);
   U10150 : AOI222_X1 port map( A1 => n11987, A2 => n11740, B1 => n11980, B2 =>
                           n11419, C1 => n11976, C2 => n11291, ZN => n10548);
   U10151 : OAI221_X1 port map( B1 => n9309, B2 => n12137, C1 => n8861, C2 => 
                           n12133, A => n10498, ZN => n10489);
   U10152 : AOI222_X1 port map( A1 => n12129, A2 => n11709, B1 => n12126, B2 =>
                           n11388, C1 => n12122, C2 => n11260, ZN => n10498);
   U10153 : OAI221_X1 port map( B1 => n9308, B2 => n12137, C1 => n8860, C2 => 
                           n12133, A => n10462, ZN => n10455);
   U10154 : AOI222_X1 port map( A1 => n12129, A2 => n11710, B1 => n12126, B2 =>
                           n11389, C1 => n12122, C2 => n11261, ZN => n10462);
   U10155 : OAI221_X1 port map( B1 => n9307, B2 => n12137, C1 => n8859, C2 => 
                           n12133, A => n10445, ZN => n10438);
   U10156 : AOI222_X1 port map( A1 => n12129, A2 => n11711, B1 => n12126, B2 =>
                           n11390, C1 => n12122, C2 => n11262, ZN => n10445);
   U10157 : OAI221_X1 port map( B1 => n9306, B2 => n12137, C1 => n8858, C2 => 
                           n12133, A => n10428, ZN => n10421);
   U10158 : AOI222_X1 port map( A1 => n12129, A2 => n11712, B1 => n12126, B2 =>
                           n11391, C1 => n12122, C2 => n11263, ZN => n10428);
   U10159 : OAI221_X1 port map( B1 => n9305, B2 => n12137, C1 => n8857, C2 => 
                           n12133, A => n10411, ZN => n10404);
   U10160 : AOI222_X1 port map( A1 => n12129, A2 => n11713, B1 => n12126, B2 =>
                           n11392, C1 => n12122, C2 => n11264, ZN => n10411);
   U10161 : OAI221_X1 port map( B1 => n9304, B2 => n12137, C1 => n8856, C2 => 
                           n12133, A => n10394, ZN => n10387);
   U10162 : AOI222_X1 port map( A1 => n12129, A2 => n11714, B1 => n12126, B2 =>
                           n11393, C1 => n12122, C2 => n11265, ZN => n10394);
   U10163 : OAI221_X1 port map( B1 => n9303, B2 => n12137, C1 => n8855, C2 => 
                           n12133, A => n10377, ZN => n10370);
   U10164 : AOI222_X1 port map( A1 => n12129, A2 => n11715, B1 => n12126, B2 =>
                           n11394, C1 => n12122, C2 => n11266, ZN => n10377);
   U10165 : OAI221_X1 port map( B1 => n9302, B2 => n12137, C1 => n8854, C2 => 
                           n12133, A => n10360, ZN => n10353);
   U10166 : AOI222_X1 port map( A1 => n12129, A2 => n11716, B1 => n12126, B2 =>
                           n11395, C1 => n12122, C2 => n11267, ZN => n10360);
   U10167 : OAI221_X1 port map( B1 => n9301, B2 => n12137, C1 => n8853, C2 => 
                           n12133, A => n10343, ZN => n10336);
   U10168 : AOI222_X1 port map( A1 => n12129, A2 => n11717, B1 => n12125, B2 =>
                           n11396, C1 => n12121, C2 => n11268, ZN => n10343);
   U10169 : OAI221_X1 port map( B1 => n9300, B2 => n12137, C1 => n8852, C2 => 
                           n12133, A => n10326, ZN => n10319);
   U10170 : AOI222_X1 port map( A1 => n12129, A2 => n11718, B1 => n12125, B2 =>
                           n11397, C1 => n12121, C2 => n11269, ZN => n10326);
   U10171 : OAI221_X1 port map( B1 => n9299, B2 => n12137, C1 => n8851, C2 => 
                           n12133, A => n10309, ZN => n10302);
   U10172 : AOI222_X1 port map( A1 => n12129, A2 => n11719, B1 => n12125, B2 =>
                           n11398, C1 => n12121, C2 => n11270, ZN => n10309);
   U10173 : OAI221_X1 port map( B1 => n9298, B2 => n12137, C1 => n8850, C2 => 
                           n12133, A => n10292, ZN => n10285);
   U10174 : AOI222_X1 port map( A1 => n12129, A2 => n11720, B1 => n12125, B2 =>
                           n11399, C1 => n12121, C2 => n11271, ZN => n10292);
   U10175 : OAI221_X1 port map( B1 => n9297, B2 => n12138, C1 => n8849, C2 => 
                           n12134, A => n10275, ZN => n10268);
   U10176 : AOI222_X1 port map( A1 => n12130, A2 => n11721, B1 => n12125, B2 =>
                           n11400, C1 => n12121, C2 => n11272, ZN => n10275);
   U10177 : OAI221_X1 port map( B1 => n9296, B2 => n12138, C1 => n8848, C2 => 
                           n12134, A => n10258, ZN => n10251);
   U10178 : AOI222_X1 port map( A1 => n12130, A2 => n11722, B1 => n12125, B2 =>
                           n11401, C1 => n12121, C2 => n11273, ZN => n10258);
   U10179 : OAI221_X1 port map( B1 => n9295, B2 => n12138, C1 => n8847, C2 => 
                           n12134, A => n10241, ZN => n10234);
   U10180 : AOI222_X1 port map( A1 => n12130, A2 => n11723, B1 => n12125, B2 =>
                           n11402, C1 => n12121, C2 => n11274, ZN => n10241);
   U10181 : OAI221_X1 port map( B1 => n9294, B2 => n12138, C1 => n8846, C2 => 
                           n12134, A => n10224, ZN => n10217);
   U10182 : AOI222_X1 port map( A1 => n12130, A2 => n11724, B1 => n12125, B2 =>
                           n11403, C1 => n12121, C2 => n11275, ZN => n10224);
   U10183 : OAI221_X1 port map( B1 => n9293, B2 => n12138, C1 => n8845, C2 => 
                           n12134, A => n10207, ZN => n10200);
   U10184 : AOI222_X1 port map( A1 => n12130, A2 => n11725, B1 => n12125, B2 =>
                           n11404, C1 => n12121, C2 => n11276, ZN => n10207);
   U10185 : OAI221_X1 port map( B1 => n9292, B2 => n12138, C1 => n8844, C2 => 
                           n12134, A => n10190, ZN => n10183);
   U10186 : AOI222_X1 port map( A1 => n12130, A2 => n11726, B1 => n12125, B2 =>
                           n11405, C1 => n12121, C2 => n11277, ZN => n10190);
   U10187 : OAI221_X1 port map( B1 => n9291, B2 => n12138, C1 => n8843, C2 => 
                           n12134, A => n10173, ZN => n10166);
   U10188 : AOI222_X1 port map( A1 => n12130, A2 => n11727, B1 => n12125, B2 =>
                           n11406, C1 => n12121, C2 => n11278, ZN => n10173);
   U10189 : OAI221_X1 port map( B1 => n9290, B2 => n12138, C1 => n8842, C2 => 
                           n12134, A => n10156, ZN => n10149);
   U10190 : AOI222_X1 port map( A1 => n12130, A2 => n11728, B1 => n12125, B2 =>
                           n11407, C1 => n12121, C2 => n11279, ZN => n10156);
   U10191 : OAI221_X1 port map( B1 => n9289, B2 => n12138, C1 => n8841, C2 => 
                           n12134, A => n10139, ZN => n10132);
   U10192 : AOI222_X1 port map( A1 => n12130, A2 => n11729, B1 => n12124, B2 =>
                           n11408, C1 => n12120, C2 => n11280, ZN => n10139);
   U10193 : OAI221_X1 port map( B1 => n9288, B2 => n12138, C1 => n8840, C2 => 
                           n12134, A => n10122, ZN => n10115);
   U10194 : AOI222_X1 port map( A1 => n12130, A2 => n11730, B1 => n12124, B2 =>
                           n11409, C1 => n12120, C2 => n11281, ZN => n10122);
   U10195 : OAI221_X1 port map( B1 => n9287, B2 => n12138, C1 => n8839, C2 => 
                           n12134, A => n10105, ZN => n10098);
   U10196 : AOI222_X1 port map( A1 => n12130, A2 => n11731, B1 => n12124, B2 =>
                           n11410, C1 => n12120, C2 => n11282, ZN => n10105);
   U10197 : OAI221_X1 port map( B1 => n9286, B2 => n12138, C1 => n8838, C2 => 
                           n12134, A => n10088, ZN => n10081);
   U10198 : AOI222_X1 port map( A1 => n12130, A2 => n11732, B1 => n12124, B2 =>
                           n11411, C1 => n12120, C2 => n11283, ZN => n10088);
   U10199 : OAI221_X1 port map( B1 => n9285, B2 => n12139, C1 => n8837, C2 => 
                           n12135, A => n10071, ZN => n10064);
   U10200 : AOI222_X1 port map( A1 => n12131, A2 => n11733, B1 => n12124, B2 =>
                           n11412, C1 => n12120, C2 => n11284, ZN => n10071);
   U10201 : OAI221_X1 port map( B1 => n9284, B2 => n12139, C1 => n8836, C2 => 
                           n12135, A => n10054, ZN => n10047);
   U10202 : AOI222_X1 port map( A1 => n12131, A2 => n11734, B1 => n12124, B2 =>
                           n11413, C1 => n12120, C2 => n11285, ZN => n10054);
   U10203 : OAI221_X1 port map( B1 => n9283, B2 => n12139, C1 => n8835, C2 => 
                           n12135, A => n10037, ZN => n10030);
   U10204 : AOI222_X1 port map( A1 => n12131, A2 => n11735, B1 => n12124, B2 =>
                           n11414, C1 => n12120, C2 => n11286, ZN => n10037);
   U10205 : OAI221_X1 port map( B1 => n9282, B2 => n12139, C1 => n8834, C2 => 
                           n12135, A => n10020, ZN => n10013);
   U10206 : AOI222_X1 port map( A1 => n12131, A2 => n11736, B1 => n12124, B2 =>
                           n11415, C1 => n12120, C2 => n11287, ZN => n10020);
   U10207 : OAI221_X1 port map( B1 => n9281, B2 => n12139, C1 => n8833, C2 => 
                           n12135, A => n10003, ZN => n9996);
   U10208 : AOI222_X1 port map( A1 => n12131, A2 => n11737, B1 => n12124, B2 =>
                           n11416, C1 => n12120, C2 => n11288, ZN => n10003);
   U10209 : OAI221_X1 port map( B1 => n9280, B2 => n12139, C1 => n8832, C2 => 
                           n12135, A => n9986, ZN => n9979);
   U10210 : AOI222_X1 port map( A1 => n12131, A2 => n11738, B1 => n12124, B2 =>
                           n11417, C1 => n12120, C2 => n11289, ZN => n9986);
   U10211 : OAI221_X1 port map( B1 => n9279, B2 => n12139, C1 => n8831, C2 => 
                           n12135, A => n9969, ZN => n9962);
   U10212 : AOI222_X1 port map( A1 => n12131, A2 => n11739, B1 => n12124, B2 =>
                           n11418, C1 => n12120, C2 => n11290, ZN => n9969);
   U10213 : OAI221_X1 port map( B1 => n9278, B2 => n12139, C1 => n8830, C2 => 
                           n12135, A => n9948, ZN => n9926);
   U10214 : AOI222_X1 port map( A1 => n12131, A2 => n11740, B1 => n12124, B2 =>
                           n11419, C1 => n12120, C2 => n11291, ZN => n9948);
   U10215 : OAI221_X1 port map( B1 => n8957, B2 => n12045, C1 => n9213, C2 => 
                           n12041, A => n11093, ZN => n11092);
   U10216 : AOI22_X1 port map( A1 => n12037, A2 => n7879, B1 => n12034, B2 => 
                           n7975, ZN => n11093);
   U10217 : OAI221_X1 port map( B1 => n8956, B2 => n12045, C1 => n9212, C2 => 
                           n12041, A => n11059, ZN => n11058);
   U10218 : AOI22_X1 port map( A1 => n12037, A2 => n7880, B1 => n12034, B2 => 
                           n7976, ZN => n11059);
   U10219 : OAI221_X1 port map( B1 => n8955, B2 => n12045, C1 => n9211, C2 => 
                           n12041, A => n11042, ZN => n11041);
   U10220 : AOI22_X1 port map( A1 => n12037, A2 => n7881, B1 => n12034, B2 => 
                           n7977, ZN => n11042);
   U10221 : OAI221_X1 port map( B1 => n8954, B2 => n12045, C1 => n9210, C2 => 
                           n12041, A => n11025, ZN => n11024);
   U10222 : AOI22_X1 port map( A1 => n12037, A2 => n7882, B1 => n12034, B2 => 
                           n7978, ZN => n11025);
   U10223 : OAI221_X1 port map( B1 => n8953, B2 => n12045, C1 => n9209, C2 => 
                           n12041, A => n11008, ZN => n11007);
   U10224 : AOI22_X1 port map( A1 => n12037, A2 => n7883, B1 => n12034, B2 => 
                           n7979, ZN => n11008);
   U10225 : OAI221_X1 port map( B1 => n8952, B2 => n12045, C1 => n9208, C2 => 
                           n12041, A => n10991, ZN => n10990);
   U10226 : AOI22_X1 port map( A1 => n12037, A2 => n7884, B1 => n12034, B2 => 
                           n7980, ZN => n10991);
   U10227 : OAI221_X1 port map( B1 => n8951, B2 => n12045, C1 => n9207, C2 => 
                           n12041, A => n10974, ZN => n10973);
   U10228 : AOI22_X1 port map( A1 => n12037, A2 => n7885, B1 => n12034, B2 => 
                           n7981, ZN => n10974);
   U10229 : OAI221_X1 port map( B1 => n8950, B2 => n12045, C1 => n9206, C2 => 
                           n12041, A => n10957, ZN => n10956);
   U10230 : AOI22_X1 port map( A1 => n12037, A2 => n7886, B1 => n12034, B2 => 
                           n7982, ZN => n10957);
   U10231 : OAI221_X1 port map( B1 => n8949, B2 => n12045, C1 => n9205, C2 => 
                           n12041, A => n10940, ZN => n10939);
   U10232 : AOI22_X1 port map( A1 => n12037, A2 => n7887, B1 => n12033, B2 => 
                           n7983, ZN => n10940);
   U10233 : OAI221_X1 port map( B1 => n8948, B2 => n12045, C1 => n9204, C2 => 
                           n12041, A => n10923, ZN => n10922);
   U10234 : AOI22_X1 port map( A1 => n12037, A2 => n7888, B1 => n12033, B2 => 
                           n7984, ZN => n10923);
   U10235 : OAI221_X1 port map( B1 => n8947, B2 => n12045, C1 => n9203, C2 => 
                           n12041, A => n10906, ZN => n10905);
   U10236 : AOI22_X1 port map( A1 => n12037, A2 => n7889, B1 => n12033, B2 => 
                           n7985, ZN => n10906);
   U10237 : OAI221_X1 port map( B1 => n8946, B2 => n12045, C1 => n9202, C2 => 
                           n12041, A => n10889, ZN => n10888);
   U10238 : AOI22_X1 port map( A1 => n12037, A2 => n7890, B1 => n12033, B2 => 
                           n7986, ZN => n10889);
   U10239 : OAI221_X1 port map( B1 => n8945, B2 => n12046, C1 => n9201, C2 => 
                           n12042, A => n10872, ZN => n10871);
   U10240 : AOI22_X1 port map( A1 => n12038, A2 => n7891, B1 => n12033, B2 => 
                           n7987, ZN => n10872);
   U10241 : OAI221_X1 port map( B1 => n8944, B2 => n12046, C1 => n9200, C2 => 
                           n12042, A => n10855, ZN => n10854);
   U10242 : AOI22_X1 port map( A1 => n12038, A2 => n7892, B1 => n12033, B2 => 
                           n7988, ZN => n10855);
   U10243 : OAI221_X1 port map( B1 => n8943, B2 => n12046, C1 => n9199, C2 => 
                           n12042, A => n10838, ZN => n10837);
   U10244 : AOI22_X1 port map( A1 => n12038, A2 => n7893, B1 => n12033, B2 => 
                           n7989, ZN => n10838);
   U10245 : OAI221_X1 port map( B1 => n8942, B2 => n12046, C1 => n9198, C2 => 
                           n12042, A => n10821, ZN => n10820);
   U10246 : AOI22_X1 port map( A1 => n12038, A2 => n7894, B1 => n12033, B2 => 
                           n7990, ZN => n10821);
   U10247 : OAI221_X1 port map( B1 => n8941, B2 => n12046, C1 => n9197, C2 => 
                           n12042, A => n10804, ZN => n10803);
   U10248 : AOI22_X1 port map( A1 => n12038, A2 => n7895, B1 => n12033, B2 => 
                           n7991, ZN => n10804);
   U10249 : OAI221_X1 port map( B1 => n8940, B2 => n12046, C1 => n9196, C2 => 
                           n12042, A => n10787, ZN => n10786);
   U10250 : AOI22_X1 port map( A1 => n12038, A2 => n7896, B1 => n12033, B2 => 
                           n7992, ZN => n10787);
   U10251 : OAI221_X1 port map( B1 => n8939, B2 => n12046, C1 => n9195, C2 => 
                           n12042, A => n10770, ZN => n10769);
   U10252 : AOI22_X1 port map( A1 => n12038, A2 => n7897, B1 => n12033, B2 => 
                           n7993, ZN => n10770);
   U10253 : OAI221_X1 port map( B1 => n8938, B2 => n12046, C1 => n9194, C2 => 
                           n12042, A => n10753, ZN => n10752);
   U10254 : AOI22_X1 port map( A1 => n12038, A2 => n7898, B1 => n12033, B2 => 
                           n7994, ZN => n10753);
   U10255 : OAI221_X1 port map( B1 => n8937, B2 => n12046, C1 => n9193, C2 => 
                           n12042, A => n10736, ZN => n10735);
   U10256 : AOI22_X1 port map( A1 => n12038, A2 => n7899, B1 => n12032, B2 => 
                           n7995, ZN => n10736);
   U10257 : OAI221_X1 port map( B1 => n8936, B2 => n12046, C1 => n9192, C2 => 
                           n12042, A => n10719, ZN => n10718);
   U10258 : AOI22_X1 port map( A1 => n12038, A2 => n7900, B1 => n12032, B2 => 
                           n7996, ZN => n10719);
   U10259 : OAI221_X1 port map( B1 => n8935, B2 => n12046, C1 => n9191, C2 => 
                           n12042, A => n10702, ZN => n10701);
   U10260 : AOI22_X1 port map( A1 => n12038, A2 => n7901, B1 => n12032, B2 => 
                           n7997, ZN => n10702);
   U10261 : OAI221_X1 port map( B1 => n8934, B2 => n12046, C1 => n9190, C2 => 
                           n12042, A => n10685, ZN => n10684);
   U10262 : AOI22_X1 port map( A1 => n12038, A2 => n7902, B1 => n12032, B2 => 
                           n7998, ZN => n10685);
   U10263 : OAI221_X1 port map( B1 => n8933, B2 => n12047, C1 => n9189, C2 => 
                           n12043, A => n10668, ZN => n10667);
   U10264 : AOI22_X1 port map( A1 => n12039, A2 => n7903, B1 => n12032, B2 => 
                           n7999, ZN => n10668);
   U10265 : OAI221_X1 port map( B1 => n8932, B2 => n12047, C1 => n9188, C2 => 
                           n12043, A => n10651, ZN => n10650);
   U10266 : AOI22_X1 port map( A1 => n12039, A2 => n7904, B1 => n12032, B2 => 
                           n8000, ZN => n10651);
   U10267 : OAI221_X1 port map( B1 => n8931, B2 => n12047, C1 => n9187, C2 => 
                           n12043, A => n10634, ZN => n10633);
   U10268 : AOI22_X1 port map( A1 => n12039, A2 => n7905, B1 => n12032, B2 => 
                           n8001, ZN => n10634);
   U10269 : OAI221_X1 port map( B1 => n8930, B2 => n12047, C1 => n9186, C2 => 
                           n12043, A => n10617, ZN => n10616);
   U10270 : AOI22_X1 port map( A1 => n12039, A2 => n7906, B1 => n12032, B2 => 
                           n8002, ZN => n10617);
   U10271 : OAI221_X1 port map( B1 => n8929, B2 => n12047, C1 => n9185, C2 => 
                           n12043, A => n10600, ZN => n10599);
   U10272 : AOI22_X1 port map( A1 => n12039, A2 => n7907, B1 => n12032, B2 => 
                           n8003, ZN => n10600);
   U10273 : OAI221_X1 port map( B1 => n8928, B2 => n12047, C1 => n9184, C2 => 
                           n12043, A => n10583, ZN => n10582);
   U10274 : AOI22_X1 port map( A1 => n12039, A2 => n7908, B1 => n12032, B2 => 
                           n8004, ZN => n10583);
   U10275 : OAI221_X1 port map( B1 => n8927, B2 => n12047, C1 => n9183, C2 => 
                           n12043, A => n10566, ZN => n10565);
   U10276 : AOI22_X1 port map( A1 => n12039, A2 => n7909, B1 => n12032, B2 => 
                           n8005, ZN => n10566);
   U10277 : OAI221_X1 port map( B1 => n8926, B2 => n12047, C1 => n9182, C2 => 
                           n12043, A => n10532, ZN => n10529);
   U10278 : AOI22_X1 port map( A1 => n12039, A2 => n7910, B1 => n12032, B2 => 
                           n8006, ZN => n10532);
   U10279 : OAI221_X1 port map( B1 => n8957, B2 => n12189, C1 => n9213, C2 => 
                           n12185, A => n10493, ZN => n10492);
   U10280 : AOI22_X1 port map( A1 => n12181, A2 => n7879, B1 => n12178, B2 => 
                           n7975, ZN => n10493);
   U10281 : OAI221_X1 port map( B1 => n8956, B2 => n12189, C1 => n9212, C2 => 
                           n12185, A => n10459, ZN => n10458);
   U10282 : AOI22_X1 port map( A1 => n12181, A2 => n7880, B1 => n12178, B2 => 
                           n7976, ZN => n10459);
   U10283 : OAI221_X1 port map( B1 => n8955, B2 => n12189, C1 => n9211, C2 => 
                           n12185, A => n10442, ZN => n10441);
   U10284 : AOI22_X1 port map( A1 => n12181, A2 => n7881, B1 => n12178, B2 => 
                           n7977, ZN => n10442);
   U10285 : OAI221_X1 port map( B1 => n8954, B2 => n12189, C1 => n9210, C2 => 
                           n12185, A => n10425, ZN => n10424);
   U10286 : AOI22_X1 port map( A1 => n12181, A2 => n7882, B1 => n12178, B2 => 
                           n7978, ZN => n10425);
   U10287 : OAI221_X1 port map( B1 => n8953, B2 => n12189, C1 => n9209, C2 => 
                           n12185, A => n10408, ZN => n10407);
   U10288 : AOI22_X1 port map( A1 => n12181, A2 => n7883, B1 => n12178, B2 => 
                           n7979, ZN => n10408);
   U10289 : OAI221_X1 port map( B1 => n8952, B2 => n12189, C1 => n9208, C2 => 
                           n12185, A => n10391, ZN => n10390);
   U10290 : AOI22_X1 port map( A1 => n12181, A2 => n7884, B1 => n12178, B2 => 
                           n7980, ZN => n10391);
   U10291 : OAI221_X1 port map( B1 => n8951, B2 => n12189, C1 => n9207, C2 => 
                           n12185, A => n10374, ZN => n10373);
   U10292 : AOI22_X1 port map( A1 => n12181, A2 => n7885, B1 => n12178, B2 => 
                           n7981, ZN => n10374);
   U10293 : OAI221_X1 port map( B1 => n8950, B2 => n12189, C1 => n9206, C2 => 
                           n12185, A => n10357, ZN => n10356);
   U10294 : AOI22_X1 port map( A1 => n12181, A2 => n7886, B1 => n12178, B2 => 
                           n7982, ZN => n10357);
   U10295 : OAI221_X1 port map( B1 => n8949, B2 => n12189, C1 => n9205, C2 => 
                           n12185, A => n10340, ZN => n10339);
   U10296 : AOI22_X1 port map( A1 => n12181, A2 => n7887, B1 => n12177, B2 => 
                           n7983, ZN => n10340);
   U10297 : OAI221_X1 port map( B1 => n8948, B2 => n12189, C1 => n9204, C2 => 
                           n12185, A => n10323, ZN => n10322);
   U10298 : AOI22_X1 port map( A1 => n12181, A2 => n7888, B1 => n12177, B2 => 
                           n7984, ZN => n10323);
   U10299 : OAI221_X1 port map( B1 => n8947, B2 => n12189, C1 => n9203, C2 => 
                           n12185, A => n10306, ZN => n10305);
   U10300 : AOI22_X1 port map( A1 => n12181, A2 => n7889, B1 => n12177, B2 => 
                           n7985, ZN => n10306);
   U10301 : OAI221_X1 port map( B1 => n8946, B2 => n12189, C1 => n9202, C2 => 
                           n12185, A => n10289, ZN => n10288);
   U10302 : AOI22_X1 port map( A1 => n12181, A2 => n7890, B1 => n12177, B2 => 
                           n7986, ZN => n10289);
   U10303 : OAI221_X1 port map( B1 => n8945, B2 => n12190, C1 => n9201, C2 => 
                           n12186, A => n10272, ZN => n10271);
   U10304 : AOI22_X1 port map( A1 => n12182, A2 => n7891, B1 => n12177, B2 => 
                           n7987, ZN => n10272);
   U10305 : OAI221_X1 port map( B1 => n8944, B2 => n12190, C1 => n9200, C2 => 
                           n12186, A => n10255, ZN => n10254);
   U10306 : AOI22_X1 port map( A1 => n12182, A2 => n7892, B1 => n12177, B2 => 
                           n7988, ZN => n10255);
   U10307 : OAI221_X1 port map( B1 => n8943, B2 => n12190, C1 => n9199, C2 => 
                           n12186, A => n10238, ZN => n10237);
   U10308 : AOI22_X1 port map( A1 => n12182, A2 => n7893, B1 => n12177, B2 => 
                           n7989, ZN => n10238);
   U10309 : OAI221_X1 port map( B1 => n8942, B2 => n12190, C1 => n9198, C2 => 
                           n12186, A => n10221, ZN => n10220);
   U10310 : AOI22_X1 port map( A1 => n12182, A2 => n7894, B1 => n12177, B2 => 
                           n7990, ZN => n10221);
   U10311 : OAI221_X1 port map( B1 => n8941, B2 => n12190, C1 => n9197, C2 => 
                           n12186, A => n10204, ZN => n10203);
   U10312 : AOI22_X1 port map( A1 => n12182, A2 => n7895, B1 => n12177, B2 => 
                           n7991, ZN => n10204);
   U10313 : OAI221_X1 port map( B1 => n8940, B2 => n12190, C1 => n9196, C2 => 
                           n12186, A => n10187, ZN => n10186);
   U10314 : AOI22_X1 port map( A1 => n12182, A2 => n7896, B1 => n12177, B2 => 
                           n7992, ZN => n10187);
   U10315 : OAI221_X1 port map( B1 => n8939, B2 => n12190, C1 => n9195, C2 => 
                           n12186, A => n10170, ZN => n10169);
   U10316 : AOI22_X1 port map( A1 => n12182, A2 => n7897, B1 => n12177, B2 => 
                           n7993, ZN => n10170);
   U10317 : OAI221_X1 port map( B1 => n8938, B2 => n12190, C1 => n9194, C2 => 
                           n12186, A => n10153, ZN => n10152);
   U10318 : AOI22_X1 port map( A1 => n12182, A2 => n7898, B1 => n12177, B2 => 
                           n7994, ZN => n10153);
   U10319 : OAI221_X1 port map( B1 => n8937, B2 => n12190, C1 => n9193, C2 => 
                           n12186, A => n10136, ZN => n10135);
   U10320 : AOI22_X1 port map( A1 => n12182, A2 => n7899, B1 => n12176, B2 => 
                           n7995, ZN => n10136);
   U10321 : OAI221_X1 port map( B1 => n8936, B2 => n12190, C1 => n9192, C2 => 
                           n12186, A => n10119, ZN => n10118);
   U10322 : AOI22_X1 port map( A1 => n12182, A2 => n7900, B1 => n12176, B2 => 
                           n7996, ZN => n10119);
   U10323 : OAI221_X1 port map( B1 => n8935, B2 => n12190, C1 => n9191, C2 => 
                           n12186, A => n10102, ZN => n10101);
   U10324 : AOI22_X1 port map( A1 => n12182, A2 => n7901, B1 => n12176, B2 => 
                           n7997, ZN => n10102);
   U10325 : OAI221_X1 port map( B1 => n8934, B2 => n12190, C1 => n9190, C2 => 
                           n12186, A => n10085, ZN => n10084);
   U10326 : AOI22_X1 port map( A1 => n12182, A2 => n7902, B1 => n12176, B2 => 
                           n7998, ZN => n10085);
   U10327 : OAI221_X1 port map( B1 => n8933, B2 => n12191, C1 => n9189, C2 => 
                           n12187, A => n10068, ZN => n10067);
   U10328 : AOI22_X1 port map( A1 => n12183, A2 => n7903, B1 => n12176, B2 => 
                           n7999, ZN => n10068);
   U10329 : OAI221_X1 port map( B1 => n8932, B2 => n12191, C1 => n9188, C2 => 
                           n12187, A => n10051, ZN => n10050);
   U10330 : AOI22_X1 port map( A1 => n12183, A2 => n7904, B1 => n12176, B2 => 
                           n8000, ZN => n10051);
   U10331 : OAI221_X1 port map( B1 => n8931, B2 => n12191, C1 => n9187, C2 => 
                           n12187, A => n10034, ZN => n10033);
   U10332 : AOI22_X1 port map( A1 => n12183, A2 => n7905, B1 => n12176, B2 => 
                           n8001, ZN => n10034);
   U10333 : OAI221_X1 port map( B1 => n8930, B2 => n12191, C1 => n9186, C2 => 
                           n12187, A => n10017, ZN => n10016);
   U10334 : AOI22_X1 port map( A1 => n12183, A2 => n7906, B1 => n12176, B2 => 
                           n8002, ZN => n10017);
   U10335 : OAI221_X1 port map( B1 => n8929, B2 => n12191, C1 => n9185, C2 => 
                           n12187, A => n10000, ZN => n9999);
   U10336 : AOI22_X1 port map( A1 => n12183, A2 => n7907, B1 => n12176, B2 => 
                           n8003, ZN => n10000);
   U10337 : OAI221_X1 port map( B1 => n8928, B2 => n12191, C1 => n9184, C2 => 
                           n12187, A => n9983, ZN => n9982);
   U10338 : AOI22_X1 port map( A1 => n12183, A2 => n7908, B1 => n12176, B2 => 
                           n8004, ZN => n9983);
   U10339 : OAI221_X1 port map( B1 => n8927, B2 => n12191, C1 => n9183, C2 => 
                           n12187, A => n9966, ZN => n9965);
   U10340 : AOI22_X1 port map( A1 => n12183, A2 => n7909, B1 => n12176, B2 => 
                           n8005, ZN => n9966);
   U10341 : OAI221_X1 port map( B1 => n8926, B2 => n12191, C1 => n9182, C2 => 
                           n12187, A => n9932, ZN => n9929);
   U10342 : AOI22_X1 port map( A1 => n12183, A2 => n7910, B1 => n12176, B2 => 
                           n8006, ZN => n9932);
   U10343 : AOI22_X1 port map( A1 => n12001, A2 => n11324, B1 => n11998, B2 => 
                           n11484, ZN => n11097);
   U10344 : AOI22_X1 port map( A1 => n12001, A2 => n11325, B1 => n11998, B2 => 
                           n11485, ZN => n11061);
   U10345 : AOI22_X1 port map( A1 => n12001, A2 => n11326, B1 => n11998, B2 => 
                           n11486, ZN => n11044);
   U10346 : AOI22_X1 port map( A1 => n12001, A2 => n11327, B1 => n11998, B2 => 
                           n11487, ZN => n11027);
   U10347 : AOI22_X1 port map( A1 => n12001, A2 => n11328, B1 => n11998, B2 => 
                           n11488, ZN => n11010);
   U10348 : AOI22_X1 port map( A1 => n12001, A2 => n11329, B1 => n11998, B2 => 
                           n11489, ZN => n10993);
   U10349 : AOI22_X1 port map( A1 => n12001, A2 => n11330, B1 => n11998, B2 => 
                           n11490, ZN => n10976);
   U10350 : AOI22_X1 port map( A1 => n12001, A2 => n11331, B1 => n11998, B2 => 
                           n11491, ZN => n10959);
   U10351 : AOI22_X1 port map( A1 => n12001, A2 => n11332, B1 => n11997, B2 => 
                           n11492, ZN => n10942);
   U10352 : AOI22_X1 port map( A1 => n12001, A2 => n11333, B1 => n11997, B2 => 
                           n11493, ZN => n10925);
   U10353 : AOI22_X1 port map( A1 => n12001, A2 => n11334, B1 => n11997, B2 => 
                           n11494, ZN => n10908);
   U10354 : AOI22_X1 port map( A1 => n12001, A2 => n11335, B1 => n11997, B2 => 
                           n11495, ZN => n10891);
   U10355 : AOI22_X1 port map( A1 => n12002, A2 => n11336, B1 => n11997, B2 => 
                           n11496, ZN => n10874);
   U10356 : AOI22_X1 port map( A1 => n12002, A2 => n11337, B1 => n11997, B2 => 
                           n11497, ZN => n10857);
   U10357 : AOI22_X1 port map( A1 => n12002, A2 => n11338, B1 => n11997, B2 => 
                           n11498, ZN => n10840);
   U10358 : AOI22_X1 port map( A1 => n12002, A2 => n11339, B1 => n11997, B2 => 
                           n11499, ZN => n10823);
   U10359 : AOI22_X1 port map( A1 => n12002, A2 => n11340, B1 => n11997, B2 => 
                           n11500, ZN => n10806);
   U10360 : AOI22_X1 port map( A1 => n12002, A2 => n11341, B1 => n11997, B2 => 
                           n11501, ZN => n10789);
   U10361 : AOI22_X1 port map( A1 => n12002, A2 => n11342, B1 => n11997, B2 => 
                           n11502, ZN => n10772);
   U10362 : AOI22_X1 port map( A1 => n12002, A2 => n11343, B1 => n11997, B2 => 
                           n11503, ZN => n10755);
   U10363 : AOI22_X1 port map( A1 => n12002, A2 => n11344, B1 => n11996, B2 => 
                           n11504, ZN => n10738);
   U10364 : AOI22_X1 port map( A1 => n12002, A2 => n11345, B1 => n11996, B2 => 
                           n11505, ZN => n10721);
   U10365 : AOI22_X1 port map( A1 => n12002, A2 => n11346, B1 => n11996, B2 => 
                           n11506, ZN => n10704);
   U10366 : AOI22_X1 port map( A1 => n12002, A2 => n11347, B1 => n11996, B2 => 
                           n11507, ZN => n10687);
   U10367 : AOI22_X1 port map( A1 => n12003, A2 => n11348, B1 => n11996, B2 => 
                           n11508, ZN => n10670);
   U10368 : AOI22_X1 port map( A1 => n12003, A2 => n11349, B1 => n11996, B2 => 
                           n11509, ZN => n10653);
   U10369 : AOI22_X1 port map( A1 => n12003, A2 => n11350, B1 => n11996, B2 => 
                           n11510, ZN => n10636);
   U10370 : AOI22_X1 port map( A1 => n12003, A2 => n11351, B1 => n11996, B2 => 
                           n11511, ZN => n10619);
   U10371 : AOI22_X1 port map( A1 => n12003, A2 => n11352, B1 => n11996, B2 => 
                           n11512, ZN => n10602);
   U10372 : AOI22_X1 port map( A1 => n12003, A2 => n11353, B1 => n11996, B2 => 
                           n11513, ZN => n10585);
   U10373 : AOI22_X1 port map( A1 => n12003, A2 => n11354, B1 => n11996, B2 => 
                           n11514, ZN => n10568);
   U10374 : AOI22_X1 port map( A1 => n12003, A2 => n11355, B1 => n11996, B2 => 
                           n11515, ZN => n10543);
   U10375 : AOI22_X1 port map( A1 => n12145, A2 => n11324, B1 => n12142, B2 => 
                           n11484, ZN => n10497);
   U10376 : AOI22_X1 port map( A1 => n12145, A2 => n11325, B1 => n12142, B2 => 
                           n11485, ZN => n10461);
   U10377 : AOI22_X1 port map( A1 => n12145, A2 => n11326, B1 => n12142, B2 => 
                           n11486, ZN => n10444);
   U10378 : AOI22_X1 port map( A1 => n12145, A2 => n11327, B1 => n12142, B2 => 
                           n11487, ZN => n10427);
   U10379 : AOI22_X1 port map( A1 => n12145, A2 => n11328, B1 => n12142, B2 => 
                           n11488, ZN => n10410);
   U10380 : AOI22_X1 port map( A1 => n12145, A2 => n11329, B1 => n12142, B2 => 
                           n11489, ZN => n10393);
   U10381 : AOI22_X1 port map( A1 => n12145, A2 => n11330, B1 => n12142, B2 => 
                           n11490, ZN => n10376);
   U10382 : AOI22_X1 port map( A1 => n12145, A2 => n11331, B1 => n12142, B2 => 
                           n11491, ZN => n10359);
   U10383 : AOI22_X1 port map( A1 => n12145, A2 => n11332, B1 => n12141, B2 => 
                           n11492, ZN => n10342);
   U10384 : AOI22_X1 port map( A1 => n12145, A2 => n11333, B1 => n12141, B2 => 
                           n11493, ZN => n10325);
   U10385 : AOI22_X1 port map( A1 => n12145, A2 => n11334, B1 => n12141, B2 => 
                           n11494, ZN => n10308);
   U10386 : AOI22_X1 port map( A1 => n12145, A2 => n11335, B1 => n12141, B2 => 
                           n11495, ZN => n10291);
   U10387 : AOI22_X1 port map( A1 => n12146, A2 => n11336, B1 => n12141, B2 => 
                           n11496, ZN => n10274);
   U10388 : AOI22_X1 port map( A1 => n12146, A2 => n11337, B1 => n12141, B2 => 
                           n11497, ZN => n10257);
   U10389 : AOI22_X1 port map( A1 => n12146, A2 => n11338, B1 => n12141, B2 => 
                           n11498, ZN => n10240);
   U10390 : AOI22_X1 port map( A1 => n12146, A2 => n11339, B1 => n12141, B2 => 
                           n11499, ZN => n10223);
   U10391 : AOI22_X1 port map( A1 => n12146, A2 => n11340, B1 => n12141, B2 => 
                           n11500, ZN => n10206);
   U10392 : AOI22_X1 port map( A1 => n12146, A2 => n11341, B1 => n12141, B2 => 
                           n11501, ZN => n10189);
   U10393 : AOI22_X1 port map( A1 => n12146, A2 => n11342, B1 => n12141, B2 => 
                           n11502, ZN => n10172);
   U10394 : AOI22_X1 port map( A1 => n12146, A2 => n11343, B1 => n12141, B2 => 
                           n11503, ZN => n10155);
   U10395 : AOI22_X1 port map( A1 => n12146, A2 => n11344, B1 => n12140, B2 => 
                           n11504, ZN => n10138);
   U10396 : AOI22_X1 port map( A1 => n12146, A2 => n11345, B1 => n12140, B2 => 
                           n11505, ZN => n10121);
   U10397 : AOI22_X1 port map( A1 => n12146, A2 => n11346, B1 => n12140, B2 => 
                           n11506, ZN => n10104);
   U10398 : AOI22_X1 port map( A1 => n12146, A2 => n11347, B1 => n12140, B2 => 
                           n11507, ZN => n10087);
   U10399 : AOI22_X1 port map( A1 => n12147, A2 => n11348, B1 => n12140, B2 => 
                           n11508, ZN => n10070);
   U10400 : AOI22_X1 port map( A1 => n12147, A2 => n11349, B1 => n12140, B2 => 
                           n11509, ZN => n10053);
   U10401 : AOI22_X1 port map( A1 => n12147, A2 => n11350, B1 => n12140, B2 => 
                           n11510, ZN => n10036);
   U10402 : AOI22_X1 port map( A1 => n12147, A2 => n11351, B1 => n12140, B2 => 
                           n11511, ZN => n10019);
   U10403 : AOI22_X1 port map( A1 => n12147, A2 => n11352, B1 => n12140, B2 => 
                           n11512, ZN => n10002);
   U10404 : AOI22_X1 port map( A1 => n12147, A2 => n11353, B1 => n12140, B2 => 
                           n11513, ZN => n9985);
   U10405 : AOI22_X1 port map( A1 => n12147, A2 => n11354, B1 => n12140, B2 => 
                           n11514, ZN => n9968);
   U10406 : AOI22_X1 port map( A1 => n12147, A2 => n11355, B1 => n12140, B2 => 
                           n11515, ZN => n9943);
   U10407 : OAI22_X1 port map( A1 => n11890, A2 => n12388, B1 => n12277, B2 => 
                           n9693, ZN => n1739);
   U10408 : OAI22_X1 port map( A1 => n11890, A2 => n12392, B1 => n12277, B2 => 
                           n9692, ZN => n1740);
   U10409 : OAI22_X1 port map( A1 => n11890, A2 => n12396, B1 => n12277, B2 => 
                           n9691, ZN => n1741);
   U10410 : OAI22_X1 port map( A1 => n11890, A2 => n12400, B1 => n12277, B2 => 
                           n9690, ZN => n1742);
   U10411 : OAI22_X1 port map( A1 => n11890, A2 => n12404, B1 => n12277, B2 => 
                           n9689, ZN => n1743);
   U10412 : OAI22_X1 port map( A1 => n11890, A2 => n12408, B1 => n12277, B2 => 
                           n9688, ZN => n1744);
   U10413 : OAI22_X1 port map( A1 => n11890, A2 => n12412, B1 => n12277, B2 => 
                           n9687, ZN => n1745);
   U10414 : OAI22_X1 port map( A1 => n11890, A2 => n12416, B1 => n12277, B2 => 
                           n9686, ZN => n1746);
   U10415 : OAI22_X1 port map( A1 => n11889, A2 => n12420, B1 => n12277, B2 => 
                           n9685, ZN => n1747);
   U10416 : OAI22_X1 port map( A1 => n11889, A2 => n12424, B1 => n12277, B2 => 
                           n9684, ZN => n1748);
   U10417 : OAI22_X1 port map( A1 => n11889, A2 => n12428, B1 => n12277, B2 => 
                           n9683, ZN => n1749);
   U10418 : OAI22_X1 port map( A1 => n11889, A2 => n12432, B1 => n12277, B2 => 
                           n9682, ZN => n1750);
   U10419 : OAI22_X1 port map( A1 => n11889, A2 => n12436, B1 => n9894, B2 => 
                           n9681, ZN => n1751);
   U10420 : OAI22_X1 port map( A1 => n11889, A2 => n12440, B1 => n9894, B2 => 
                           n9680, ZN => n1752);
   U10421 : OAI22_X1 port map( A1 => n11889, A2 => n12444, B1 => n9894, B2 => 
                           n9679, ZN => n1753);
   U10422 : OAI22_X1 port map( A1 => n11889, A2 => n12448, B1 => n12277, B2 => 
                           n9678, ZN => n1754);
   U10423 : OAI22_X1 port map( A1 => n11889, A2 => n12452, B1 => n12277, B2 => 
                           n9677, ZN => n1755);
   U10424 : OAI22_X1 port map( A1 => n11889, A2 => n12456, B1 => n12277, B2 => 
                           n9676, ZN => n1756);
   U10425 : OAI22_X1 port map( A1 => n11889, A2 => n12460, B1 => n12277, B2 => 
                           n9675, ZN => n1757);
   U10426 : OAI22_X1 port map( A1 => n11889, A2 => n12464, B1 => n12277, B2 => 
                           n9674, ZN => n1758);
   U10427 : OAI22_X1 port map( A1 => n11888, A2 => n12468, B1 => n12277, B2 => 
                           n9673, ZN => n1759);
   U10428 : OAI22_X1 port map( A1 => n11888, A2 => n12472, B1 => n12277, B2 => 
                           n9672, ZN => n1760);
   U10429 : OAI22_X1 port map( A1 => n11888, A2 => n12476, B1 => n12277, B2 => 
                           n9671, ZN => n1761);
   U10430 : OAI22_X1 port map( A1 => n11888, A2 => n12480, B1 => n12277, B2 => 
                           n9670, ZN => n1762);
   U10431 : OAI22_X1 port map( A1 => n11888, A2 => n12484, B1 => n9894, B2 => 
                           n9669, ZN => n1763);
   U10432 : OAI22_X1 port map( A1 => n11888, A2 => n12488, B1 => n9894, B2 => 
                           n9668, ZN => n1764);
   U10433 : OAI22_X1 port map( A1 => n11888, A2 => n12492, B1 => n9894, B2 => 
                           n9667, ZN => n1765);
   U10434 : OAI22_X1 port map( A1 => n11888, A2 => n12496, B1 => n9894, B2 => 
                           n9666, ZN => n1766);
   U10435 : OAI22_X1 port map( A1 => n11888, A2 => n12500, B1 => n9894, B2 => 
                           n9665, ZN => n1767);
   U10436 : OAI22_X1 port map( A1 => n11888, A2 => n12504, B1 => n9894, B2 => 
                           n9664, ZN => n1768);
   U10437 : OAI22_X1 port map( A1 => n11888, A2 => n12508, B1 => n9894, B2 => 
                           n9663, ZN => n1769);
   U10438 : OAI22_X1 port map( A1 => n11888, A2 => n12516, B1 => n9894, B2 => 
                           n9662, ZN => n1770);
   U10439 : OAI22_X1 port map( A1 => n11896, A2 => n12388, B1 => n12285, B2 => 
                           n9629, ZN => n1803);
   U10440 : OAI22_X1 port map( A1 => n11896, A2 => n12392, B1 => n12285, B2 => 
                           n9628, ZN => n1804);
   U10441 : OAI22_X1 port map( A1 => n11896, A2 => n12396, B1 => n12285, B2 => 
                           n9627, ZN => n1805);
   U10442 : OAI22_X1 port map( A1 => n11896, A2 => n12400, B1 => n12285, B2 => 
                           n9626, ZN => n1806);
   U10443 : OAI22_X1 port map( A1 => n11896, A2 => n12404, B1 => n12285, B2 => 
                           n9625, ZN => n1807);
   U10444 : OAI22_X1 port map( A1 => n11896, A2 => n12408, B1 => n12285, B2 => 
                           n9624, ZN => n1808);
   U10445 : OAI22_X1 port map( A1 => n11896, A2 => n12412, B1 => n12285, B2 => 
                           n9623, ZN => n1809);
   U10446 : OAI22_X1 port map( A1 => n11896, A2 => n12416, B1 => n12285, B2 => 
                           n9622, ZN => n1810);
   U10447 : OAI22_X1 port map( A1 => n11895, A2 => n12420, B1 => n12285, B2 => 
                           n9621, ZN => n1811);
   U10448 : OAI22_X1 port map( A1 => n11895, A2 => n12424, B1 => n12285, B2 => 
                           n9620, ZN => n1812);
   U10449 : OAI22_X1 port map( A1 => n11895, A2 => n12428, B1 => n12285, B2 => 
                           n9619, ZN => n1813);
   U10450 : OAI22_X1 port map( A1 => n11895, A2 => n12432, B1 => n12285, B2 => 
                           n9618, ZN => n1814);
   U10451 : OAI22_X1 port map( A1 => n11895, A2 => n12436, B1 => n9892, B2 => 
                           n9617, ZN => n1815);
   U10452 : OAI22_X1 port map( A1 => n11895, A2 => n12440, B1 => n9892, B2 => 
                           n9616, ZN => n1816);
   U10453 : OAI22_X1 port map( A1 => n11895, A2 => n12444, B1 => n9892, B2 => 
                           n9615, ZN => n1817);
   U10454 : OAI22_X1 port map( A1 => n11895, A2 => n12448, B1 => n12285, B2 => 
                           n9614, ZN => n1818);
   U10455 : OAI22_X1 port map( A1 => n11895, A2 => n12452, B1 => n12285, B2 => 
                           n9613, ZN => n1819);
   U10456 : OAI22_X1 port map( A1 => n11895, A2 => n12456, B1 => n12285, B2 => 
                           n9612, ZN => n1820);
   U10457 : OAI22_X1 port map( A1 => n11895, A2 => n12460, B1 => n12285, B2 => 
                           n9611, ZN => n1821);
   U10458 : OAI22_X1 port map( A1 => n11895, A2 => n12464, B1 => n12285, B2 => 
                           n9610, ZN => n1822);
   U10459 : OAI22_X1 port map( A1 => n11894, A2 => n12468, B1 => n12285, B2 => 
                           n9609, ZN => n1823);
   U10460 : OAI22_X1 port map( A1 => n11894, A2 => n12472, B1 => n12285, B2 => 
                           n9608, ZN => n1824);
   U10461 : OAI22_X1 port map( A1 => n11894, A2 => n12476, B1 => n12285, B2 => 
                           n9607, ZN => n1825);
   U10462 : OAI22_X1 port map( A1 => n11894, A2 => n12480, B1 => n12285, B2 => 
                           n9606, ZN => n1826);
   U10463 : OAI22_X1 port map( A1 => n11894, A2 => n12484, B1 => n9892, B2 => 
                           n9605, ZN => n1827);
   U10464 : OAI22_X1 port map( A1 => n11894, A2 => n12488, B1 => n9892, B2 => 
                           n9604, ZN => n1828);
   U10465 : OAI22_X1 port map( A1 => n11894, A2 => n12492, B1 => n9892, B2 => 
                           n9603, ZN => n1829);
   U10466 : OAI22_X1 port map( A1 => n11894, A2 => n12496, B1 => n9892, B2 => 
                           n9602, ZN => n1830);
   U10467 : OAI22_X1 port map( A1 => n11894, A2 => n12500, B1 => n9892, B2 => 
                           n9601, ZN => n1831);
   U10468 : OAI22_X1 port map( A1 => n11894, A2 => n12504, B1 => n9892, B2 => 
                           n9600, ZN => n1832);
   U10469 : OAI22_X1 port map( A1 => n11894, A2 => n12508, B1 => n9892, B2 => 
                           n9599, ZN => n1833);
   U10470 : OAI22_X1 port map( A1 => n11894, A2 => n12516, B1 => n9892, B2 => 
                           n9598, ZN => n1834);
   U10471 : OAI22_X1 port map( A1 => n11914, A2 => n12387, B1 => n12309, B2 => 
                           n9437, ZN => n1995);
   U10472 : OAI22_X1 port map( A1 => n11914, A2 => n12391, B1 => n12309, B2 => 
                           n9436, ZN => n1996);
   U10473 : OAI22_X1 port map( A1 => n11914, A2 => n12395, B1 => n12309, B2 => 
                           n9435, ZN => n1997);
   U10474 : OAI22_X1 port map( A1 => n11914, A2 => n12399, B1 => n12309, B2 => 
                           n9434, ZN => n1998);
   U10475 : OAI22_X1 port map( A1 => n11914, A2 => n12403, B1 => n12309, B2 => 
                           n9433, ZN => n1999);
   U10476 : OAI22_X1 port map( A1 => n11914, A2 => n12407, B1 => n12309, B2 => 
                           n9432, ZN => n2000);
   U10477 : OAI22_X1 port map( A1 => n11914, A2 => n12411, B1 => n12309, B2 => 
                           n9431, ZN => n2001);
   U10478 : OAI22_X1 port map( A1 => n11914, A2 => n12415, B1 => n12309, B2 => 
                           n9430, ZN => n2002);
   U10479 : OAI22_X1 port map( A1 => n11913, A2 => n12419, B1 => n12309, B2 => 
                           n9429, ZN => n2003);
   U10480 : OAI22_X1 port map( A1 => n11913, A2 => n12423, B1 => n12309, B2 => 
                           n9428, ZN => n2004);
   U10481 : OAI22_X1 port map( A1 => n11913, A2 => n12427, B1 => n12309, B2 => 
                           n9427, ZN => n2005);
   U10482 : OAI22_X1 port map( A1 => n11913, A2 => n12431, B1 => n12309, B2 => 
                           n9426, ZN => n2006);
   U10483 : OAI22_X1 port map( A1 => n11913, A2 => n12435, B1 => n9883, B2 => 
                           n9425, ZN => n2007);
   U10484 : OAI22_X1 port map( A1 => n11913, A2 => n12439, B1 => n9883, B2 => 
                           n9424, ZN => n2008);
   U10485 : OAI22_X1 port map( A1 => n11913, A2 => n12443, B1 => n9883, B2 => 
                           n9423, ZN => n2009);
   U10486 : OAI22_X1 port map( A1 => n11913, A2 => n12447, B1 => n12309, B2 => 
                           n9422, ZN => n2010);
   U10487 : OAI22_X1 port map( A1 => n11913, A2 => n12451, B1 => n12309, B2 => 
                           n9421, ZN => n2011);
   U10488 : OAI22_X1 port map( A1 => n11913, A2 => n12455, B1 => n12309, B2 => 
                           n9420, ZN => n2012);
   U10489 : OAI22_X1 port map( A1 => n11913, A2 => n12459, B1 => n12309, B2 => 
                           n9419, ZN => n2013);
   U10490 : OAI22_X1 port map( A1 => n11913, A2 => n12463, B1 => n12309, B2 => 
                           n9418, ZN => n2014);
   U10491 : OAI22_X1 port map( A1 => n11912, A2 => n12467, B1 => n12309, B2 => 
                           n9417, ZN => n2015);
   U10492 : OAI22_X1 port map( A1 => n11912, A2 => n12471, B1 => n12309, B2 => 
                           n9416, ZN => n2016);
   U10493 : OAI22_X1 port map( A1 => n11912, A2 => n12475, B1 => n12309, B2 => 
                           n9415, ZN => n2017);
   U10494 : OAI22_X1 port map( A1 => n11912, A2 => n12479, B1 => n12309, B2 => 
                           n9414, ZN => n2018);
   U10495 : OAI22_X1 port map( A1 => n11912, A2 => n12483, B1 => n9883, B2 => 
                           n9413, ZN => n2019);
   U10496 : OAI22_X1 port map( A1 => n11912, A2 => n12487, B1 => n9883, B2 => 
                           n9412, ZN => n2020);
   U10497 : OAI22_X1 port map( A1 => n11912, A2 => n12491, B1 => n9883, B2 => 
                           n9411, ZN => n2021);
   U10498 : OAI22_X1 port map( A1 => n11912, A2 => n12495, B1 => n9883, B2 => 
                           n9410, ZN => n2022);
   U10499 : OAI22_X1 port map( A1 => n11912, A2 => n12499, B1 => n9883, B2 => 
                           n9409, ZN => n2023);
   U10500 : OAI22_X1 port map( A1 => n11912, A2 => n12503, B1 => n9883, B2 => 
                           n9408, ZN => n2024);
   U10501 : OAI22_X1 port map( A1 => n11912, A2 => n12507, B1 => n9883, B2 => 
                           n9407, ZN => n2025);
   U10502 : OAI22_X1 port map( A1 => n11912, A2 => n12515, B1 => n9883, B2 => 
                           n9406, ZN => n2026);
   U10503 : OAI22_X1 port map( A1 => n11908, A2 => n12387, B1 => n12301, B2 => 
                           n9501, ZN => n1931);
   U10504 : OAI22_X1 port map( A1 => n11908, A2 => n12391, B1 => n12301, B2 => 
                           n9500, ZN => n1932);
   U10505 : OAI22_X1 port map( A1 => n11908, A2 => n12395, B1 => n12301, B2 => 
                           n9499, ZN => n1933);
   U10506 : OAI22_X1 port map( A1 => n11908, A2 => n12399, B1 => n12301, B2 => 
                           n9498, ZN => n1934);
   U10507 : OAI22_X1 port map( A1 => n11908, A2 => n12403, B1 => n12301, B2 => 
                           n9497, ZN => n1935);
   U10508 : OAI22_X1 port map( A1 => n11908, A2 => n12407, B1 => n12301, B2 => 
                           n9496, ZN => n1936);
   U10509 : OAI22_X1 port map( A1 => n11908, A2 => n12411, B1 => n12301, B2 => 
                           n9495, ZN => n1937);
   U10510 : OAI22_X1 port map( A1 => n11908, A2 => n12415, B1 => n12301, B2 => 
                           n9494, ZN => n1938);
   U10511 : OAI22_X1 port map( A1 => n11907, A2 => n12419, B1 => n12301, B2 => 
                           n9493, ZN => n1939);
   U10512 : OAI22_X1 port map( A1 => n11907, A2 => n12423, B1 => n12301, B2 => 
                           n9492, ZN => n1940);
   U10513 : OAI22_X1 port map( A1 => n11907, A2 => n12427, B1 => n12301, B2 => 
                           n9491, ZN => n1941);
   U10514 : OAI22_X1 port map( A1 => n11907, A2 => n12431, B1 => n12301, B2 => 
                           n9490, ZN => n1942);
   U10515 : OAI22_X1 port map( A1 => n11907, A2 => n12435, B1 => n9887, B2 => 
                           n9489, ZN => n1943);
   U10516 : OAI22_X1 port map( A1 => n11907, A2 => n12439, B1 => n9887, B2 => 
                           n9488, ZN => n1944);
   U10517 : OAI22_X1 port map( A1 => n11907, A2 => n12443, B1 => n9887, B2 => 
                           n9487, ZN => n1945);
   U10518 : OAI22_X1 port map( A1 => n11907, A2 => n12447, B1 => n12301, B2 => 
                           n9486, ZN => n1946);
   U10519 : OAI22_X1 port map( A1 => n11907, A2 => n12451, B1 => n12301, B2 => 
                           n9485, ZN => n1947);
   U10520 : OAI22_X1 port map( A1 => n11907, A2 => n12455, B1 => n12301, B2 => 
                           n9484, ZN => n1948);
   U10521 : OAI22_X1 port map( A1 => n11907, A2 => n12459, B1 => n12301, B2 => 
                           n9483, ZN => n1949);
   U10522 : OAI22_X1 port map( A1 => n11907, A2 => n12463, B1 => n12301, B2 => 
                           n9482, ZN => n1950);
   U10523 : OAI22_X1 port map( A1 => n11906, A2 => n12467, B1 => n12301, B2 => 
                           n9481, ZN => n1951);
   U10524 : OAI22_X1 port map( A1 => n11906, A2 => n12471, B1 => n12301, B2 => 
                           n9480, ZN => n1952);
   U10525 : OAI22_X1 port map( A1 => n11906, A2 => n12475, B1 => n12301, B2 => 
                           n9479, ZN => n1953);
   U10526 : OAI22_X1 port map( A1 => n11906, A2 => n12479, B1 => n12301, B2 => 
                           n9478, ZN => n1954);
   U10527 : OAI22_X1 port map( A1 => n11906, A2 => n12483, B1 => n9887, B2 => 
                           n9477, ZN => n1955);
   U10528 : OAI22_X1 port map( A1 => n11906, A2 => n12487, B1 => n9887, B2 => 
                           n9476, ZN => n1956);
   U10529 : OAI22_X1 port map( A1 => n11906, A2 => n12491, B1 => n9887, B2 => 
                           n9475, ZN => n1957);
   U10530 : OAI22_X1 port map( A1 => n11906, A2 => n12495, B1 => n9887, B2 => 
                           n9474, ZN => n1958);
   U10531 : OAI22_X1 port map( A1 => n11906, A2 => n12499, B1 => n9887, B2 => 
                           n9473, ZN => n1959);
   U10532 : OAI22_X1 port map( A1 => n11906, A2 => n12503, B1 => n9887, B2 => 
                           n9472, ZN => n1960);
   U10533 : OAI22_X1 port map( A1 => n11906, A2 => n12507, B1 => n9887, B2 => 
                           n9471, ZN => n1961);
   U10534 : OAI22_X1 port map( A1 => n11906, A2 => n12515, B1 => n9887, B2 => 
                           n9470, ZN => n1962);
   U10535 : OAI22_X1 port map( A1 => n11944, A2 => n12386, B1 => n12349, B2 => 
                           n9117, ZN => n2315);
   U10536 : OAI22_X1 port map( A1 => n11944, A2 => n12390, B1 => n12349, B2 => 
                           n9116, ZN => n2316);
   U10537 : OAI22_X1 port map( A1 => n11944, A2 => n12394, B1 => n12349, B2 => 
                           n9115, ZN => n2317);
   U10538 : OAI22_X1 port map( A1 => n11944, A2 => n12398, B1 => n12349, B2 => 
                           n9114, ZN => n2318);
   U10539 : OAI22_X1 port map( A1 => n11944, A2 => n12402, B1 => n12349, B2 => 
                           n9113, ZN => n2319);
   U10540 : OAI22_X1 port map( A1 => n11944, A2 => n12406, B1 => n12349, B2 => 
                           n9112, ZN => n2320);
   U10541 : OAI22_X1 port map( A1 => n11944, A2 => n12410, B1 => n12349, B2 => 
                           n9111, ZN => n2321);
   U10542 : OAI22_X1 port map( A1 => n11944, A2 => n12414, B1 => n12349, B2 => 
                           n9110, ZN => n2322);
   U10543 : OAI22_X1 port map( A1 => n11943, A2 => n12418, B1 => n12349, B2 => 
                           n9109, ZN => n2323);
   U10544 : OAI22_X1 port map( A1 => n11943, A2 => n12422, B1 => n12349, B2 => 
                           n9108, ZN => n2324);
   U10545 : OAI22_X1 port map( A1 => n11943, A2 => n12426, B1 => n12349, B2 => 
                           n9107, ZN => n2325);
   U10546 : OAI22_X1 port map( A1 => n11943, A2 => n12430, B1 => n12349, B2 => 
                           n9106, ZN => n2326);
   U10547 : OAI22_X1 port map( A1 => n11943, A2 => n12434, B1 => n9871, B2 => 
                           n9105, ZN => n2327);
   U10548 : OAI22_X1 port map( A1 => n11943, A2 => n12438, B1 => n9871, B2 => 
                           n9104, ZN => n2328);
   U10549 : OAI22_X1 port map( A1 => n11943, A2 => n12442, B1 => n9871, B2 => 
                           n9103, ZN => n2329);
   U10550 : OAI22_X1 port map( A1 => n11943, A2 => n12446, B1 => n12349, B2 => 
                           n9102, ZN => n2330);
   U10551 : OAI22_X1 port map( A1 => n11943, A2 => n12450, B1 => n12349, B2 => 
                           n9101, ZN => n2331);
   U10552 : OAI22_X1 port map( A1 => n11943, A2 => n12454, B1 => n12349, B2 => 
                           n9100, ZN => n2332);
   U10553 : OAI22_X1 port map( A1 => n11943, A2 => n12458, B1 => n12349, B2 => 
                           n9099, ZN => n2333);
   U10554 : OAI22_X1 port map( A1 => n11943, A2 => n12462, B1 => n12349, B2 => 
                           n9098, ZN => n2334);
   U10555 : OAI22_X1 port map( A1 => n11942, A2 => n12466, B1 => n12349, B2 => 
                           n9097, ZN => n2335);
   U10556 : OAI22_X1 port map( A1 => n11942, A2 => n12470, B1 => n12349, B2 => 
                           n9096, ZN => n2336);
   U10557 : OAI22_X1 port map( A1 => n11942, A2 => n12474, B1 => n12349, B2 => 
                           n9095, ZN => n2337);
   U10558 : OAI22_X1 port map( A1 => n11942, A2 => n12478, B1 => n12349, B2 => 
                           n9094, ZN => n2338);
   U10559 : OAI22_X1 port map( A1 => n11942, A2 => n12482, B1 => n9871, B2 => 
                           n9093, ZN => n2339);
   U10560 : OAI22_X1 port map( A1 => n11942, A2 => n12486, B1 => n9871, B2 => 
                           n9092, ZN => n2340);
   U10561 : OAI22_X1 port map( A1 => n11942, A2 => n12490, B1 => n9871, B2 => 
                           n9091, ZN => n2341);
   U10562 : OAI22_X1 port map( A1 => n11942, A2 => n12494, B1 => n9871, B2 => 
                           n9090, ZN => n2342);
   U10563 : OAI22_X1 port map( A1 => n11942, A2 => n12498, B1 => n9871, B2 => 
                           n9089, ZN => n2343);
   U10564 : OAI22_X1 port map( A1 => n11942, A2 => n12502, B1 => n9871, B2 => 
                           n9088, ZN => n2344);
   U10565 : OAI22_X1 port map( A1 => n11942, A2 => n12506, B1 => n9871, B2 => 
                           n9087, ZN => n2345);
   U10566 : OAI22_X1 port map( A1 => n11942, A2 => n12514, B1 => n9871, B2 => 
                           n9086, ZN => n2346);
   U10567 : OAI22_X1 port map( A1 => n11902, A2 => n12387, B1 => n12293, B2 => 
                           n9565, ZN => n1867);
   U10568 : OAI22_X1 port map( A1 => n11902, A2 => n12391, B1 => n12293, B2 => 
                           n9564, ZN => n1868);
   U10569 : OAI22_X1 port map( A1 => n11902, A2 => n12395, B1 => n12293, B2 => 
                           n9563, ZN => n1869);
   U10570 : OAI22_X1 port map( A1 => n11902, A2 => n12399, B1 => n12293, B2 => 
                           n9562, ZN => n1870);
   U10571 : OAI22_X1 port map( A1 => n11902, A2 => n12403, B1 => n12293, B2 => 
                           n9561, ZN => n1871);
   U10572 : OAI22_X1 port map( A1 => n11902, A2 => n12407, B1 => n12293, B2 => 
                           n9560, ZN => n1872);
   U10573 : OAI22_X1 port map( A1 => n11902, A2 => n12411, B1 => n12293, B2 => 
                           n9559, ZN => n1873);
   U10574 : OAI22_X1 port map( A1 => n11902, A2 => n12415, B1 => n12293, B2 => 
                           n9558, ZN => n1874);
   U10575 : OAI22_X1 port map( A1 => n11901, A2 => n12419, B1 => n12293, B2 => 
                           n9557, ZN => n1875);
   U10576 : OAI22_X1 port map( A1 => n11901, A2 => n12423, B1 => n12293, B2 => 
                           n9556, ZN => n1876);
   U10577 : OAI22_X1 port map( A1 => n11901, A2 => n12427, B1 => n12293, B2 => 
                           n9555, ZN => n1877);
   U10578 : OAI22_X1 port map( A1 => n11901, A2 => n12431, B1 => n12293, B2 => 
                           n9554, ZN => n1878);
   U10579 : OAI22_X1 port map( A1 => n11901, A2 => n12435, B1 => n9889, B2 => 
                           n9553, ZN => n1879);
   U10580 : OAI22_X1 port map( A1 => n11901, A2 => n12439, B1 => n9889, B2 => 
                           n9552, ZN => n1880);
   U10581 : OAI22_X1 port map( A1 => n11901, A2 => n12443, B1 => n9889, B2 => 
                           n9551, ZN => n1881);
   U10582 : OAI22_X1 port map( A1 => n11901, A2 => n12447, B1 => n12293, B2 => 
                           n9550, ZN => n1882);
   U10583 : OAI22_X1 port map( A1 => n11901, A2 => n12451, B1 => n12293, B2 => 
                           n9549, ZN => n1883);
   U10584 : OAI22_X1 port map( A1 => n11901, A2 => n12455, B1 => n12293, B2 => 
                           n9548, ZN => n1884);
   U10585 : OAI22_X1 port map( A1 => n11901, A2 => n12459, B1 => n12293, B2 => 
                           n9547, ZN => n1885);
   U10586 : OAI22_X1 port map( A1 => n11901, A2 => n12463, B1 => n12293, B2 => 
                           n9546, ZN => n1886);
   U10587 : OAI22_X1 port map( A1 => n11900, A2 => n12467, B1 => n12293, B2 => 
                           n9545, ZN => n1887);
   U10588 : OAI22_X1 port map( A1 => n11900, A2 => n12471, B1 => n12293, B2 => 
                           n9544, ZN => n1888);
   U10589 : OAI22_X1 port map( A1 => n11900, A2 => n12475, B1 => n12293, B2 => 
                           n9543, ZN => n1889);
   U10590 : OAI22_X1 port map( A1 => n11900, A2 => n12479, B1 => n12293, B2 => 
                           n9542, ZN => n1890);
   U10591 : OAI22_X1 port map( A1 => n11900, A2 => n12483, B1 => n9889, B2 => 
                           n9541, ZN => n1891);
   U10592 : OAI22_X1 port map( A1 => n11900, A2 => n12487, B1 => n9889, B2 => 
                           n9540, ZN => n1892);
   U10593 : OAI22_X1 port map( A1 => n11900, A2 => n12491, B1 => n9889, B2 => 
                           n9539, ZN => n1893);
   U10594 : OAI22_X1 port map( A1 => n11900, A2 => n12495, B1 => n9889, B2 => 
                           n9538, ZN => n1894);
   U10595 : OAI22_X1 port map( A1 => n11900, A2 => n12499, B1 => n9889, B2 => 
                           n9537, ZN => n1895);
   U10596 : OAI22_X1 port map( A1 => n11900, A2 => n12503, B1 => n9889, B2 => 
                           n9536, ZN => n1896);
   U10597 : OAI22_X1 port map( A1 => n11900, A2 => n12507, B1 => n9889, B2 => 
                           n9535, ZN => n1897);
   U10598 : OAI22_X1 port map( A1 => n11900, A2 => n12515, B1 => n9889, B2 => 
                           n9534, ZN => n1898);
   U10599 : OAI22_X1 port map( A1 => n11971, A2 => n12386, B1 => n12509, B2 => 
                           n8829, ZN => n2603);
   U10600 : OAI22_X1 port map( A1 => n11971, A2 => n12390, B1 => n12509, B2 => 
                           n8828, ZN => n2604);
   U10601 : OAI22_X1 port map( A1 => n11971, A2 => n12394, B1 => n12509, B2 => 
                           n8827, ZN => n2605);
   U10602 : OAI22_X1 port map( A1 => n11971, A2 => n12398, B1 => n12509, B2 => 
                           n8826, ZN => n2606);
   U10603 : OAI22_X1 port map( A1 => n11971, A2 => n12402, B1 => n12509, B2 => 
                           n8825, ZN => n2607);
   U10604 : OAI22_X1 port map( A1 => n11971, A2 => n12406, B1 => n12509, B2 => 
                           n8824, ZN => n2608);
   U10605 : OAI22_X1 port map( A1 => n11971, A2 => n12410, B1 => n12509, B2 => 
                           n8823, ZN => n2609);
   U10606 : OAI22_X1 port map( A1 => n11971, A2 => n12414, B1 => n12509, B2 => 
                           n8822, ZN => n2610);
   U10607 : OAI22_X1 port map( A1 => n11970, A2 => n12418, B1 => n12509, B2 => 
                           n8821, ZN => n2611);
   U10608 : OAI22_X1 port map( A1 => n11970, A2 => n12422, B1 => n12509, B2 => 
                           n8820, ZN => n2612);
   U10609 : OAI22_X1 port map( A1 => n11970, A2 => n12426, B1 => n12509, B2 => 
                           n8819, ZN => n2613);
   U10610 : OAI22_X1 port map( A1 => n11970, A2 => n12430, B1 => n12509, B2 => 
                           n8818, ZN => n2614);
   U10611 : OAI22_X1 port map( A1 => n11970, A2 => n12434, B1 => n9823, B2 => 
                           n8817, ZN => n2615);
   U10612 : OAI22_X1 port map( A1 => n11970, A2 => n12438, B1 => n9823, B2 => 
                           n8816, ZN => n2616);
   U10613 : OAI22_X1 port map( A1 => n11970, A2 => n12442, B1 => n9823, B2 => 
                           n8815, ZN => n2617);
   U10614 : OAI22_X1 port map( A1 => n11970, A2 => n12446, B1 => n12509, B2 => 
                           n8814, ZN => n2618);
   U10615 : OAI22_X1 port map( A1 => n11970, A2 => n12450, B1 => n12509, B2 => 
                           n8813, ZN => n2619);
   U10616 : OAI22_X1 port map( A1 => n11970, A2 => n12454, B1 => n12509, B2 => 
                           n8812, ZN => n2620);
   U10617 : OAI22_X1 port map( A1 => n11970, A2 => n12458, B1 => n12509, B2 => 
                           n8811, ZN => n2621);
   U10618 : OAI22_X1 port map( A1 => n11970, A2 => n12462, B1 => n12509, B2 => 
                           n8810, ZN => n2622);
   U10619 : OAI22_X1 port map( A1 => n11969, A2 => n12466, B1 => n12509, B2 => 
                           n8809, ZN => n2623);
   U10620 : OAI22_X1 port map( A1 => n11969, A2 => n12470, B1 => n12509, B2 => 
                           n8808, ZN => n2624);
   U10621 : OAI22_X1 port map( A1 => n11969, A2 => n12474, B1 => n12509, B2 => 
                           n8807, ZN => n2625);
   U10622 : OAI22_X1 port map( A1 => n11969, A2 => n12478, B1 => n12509, B2 => 
                           n8806, ZN => n2626);
   U10623 : OAI22_X1 port map( A1 => n11969, A2 => n12482, B1 => n9823, B2 => 
                           n8805, ZN => n2627);
   U10624 : OAI22_X1 port map( A1 => n11969, A2 => n12486, B1 => n9823, B2 => 
                           n8804, ZN => n2628);
   U10625 : OAI22_X1 port map( A1 => n11969, A2 => n12490, B1 => n9823, B2 => 
                           n8803, ZN => n2629);
   U10626 : OAI22_X1 port map( A1 => n11969, A2 => n12494, B1 => n9823, B2 => 
                           n8802, ZN => n2630);
   U10627 : OAI22_X1 port map( A1 => n11969, A2 => n12498, B1 => n9823, B2 => 
                           n8801, ZN => n2631);
   U10628 : OAI22_X1 port map( A1 => n11969, A2 => n12502, B1 => n9823, B2 => 
                           n8800, ZN => n2632);
   U10629 : OAI22_X1 port map( A1 => n11969, A2 => n12506, B1 => n9823, B2 => 
                           n8799, ZN => n2633);
   U10630 : OAI22_X1 port map( A1 => n11969, A2 => n12514, B1 => n9823, B2 => 
                           n8798, ZN => n2634);
   U10631 : OAI22_X1 port map( A1 => n11941, A2 => n12386, B1 => n12345, B2 => 
                           n9149, ZN => n2283);
   U10632 : OAI22_X1 port map( A1 => n11941, A2 => n12390, B1 => n12345, B2 => 
                           n9148, ZN => n2284);
   U10633 : OAI22_X1 port map( A1 => n11941, A2 => n12394, B1 => n12345, B2 => 
                           n9147, ZN => n2285);
   U10634 : OAI22_X1 port map( A1 => n11941, A2 => n12398, B1 => n12345, B2 => 
                           n9146, ZN => n2286);
   U10635 : OAI22_X1 port map( A1 => n11941, A2 => n12402, B1 => n12345, B2 => 
                           n9145, ZN => n2287);
   U10636 : OAI22_X1 port map( A1 => n11941, A2 => n12406, B1 => n12345, B2 => 
                           n9144, ZN => n2288);
   U10637 : OAI22_X1 port map( A1 => n11941, A2 => n12410, B1 => n12345, B2 => 
                           n9143, ZN => n2289);
   U10638 : OAI22_X1 port map( A1 => n11941, A2 => n12414, B1 => n12345, B2 => 
                           n9142, ZN => n2290);
   U10639 : OAI22_X1 port map( A1 => n11940, A2 => n12418, B1 => n12345, B2 => 
                           n9141, ZN => n2291);
   U10640 : OAI22_X1 port map( A1 => n11940, A2 => n12422, B1 => n12345, B2 => 
                           n9140, ZN => n2292);
   U10641 : OAI22_X1 port map( A1 => n11940, A2 => n12426, B1 => n12345, B2 => 
                           n9139, ZN => n2293);
   U10642 : OAI22_X1 port map( A1 => n11940, A2 => n12430, B1 => n12345, B2 => 
                           n9138, ZN => n2294);
   U10643 : OAI22_X1 port map( A1 => n11940, A2 => n12434, B1 => n9872, B2 => 
                           n9137, ZN => n2295);
   U10644 : OAI22_X1 port map( A1 => n11940, A2 => n12438, B1 => n9872, B2 => 
                           n9136, ZN => n2296);
   U10645 : OAI22_X1 port map( A1 => n11940, A2 => n12442, B1 => n9872, B2 => 
                           n9135, ZN => n2297);
   U10646 : OAI22_X1 port map( A1 => n11940, A2 => n12446, B1 => n12345, B2 => 
                           n9134, ZN => n2298);
   U10647 : OAI22_X1 port map( A1 => n11940, A2 => n12450, B1 => n12345, B2 => 
                           n9133, ZN => n2299);
   U10648 : OAI22_X1 port map( A1 => n11940, A2 => n12454, B1 => n12345, B2 => 
                           n9132, ZN => n2300);
   U10649 : OAI22_X1 port map( A1 => n11940, A2 => n12458, B1 => n12345, B2 => 
                           n9131, ZN => n2301);
   U10650 : OAI22_X1 port map( A1 => n11940, A2 => n12462, B1 => n12345, B2 => 
                           n9130, ZN => n2302);
   U10651 : OAI22_X1 port map( A1 => n11939, A2 => n12466, B1 => n12345, B2 => 
                           n9129, ZN => n2303);
   U10652 : OAI22_X1 port map( A1 => n11939, A2 => n12470, B1 => n12345, B2 => 
                           n9128, ZN => n2304);
   U10653 : OAI22_X1 port map( A1 => n11939, A2 => n12474, B1 => n12345, B2 => 
                           n9127, ZN => n2305);
   U10654 : OAI22_X1 port map( A1 => n11939, A2 => n12478, B1 => n12345, B2 => 
                           n9126, ZN => n2306);
   U10655 : OAI22_X1 port map( A1 => n11939, A2 => n12482, B1 => n9872, B2 => 
                           n9125, ZN => n2307);
   U10656 : OAI22_X1 port map( A1 => n11939, A2 => n12486, B1 => n9872, B2 => 
                           n9124, ZN => n2308);
   U10657 : OAI22_X1 port map( A1 => n11939, A2 => n12490, B1 => n9872, B2 => 
                           n9123, ZN => n2309);
   U10658 : OAI22_X1 port map( A1 => n11939, A2 => n12494, B1 => n9872, B2 => 
                           n9122, ZN => n2310);
   U10659 : OAI22_X1 port map( A1 => n11939, A2 => n12498, B1 => n9872, B2 => 
                           n9121, ZN => n2311);
   U10660 : OAI22_X1 port map( A1 => n11939, A2 => n12502, B1 => n9872, B2 => 
                           n9120, ZN => n2312);
   U10661 : OAI22_X1 port map( A1 => n11939, A2 => n12506, B1 => n9872, B2 => 
                           n9119, ZN => n2313);
   U10662 : OAI22_X1 port map( A1 => n11939, A2 => n12514, B1 => n9872, B2 => 
                           n9118, ZN => n2314);
   U10663 : OAI22_X1 port map( A1 => n11956, A2 => n12386, B1 => n12365, B2 => 
                           n8989, ZN => n2443);
   U10664 : OAI22_X1 port map( A1 => n11956, A2 => n12390, B1 => n12365, B2 => 
                           n8988, ZN => n2444);
   U10665 : OAI22_X1 port map( A1 => n11956, A2 => n12394, B1 => n12365, B2 => 
                           n8987, ZN => n2445);
   U10666 : OAI22_X1 port map( A1 => n11956, A2 => n12398, B1 => n12365, B2 => 
                           n8986, ZN => n2446);
   U10667 : OAI22_X1 port map( A1 => n11956, A2 => n12402, B1 => n12365, B2 => 
                           n8985, ZN => n2447);
   U10668 : OAI22_X1 port map( A1 => n11956, A2 => n12406, B1 => n12365, B2 => 
                           n8984, ZN => n2448);
   U10669 : OAI22_X1 port map( A1 => n11956, A2 => n12410, B1 => n12365, B2 => 
                           n8983, ZN => n2449);
   U10670 : OAI22_X1 port map( A1 => n11956, A2 => n12414, B1 => n12365, B2 => 
                           n8982, ZN => n2450);
   U10671 : OAI22_X1 port map( A1 => n11955, A2 => n12418, B1 => n12365, B2 => 
                           n8981, ZN => n2451);
   U10672 : OAI22_X1 port map( A1 => n11955, A2 => n12422, B1 => n12365, B2 => 
                           n8980, ZN => n2452);
   U10673 : OAI22_X1 port map( A1 => n11955, A2 => n12426, B1 => n12365, B2 => 
                           n8979, ZN => n2453);
   U10674 : OAI22_X1 port map( A1 => n11955, A2 => n12430, B1 => n12365, B2 => 
                           n8978, ZN => n2454);
   U10675 : OAI22_X1 port map( A1 => n11955, A2 => n12434, B1 => n9866, B2 => 
                           n8977, ZN => n2455);
   U10676 : OAI22_X1 port map( A1 => n11955, A2 => n12438, B1 => n9866, B2 => 
                           n8976, ZN => n2456);
   U10677 : OAI22_X1 port map( A1 => n11955, A2 => n12442, B1 => n9866, B2 => 
                           n8975, ZN => n2457);
   U10678 : OAI22_X1 port map( A1 => n11955, A2 => n12446, B1 => n12365, B2 => 
                           n8974, ZN => n2458);
   U10679 : OAI22_X1 port map( A1 => n11955, A2 => n12450, B1 => n12365, B2 => 
                           n8973, ZN => n2459);
   U10680 : OAI22_X1 port map( A1 => n11955, A2 => n12454, B1 => n12365, B2 => 
                           n8972, ZN => n2460);
   U10681 : OAI22_X1 port map( A1 => n11955, A2 => n12458, B1 => n12365, B2 => 
                           n8971, ZN => n2461);
   U10682 : OAI22_X1 port map( A1 => n11955, A2 => n12462, B1 => n12365, B2 => 
                           n8970, ZN => n2462);
   U10683 : OAI22_X1 port map( A1 => n11954, A2 => n12466, B1 => n12365, B2 => 
                           n8969, ZN => n2463);
   U10684 : OAI22_X1 port map( A1 => n11954, A2 => n12470, B1 => n12365, B2 => 
                           n8968, ZN => n2464);
   U10685 : OAI22_X1 port map( A1 => n11954, A2 => n12474, B1 => n12365, B2 => 
                           n8967, ZN => n2465);
   U10686 : OAI22_X1 port map( A1 => n11954, A2 => n12478, B1 => n12365, B2 => 
                           n8966, ZN => n2466);
   U10687 : OAI22_X1 port map( A1 => n11954, A2 => n12482, B1 => n9866, B2 => 
                           n8965, ZN => n2467);
   U10688 : OAI22_X1 port map( A1 => n11954, A2 => n12486, B1 => n9866, B2 => 
                           n8964, ZN => n2468);
   U10689 : OAI22_X1 port map( A1 => n11954, A2 => n12490, B1 => n9866, B2 => 
                           n8963, ZN => n2469);
   U10690 : OAI22_X1 port map( A1 => n11954, A2 => n12494, B1 => n9866, B2 => 
                           n8962, ZN => n2470);
   U10691 : OAI22_X1 port map( A1 => n11954, A2 => n12498, B1 => n9866, B2 => 
                           n8961, ZN => n2471);
   U10692 : OAI22_X1 port map( A1 => n11954, A2 => n12502, B1 => n9866, B2 => 
                           n8960, ZN => n2472);
   U10693 : OAI22_X1 port map( A1 => n11954, A2 => n12506, B1 => n9866, B2 => 
                           n8959, ZN => n2473);
   U10694 : OAI22_X1 port map( A1 => n11954, A2 => n12514, B1 => n9866, B2 => 
                           n8958, ZN => n2474);
   U10695 : OAI22_X1 port map( A1 => n11932, A2 => n12387, B1 => n12333, B2 => 
                           n9245, ZN => n2187);
   U10696 : OAI22_X1 port map( A1 => n11932, A2 => n12391, B1 => n12333, B2 => 
                           n9244, ZN => n2188);
   U10697 : OAI22_X1 port map( A1 => n11932, A2 => n12395, B1 => n12333, B2 => 
                           n9243, ZN => n2189);
   U10698 : OAI22_X1 port map( A1 => n11932, A2 => n12399, B1 => n12333, B2 => 
                           n9242, ZN => n2190);
   U10699 : OAI22_X1 port map( A1 => n11932, A2 => n12403, B1 => n12333, B2 => 
                           n9241, ZN => n2191);
   U10700 : OAI22_X1 port map( A1 => n11932, A2 => n12407, B1 => n12333, B2 => 
                           n9240, ZN => n2192);
   U10701 : OAI22_X1 port map( A1 => n11932, A2 => n12411, B1 => n12333, B2 => 
                           n9239, ZN => n2193);
   U10702 : OAI22_X1 port map( A1 => n11932, A2 => n12415, B1 => n12333, B2 => 
                           n9238, ZN => n2194);
   U10703 : OAI22_X1 port map( A1 => n11931, A2 => n12419, B1 => n12333, B2 => 
                           n9237, ZN => n2195);
   U10704 : OAI22_X1 port map( A1 => n11931, A2 => n12423, B1 => n12333, B2 => 
                           n9236, ZN => n2196);
   U10705 : OAI22_X1 port map( A1 => n11931, A2 => n12427, B1 => n12333, B2 => 
                           n9235, ZN => n2197);
   U10706 : OAI22_X1 port map( A1 => n11931, A2 => n12431, B1 => n12333, B2 => 
                           n9234, ZN => n2198);
   U10707 : OAI22_X1 port map( A1 => n11931, A2 => n12435, B1 => n9876, B2 => 
                           n9233, ZN => n2199);
   U10708 : OAI22_X1 port map( A1 => n11931, A2 => n12439, B1 => n9876, B2 => 
                           n9232, ZN => n2200);
   U10709 : OAI22_X1 port map( A1 => n11931, A2 => n12443, B1 => n9876, B2 => 
                           n9231, ZN => n2201);
   U10710 : OAI22_X1 port map( A1 => n11931, A2 => n12447, B1 => n12333, B2 => 
                           n9230, ZN => n2202);
   U10711 : OAI22_X1 port map( A1 => n11931, A2 => n12451, B1 => n12333, B2 => 
                           n9229, ZN => n2203);
   U10712 : OAI22_X1 port map( A1 => n11931, A2 => n12455, B1 => n12333, B2 => 
                           n9228, ZN => n2204);
   U10713 : OAI22_X1 port map( A1 => n11931, A2 => n12459, B1 => n12333, B2 => 
                           n9227, ZN => n2205);
   U10714 : OAI22_X1 port map( A1 => n11931, A2 => n12463, B1 => n12333, B2 => 
                           n9226, ZN => n2206);
   U10715 : OAI22_X1 port map( A1 => n11930, A2 => n12467, B1 => n12333, B2 => 
                           n9225, ZN => n2207);
   U10716 : OAI22_X1 port map( A1 => n11930, A2 => n12471, B1 => n12333, B2 => 
                           n9224, ZN => n2208);
   U10717 : OAI22_X1 port map( A1 => n11930, A2 => n12475, B1 => n12333, B2 => 
                           n9223, ZN => n2209);
   U10718 : OAI22_X1 port map( A1 => n11930, A2 => n12479, B1 => n12333, B2 => 
                           n9222, ZN => n2210);
   U10719 : OAI22_X1 port map( A1 => n11930, A2 => n12483, B1 => n9876, B2 => 
                           n9221, ZN => n2211);
   U10720 : OAI22_X1 port map( A1 => n11930, A2 => n12487, B1 => n9876, B2 => 
                           n9220, ZN => n2212);
   U10721 : OAI22_X1 port map( A1 => n11930, A2 => n12491, B1 => n9876, B2 => 
                           n9219, ZN => n2213);
   U10722 : OAI22_X1 port map( A1 => n11930, A2 => n12495, B1 => n9876, B2 => 
                           n9218, ZN => n2214);
   U10723 : OAI22_X1 port map( A1 => n11930, A2 => n12499, B1 => n9876, B2 => 
                           n9217, ZN => n2215);
   U10724 : OAI22_X1 port map( A1 => n11930, A2 => n12503, B1 => n9876, B2 => 
                           n9216, ZN => n2216);
   U10725 : OAI22_X1 port map( A1 => n11930, A2 => n12507, B1 => n9876, B2 => 
                           n9215, ZN => n2217);
   U10726 : OAI22_X1 port map( A1 => n11930, A2 => n12515, B1 => n9876, B2 => 
                           n9214, ZN => n2218);
   U10727 : OAI22_X1 port map( A1 => n11953, A2 => n12386, B1 => n12361, B2 => 
                           n9021, ZN => n2411);
   U10728 : OAI22_X1 port map( A1 => n11953, A2 => n12390, B1 => n12361, B2 => 
                           n9020, ZN => n2412);
   U10729 : OAI22_X1 port map( A1 => n11953, A2 => n12394, B1 => n12361, B2 => 
                           n9019, ZN => n2413);
   U10730 : OAI22_X1 port map( A1 => n11953, A2 => n12398, B1 => n12361, B2 => 
                           n9018, ZN => n2414);
   U10731 : OAI22_X1 port map( A1 => n11953, A2 => n12402, B1 => n12361, B2 => 
                           n9017, ZN => n2415);
   U10732 : OAI22_X1 port map( A1 => n11953, A2 => n12406, B1 => n12361, B2 => 
                           n9016, ZN => n2416);
   U10733 : OAI22_X1 port map( A1 => n11953, A2 => n12410, B1 => n12361, B2 => 
                           n9015, ZN => n2417);
   U10734 : OAI22_X1 port map( A1 => n11953, A2 => n12414, B1 => n12361, B2 => 
                           n9014, ZN => n2418);
   U10735 : OAI22_X1 port map( A1 => n11952, A2 => n12418, B1 => n12361, B2 => 
                           n9013, ZN => n2419);
   U10736 : OAI22_X1 port map( A1 => n11952, A2 => n12422, B1 => n12361, B2 => 
                           n9012, ZN => n2420);
   U10737 : OAI22_X1 port map( A1 => n11952, A2 => n12426, B1 => n12361, B2 => 
                           n9011, ZN => n2421);
   U10738 : OAI22_X1 port map( A1 => n11952, A2 => n12430, B1 => n12361, B2 => 
                           n9010, ZN => n2422);
   U10739 : OAI22_X1 port map( A1 => n11952, A2 => n12434, B1 => n9867, B2 => 
                           n9009, ZN => n2423);
   U10740 : OAI22_X1 port map( A1 => n11952, A2 => n12438, B1 => n9867, B2 => 
                           n9008, ZN => n2424);
   U10741 : OAI22_X1 port map( A1 => n11952, A2 => n12442, B1 => n9867, B2 => 
                           n9007, ZN => n2425);
   U10742 : OAI22_X1 port map( A1 => n11952, A2 => n12446, B1 => n12361, B2 => 
                           n9006, ZN => n2426);
   U10743 : OAI22_X1 port map( A1 => n11952, A2 => n12450, B1 => n12361, B2 => 
                           n9005, ZN => n2427);
   U10744 : OAI22_X1 port map( A1 => n11952, A2 => n12454, B1 => n12361, B2 => 
                           n9004, ZN => n2428);
   U10745 : OAI22_X1 port map( A1 => n11952, A2 => n12458, B1 => n12361, B2 => 
                           n9003, ZN => n2429);
   U10746 : OAI22_X1 port map( A1 => n11952, A2 => n12462, B1 => n12361, B2 => 
                           n9002, ZN => n2430);
   U10747 : OAI22_X1 port map( A1 => n11951, A2 => n12466, B1 => n12361, B2 => 
                           n9001, ZN => n2431);
   U10748 : OAI22_X1 port map( A1 => n11951, A2 => n12470, B1 => n12361, B2 => 
                           n9000, ZN => n2432);
   U10749 : OAI22_X1 port map( A1 => n11951, A2 => n12474, B1 => n12361, B2 => 
                           n8999, ZN => n2433);
   U10750 : OAI22_X1 port map( A1 => n11951, A2 => n12478, B1 => n12361, B2 => 
                           n8998, ZN => n2434);
   U10751 : OAI22_X1 port map( A1 => n11951, A2 => n12482, B1 => n9867, B2 => 
                           n8997, ZN => n2435);
   U10752 : OAI22_X1 port map( A1 => n11951, A2 => n12486, B1 => n9867, B2 => 
                           n8996, ZN => n2436);
   U10753 : OAI22_X1 port map( A1 => n11951, A2 => n12490, B1 => n9867, B2 => 
                           n8995, ZN => n2437);
   U10754 : OAI22_X1 port map( A1 => n11951, A2 => n12494, B1 => n9867, B2 => 
                           n8994, ZN => n2438);
   U10755 : OAI22_X1 port map( A1 => n11951, A2 => n12498, B1 => n9867, B2 => 
                           n8993, ZN => n2439);
   U10756 : OAI22_X1 port map( A1 => n11951, A2 => n12502, B1 => n9867, B2 => 
                           n8992, ZN => n2440);
   U10757 : OAI22_X1 port map( A1 => n11951, A2 => n12506, B1 => n9867, B2 => 
                           n8991, ZN => n2441);
   U10758 : OAI22_X1 port map( A1 => n11951, A2 => n12514, B1 => n9867, B2 => 
                           n8990, ZN => n2442);
   U10759 : OAI22_X1 port map( A1 => n11929, A2 => n12387, B1 => n12329, B2 => 
                           n9277, ZN => n2155);
   U10760 : OAI22_X1 port map( A1 => n11929, A2 => n12391, B1 => n12329, B2 => 
                           n9276, ZN => n2156);
   U10761 : OAI22_X1 port map( A1 => n11929, A2 => n12395, B1 => n12329, B2 => 
                           n9275, ZN => n2157);
   U10762 : OAI22_X1 port map( A1 => n11929, A2 => n12399, B1 => n12329, B2 => 
                           n9274, ZN => n2158);
   U10763 : OAI22_X1 port map( A1 => n11929, A2 => n12403, B1 => n12329, B2 => 
                           n9273, ZN => n2159);
   U10764 : OAI22_X1 port map( A1 => n11929, A2 => n12407, B1 => n12329, B2 => 
                           n9272, ZN => n2160);
   U10765 : OAI22_X1 port map( A1 => n11929, A2 => n12411, B1 => n12329, B2 => 
                           n9271, ZN => n2161);
   U10766 : OAI22_X1 port map( A1 => n11929, A2 => n12415, B1 => n12329, B2 => 
                           n9270, ZN => n2162);
   U10767 : OAI22_X1 port map( A1 => n11928, A2 => n12419, B1 => n12329, B2 => 
                           n9269, ZN => n2163);
   U10768 : OAI22_X1 port map( A1 => n11928, A2 => n12423, B1 => n12329, B2 => 
                           n9268, ZN => n2164);
   U10769 : OAI22_X1 port map( A1 => n11928, A2 => n12427, B1 => n12329, B2 => 
                           n9267, ZN => n2165);
   U10770 : OAI22_X1 port map( A1 => n11928, A2 => n12431, B1 => n12329, B2 => 
                           n9266, ZN => n2166);
   U10771 : OAI22_X1 port map( A1 => n11928, A2 => n12435, B1 => n9877, B2 => 
                           n9265, ZN => n2167);
   U10772 : OAI22_X1 port map( A1 => n11928, A2 => n12439, B1 => n9877, B2 => 
                           n9264, ZN => n2168);
   U10773 : OAI22_X1 port map( A1 => n11928, A2 => n12443, B1 => n9877, B2 => 
                           n9263, ZN => n2169);
   U10774 : OAI22_X1 port map( A1 => n11928, A2 => n12447, B1 => n12329, B2 => 
                           n9262, ZN => n2170);
   U10775 : OAI22_X1 port map( A1 => n11928, A2 => n12451, B1 => n12329, B2 => 
                           n9261, ZN => n2171);
   U10776 : OAI22_X1 port map( A1 => n11928, A2 => n12455, B1 => n12329, B2 => 
                           n9260, ZN => n2172);
   U10777 : OAI22_X1 port map( A1 => n11928, A2 => n12459, B1 => n12329, B2 => 
                           n9259, ZN => n2173);
   U10778 : OAI22_X1 port map( A1 => n11928, A2 => n12463, B1 => n12329, B2 => 
                           n9258, ZN => n2174);
   U10779 : OAI22_X1 port map( A1 => n11927, A2 => n12467, B1 => n12329, B2 => 
                           n9257, ZN => n2175);
   U10780 : OAI22_X1 port map( A1 => n11927, A2 => n12471, B1 => n12329, B2 => 
                           n9256, ZN => n2176);
   U10781 : OAI22_X1 port map( A1 => n11927, A2 => n12475, B1 => n12329, B2 => 
                           n9255, ZN => n2177);
   U10782 : OAI22_X1 port map( A1 => n11927, A2 => n12479, B1 => n12329, B2 => 
                           n9254, ZN => n2178);
   U10783 : OAI22_X1 port map( A1 => n11927, A2 => n12483, B1 => n9877, B2 => 
                           n9253, ZN => n2179);
   U10784 : OAI22_X1 port map( A1 => n11927, A2 => n12487, B1 => n9877, B2 => 
                           n9252, ZN => n2180);
   U10785 : OAI22_X1 port map( A1 => n11927, A2 => n12491, B1 => n9877, B2 => 
                           n9251, ZN => n2181);
   U10786 : OAI22_X1 port map( A1 => n11927, A2 => n12495, B1 => n9877, B2 => 
                           n9250, ZN => n2182);
   U10787 : OAI22_X1 port map( A1 => n11927, A2 => n12499, B1 => n9877, B2 => 
                           n9249, ZN => n2183);
   U10788 : OAI22_X1 port map( A1 => n11927, A2 => n12503, B1 => n9877, B2 => 
                           n9248, ZN => n2184);
   U10789 : OAI22_X1 port map( A1 => n11927, A2 => n12507, B1 => n9877, B2 => 
                           n9247, ZN => n2185);
   U10790 : OAI22_X1 port map( A1 => n11927, A2 => n12515, B1 => n9877, B2 => 
                           n9246, ZN => n2186);
   U10791 : OAI22_X1 port map( A1 => n11950, A2 => n12386, B1 => n12357, B2 => 
                           n9053, ZN => n2379);
   U10792 : OAI22_X1 port map( A1 => n11950, A2 => n12390, B1 => n12357, B2 => 
                           n9052, ZN => n2380);
   U10793 : OAI22_X1 port map( A1 => n11950, A2 => n12394, B1 => n12357, B2 => 
                           n9051, ZN => n2381);
   U10794 : OAI22_X1 port map( A1 => n11950, A2 => n12398, B1 => n12357, B2 => 
                           n9050, ZN => n2382);
   U10795 : OAI22_X1 port map( A1 => n11950, A2 => n12402, B1 => n12357, B2 => 
                           n9049, ZN => n2383);
   U10796 : OAI22_X1 port map( A1 => n11950, A2 => n12406, B1 => n12357, B2 => 
                           n9048, ZN => n2384);
   U10797 : OAI22_X1 port map( A1 => n11950, A2 => n12410, B1 => n12357, B2 => 
                           n9047, ZN => n2385);
   U10798 : OAI22_X1 port map( A1 => n11950, A2 => n12414, B1 => n12357, B2 => 
                           n9046, ZN => n2386);
   U10799 : OAI22_X1 port map( A1 => n11949, A2 => n12418, B1 => n12357, B2 => 
                           n9045, ZN => n2387);
   U10800 : OAI22_X1 port map( A1 => n11949, A2 => n12422, B1 => n12357, B2 => 
                           n9044, ZN => n2388);
   U10801 : OAI22_X1 port map( A1 => n11949, A2 => n12426, B1 => n12357, B2 => 
                           n9043, ZN => n2389);
   U10802 : OAI22_X1 port map( A1 => n11949, A2 => n12430, B1 => n12357, B2 => 
                           n9042, ZN => n2390);
   U10803 : OAI22_X1 port map( A1 => n11949, A2 => n12434, B1 => n9868, B2 => 
                           n9041, ZN => n2391);
   U10804 : OAI22_X1 port map( A1 => n11949, A2 => n12438, B1 => n9868, B2 => 
                           n9040, ZN => n2392);
   U10805 : OAI22_X1 port map( A1 => n11949, A2 => n12442, B1 => n9868, B2 => 
                           n9039, ZN => n2393);
   U10806 : OAI22_X1 port map( A1 => n11949, A2 => n12446, B1 => n12357, B2 => 
                           n9038, ZN => n2394);
   U10807 : OAI22_X1 port map( A1 => n11949, A2 => n12450, B1 => n12357, B2 => 
                           n9037, ZN => n2395);
   U10808 : OAI22_X1 port map( A1 => n11949, A2 => n12454, B1 => n12357, B2 => 
                           n9036, ZN => n2396);
   U10809 : OAI22_X1 port map( A1 => n11949, A2 => n12458, B1 => n12357, B2 => 
                           n9035, ZN => n2397);
   U10810 : OAI22_X1 port map( A1 => n11949, A2 => n12462, B1 => n12357, B2 => 
                           n9034, ZN => n2398);
   U10811 : OAI22_X1 port map( A1 => n11948, A2 => n12466, B1 => n12357, B2 => 
                           n9033, ZN => n2399);
   U10812 : OAI22_X1 port map( A1 => n11948, A2 => n12470, B1 => n12357, B2 => 
                           n9032, ZN => n2400);
   U10813 : OAI22_X1 port map( A1 => n11948, A2 => n12474, B1 => n12357, B2 => 
                           n9031, ZN => n2401);
   U10814 : OAI22_X1 port map( A1 => n11948, A2 => n12478, B1 => n12357, B2 => 
                           n9030, ZN => n2402);
   U10815 : OAI22_X1 port map( A1 => n11948, A2 => n12482, B1 => n9868, B2 => 
                           n9029, ZN => n2403);
   U10816 : OAI22_X1 port map( A1 => n11948, A2 => n12486, B1 => n9868, B2 => 
                           n9028, ZN => n2404);
   U10817 : OAI22_X1 port map( A1 => n11948, A2 => n12490, B1 => n9868, B2 => 
                           n9027, ZN => n2405);
   U10818 : OAI22_X1 port map( A1 => n11948, A2 => n12494, B1 => n9868, B2 => 
                           n9026, ZN => n2406);
   U10819 : OAI22_X1 port map( A1 => n11948, A2 => n12498, B1 => n9868, B2 => 
                           n9025, ZN => n2407);
   U10820 : OAI22_X1 port map( A1 => n11948, A2 => n12502, B1 => n9868, B2 => 
                           n9024, ZN => n2408);
   U10821 : OAI22_X1 port map( A1 => n11948, A2 => n12506, B1 => n9868, B2 => 
                           n9023, ZN => n2409);
   U10822 : OAI22_X1 port map( A1 => n11948, A2 => n12514, B1 => n9868, B2 => 
                           n9022, ZN => n2410);
   U10823 : OAI22_X1 port map( A1 => n11881, A2 => n12388, B1 => n12265, B2 => 
                           n9789, ZN => n1643);
   U10824 : OAI22_X1 port map( A1 => n11881, A2 => n12392, B1 => n12265, B2 => 
                           n9788, ZN => n1644);
   U10825 : OAI22_X1 port map( A1 => n11881, A2 => n12396, B1 => n12265, B2 => 
                           n9787, ZN => n1645);
   U10826 : OAI22_X1 port map( A1 => n11881, A2 => n12400, B1 => n12265, B2 => 
                           n9786, ZN => n1646);
   U10827 : OAI22_X1 port map( A1 => n11881, A2 => n12404, B1 => n12265, B2 => 
                           n9785, ZN => n1647);
   U10828 : OAI22_X1 port map( A1 => n11881, A2 => n12408, B1 => n12265, B2 => 
                           n9784, ZN => n1648);
   U10829 : OAI22_X1 port map( A1 => n11881, A2 => n12412, B1 => n12265, B2 => 
                           n9783, ZN => n1649);
   U10830 : OAI22_X1 port map( A1 => n11881, A2 => n12416, B1 => n12265, B2 => 
                           n9782, ZN => n1650);
   U10831 : OAI22_X1 port map( A1 => n11880, A2 => n12420, B1 => n12265, B2 => 
                           n9781, ZN => n1651);
   U10832 : OAI22_X1 port map( A1 => n11880, A2 => n12424, B1 => n12265, B2 => 
                           n9780, ZN => n1652);
   U10833 : OAI22_X1 port map( A1 => n11880, A2 => n12428, B1 => n12265, B2 => 
                           n9779, ZN => n1653);
   U10834 : OAI22_X1 port map( A1 => n11880, A2 => n12432, B1 => n12265, B2 => 
                           n9778, ZN => n1654);
   U10835 : OAI22_X1 port map( A1 => n11880, A2 => n12436, B1 => n9898, B2 => 
                           n9777, ZN => n1655);
   U10836 : OAI22_X1 port map( A1 => n11880, A2 => n12440, B1 => n9898, B2 => 
                           n9776, ZN => n1656);
   U10837 : OAI22_X1 port map( A1 => n11880, A2 => n12444, B1 => n9898, B2 => 
                           n9775, ZN => n1657);
   U10838 : OAI22_X1 port map( A1 => n11880, A2 => n12448, B1 => n12265, B2 => 
                           n9774, ZN => n1658);
   U10839 : OAI22_X1 port map( A1 => n11880, A2 => n12452, B1 => n12265, B2 => 
                           n9773, ZN => n1659);
   U10840 : OAI22_X1 port map( A1 => n11880, A2 => n12456, B1 => n12265, B2 => 
                           n9772, ZN => n1660);
   U10841 : OAI22_X1 port map( A1 => n11880, A2 => n12460, B1 => n12265, B2 => 
                           n9771, ZN => n1661);
   U10842 : OAI22_X1 port map( A1 => n11880, A2 => n12464, B1 => n12265, B2 => 
                           n9770, ZN => n1662);
   U10843 : OAI22_X1 port map( A1 => n11879, A2 => n12468, B1 => n12265, B2 => 
                           n9769, ZN => n1663);
   U10844 : OAI22_X1 port map( A1 => n11879, A2 => n12472, B1 => n12265, B2 => 
                           n9768, ZN => n1664);
   U10845 : OAI22_X1 port map( A1 => n11879, A2 => n12476, B1 => n12265, B2 => 
                           n9767, ZN => n1665);
   U10846 : OAI22_X1 port map( A1 => n11879, A2 => n12480, B1 => n12265, B2 => 
                           n9766, ZN => n1666);
   U10847 : OAI22_X1 port map( A1 => n11879, A2 => n12484, B1 => n9898, B2 => 
                           n9765, ZN => n1667);
   U10848 : OAI22_X1 port map( A1 => n11879, A2 => n12488, B1 => n9898, B2 => 
                           n9764, ZN => n1668);
   U10849 : OAI22_X1 port map( A1 => n11879, A2 => n12492, B1 => n9898, B2 => 
                           n9763, ZN => n1669);
   U10850 : OAI22_X1 port map( A1 => n11879, A2 => n12496, B1 => n9898, B2 => 
                           n9762, ZN => n1670);
   U10851 : OAI22_X1 port map( A1 => n11879, A2 => n12500, B1 => n9898, B2 => 
                           n9761, ZN => n1671);
   U10852 : OAI22_X1 port map( A1 => n11879, A2 => n12504, B1 => n9898, B2 => 
                           n9760, ZN => n1672);
   U10853 : OAI22_X1 port map( A1 => n11879, A2 => n12508, B1 => n9898, B2 => 
                           n9759, ZN => n1673);
   U10854 : OAI22_X1 port map( A1 => n11879, A2 => n12516, B1 => n9898, B2 => 
                           n9758, ZN => n1674);
   U10855 : OAI22_X1 port map( A1 => n11920, A2 => n12387, B1 => n12317, B2 => 
                           n9373, ZN => n2059);
   U10856 : OAI22_X1 port map( A1 => n11920, A2 => n12391, B1 => n12317, B2 => 
                           n9372, ZN => n2060);
   U10857 : OAI22_X1 port map( A1 => n11920, A2 => n12395, B1 => n12317, B2 => 
                           n9371, ZN => n2061);
   U10858 : OAI22_X1 port map( A1 => n11920, A2 => n12399, B1 => n12317, B2 => 
                           n9370, ZN => n2062);
   U10859 : OAI22_X1 port map( A1 => n11920, A2 => n12403, B1 => n12317, B2 => 
                           n9369, ZN => n2063);
   U10860 : OAI22_X1 port map( A1 => n11920, A2 => n12407, B1 => n12317, B2 => 
                           n9368, ZN => n2064);
   U10861 : OAI22_X1 port map( A1 => n11920, A2 => n12411, B1 => n12317, B2 => 
                           n9367, ZN => n2065);
   U10862 : OAI22_X1 port map( A1 => n11920, A2 => n12415, B1 => n12317, B2 => 
                           n9366, ZN => n2066);
   U10863 : OAI22_X1 port map( A1 => n11919, A2 => n12419, B1 => n12317, B2 => 
                           n9365, ZN => n2067);
   U10864 : OAI22_X1 port map( A1 => n11919, A2 => n12423, B1 => n12317, B2 => 
                           n9364, ZN => n2068);
   U10865 : OAI22_X1 port map( A1 => n11919, A2 => n12427, B1 => n12317, B2 => 
                           n9363, ZN => n2069);
   U10866 : OAI22_X1 port map( A1 => n11919, A2 => n12431, B1 => n12317, B2 => 
                           n9362, ZN => n2070);
   U10867 : OAI22_X1 port map( A1 => n11919, A2 => n12435, B1 => n9881, B2 => 
                           n9361, ZN => n2071);
   U10868 : OAI22_X1 port map( A1 => n11919, A2 => n12439, B1 => n9881, B2 => 
                           n9360, ZN => n2072);
   U10869 : OAI22_X1 port map( A1 => n11919, A2 => n12443, B1 => n9881, B2 => 
                           n9359, ZN => n2073);
   U10870 : OAI22_X1 port map( A1 => n11919, A2 => n12447, B1 => n12317, B2 => 
                           n9358, ZN => n2074);
   U10871 : OAI22_X1 port map( A1 => n11919, A2 => n12451, B1 => n12317, B2 => 
                           n9357, ZN => n2075);
   U10872 : OAI22_X1 port map( A1 => n11919, A2 => n12455, B1 => n12317, B2 => 
                           n9356, ZN => n2076);
   U10873 : OAI22_X1 port map( A1 => n11919, A2 => n12459, B1 => n12317, B2 => 
                           n9355, ZN => n2077);
   U10874 : OAI22_X1 port map( A1 => n11919, A2 => n12463, B1 => n12317, B2 => 
                           n9354, ZN => n2078);
   U10875 : OAI22_X1 port map( A1 => n11918, A2 => n12467, B1 => n12317, B2 => 
                           n9353, ZN => n2079);
   U10876 : OAI22_X1 port map( A1 => n11918, A2 => n12471, B1 => n12317, B2 => 
                           n9352, ZN => n2080);
   U10877 : OAI22_X1 port map( A1 => n11918, A2 => n12475, B1 => n12317, B2 => 
                           n9351, ZN => n2081);
   U10878 : OAI22_X1 port map( A1 => n11918, A2 => n12479, B1 => n12317, B2 => 
                           n9350, ZN => n2082);
   U10879 : OAI22_X1 port map( A1 => n11918, A2 => n12483, B1 => n9881, B2 => 
                           n9349, ZN => n2083);
   U10880 : OAI22_X1 port map( A1 => n11918, A2 => n12487, B1 => n9881, B2 => 
                           n9348, ZN => n2084);
   U10881 : OAI22_X1 port map( A1 => n11918, A2 => n12491, B1 => n9881, B2 => 
                           n9347, ZN => n2085);
   U10882 : OAI22_X1 port map( A1 => n11918, A2 => n12495, B1 => n9881, B2 => 
                           n9346, ZN => n2086);
   U10883 : OAI22_X1 port map( A1 => n11918, A2 => n12499, B1 => n9881, B2 => 
                           n9345, ZN => n2087);
   U10884 : OAI22_X1 port map( A1 => n11918, A2 => n12503, B1 => n9881, B2 => 
                           n9344, ZN => n2088);
   U10885 : OAI22_X1 port map( A1 => n11918, A2 => n12507, B1 => n9881, B2 => 
                           n9343, ZN => n2089);
   U10886 : OAI22_X1 port map( A1 => n11918, A2 => n12515, B1 => n9881, B2 => 
                           n9342, ZN => n2090);
   U10887 : OAI22_X1 port map( A1 => n11876, A2 => n9821, B1 => n12261, B2 => 
                           n12388, ZN => n1611);
   U10888 : OAI22_X1 port map( A1 => n11876, A2 => n9820, B1 => n12260, B2 => 
                           n12392, ZN => n1612);
   U10889 : OAI22_X1 port map( A1 => n11876, A2 => n9819, B1 => n12261, B2 => 
                           n12396, ZN => n1613);
   U10890 : OAI22_X1 port map( A1 => n11876, A2 => n9818, B1 => n12260, B2 => 
                           n12400, ZN => n1614);
   U10891 : OAI22_X1 port map( A1 => n11876, A2 => n9817, B1 => n12261, B2 => 
                           n12404, ZN => n1615);
   U10892 : OAI22_X1 port map( A1 => n11876, A2 => n9816, B1 => n12260, B2 => 
                           n12408, ZN => n1616);
   U10893 : OAI22_X1 port map( A1 => n11876, A2 => n9815, B1 => n12261, B2 => 
                           n12412, ZN => n1617);
   U10894 : OAI22_X1 port map( A1 => n11876, A2 => n9814, B1 => n12260, B2 => 
                           n12416, ZN => n1618);
   U10895 : OAI22_X1 port map( A1 => n11876, A2 => n9813, B1 => n12261, B2 => 
                           n12420, ZN => n1619);
   U10896 : OAI22_X1 port map( A1 => n11876, A2 => n9812, B1 => n12261, B2 => 
                           n12424, ZN => n1620);
   U10897 : OAI22_X1 port map( A1 => n11876, A2 => n9811, B1 => n12261, B2 => 
                           n12428, ZN => n1621);
   U10898 : OAI22_X1 port map( A1 => n11876, A2 => n9810, B1 => n12261, B2 => 
                           n12432, ZN => n1622);
   U10899 : OAI22_X1 port map( A1 => n11877, A2 => n9809, B1 => n12261, B2 => 
                           n12436, ZN => n1623);
   U10900 : OAI22_X1 port map( A1 => n11877, A2 => n9808, B1 => n12261, B2 => 
                           n12440, ZN => n1624);
   U10901 : OAI22_X1 port map( A1 => n11877, A2 => n9807, B1 => n12261, B2 => 
                           n12444, ZN => n1625);
   U10902 : OAI22_X1 port map( A1 => n11877, A2 => n9806, B1 => n12261, B2 => 
                           n12448, ZN => n1626);
   U10903 : OAI22_X1 port map( A1 => n11877, A2 => n9805, B1 => n12261, B2 => 
                           n12452, ZN => n1627);
   U10904 : OAI22_X1 port map( A1 => n11877, A2 => n9804, B1 => n12261, B2 => 
                           n12456, ZN => n1628);
   U10905 : OAI22_X1 port map( A1 => n11877, A2 => n9803, B1 => n12261, B2 => 
                           n12460, ZN => n1629);
   U10906 : OAI22_X1 port map( A1 => n11877, A2 => n9802, B1 => n12261, B2 => 
                           n12464, ZN => n1630);
   U10907 : OAI22_X1 port map( A1 => n11877, A2 => n9801, B1 => n12260, B2 => 
                           n12468, ZN => n1631);
   U10908 : OAI22_X1 port map( A1 => n11877, A2 => n9800, B1 => n12260, B2 => 
                           n12472, ZN => n1632);
   U10909 : OAI22_X1 port map( A1 => n11877, A2 => n9799, B1 => n12260, B2 => 
                           n12476, ZN => n1633);
   U10910 : OAI22_X1 port map( A1 => n11877, A2 => n9798, B1 => n12260, B2 => 
                           n12480, ZN => n1634);
   U10911 : OAI22_X1 port map( A1 => n11878, A2 => n9797, B1 => n12260, B2 => 
                           n12484, ZN => n1635);
   U10912 : OAI22_X1 port map( A1 => n11878, A2 => n9796, B1 => n12260, B2 => 
                           n12488, ZN => n1636);
   U10913 : OAI22_X1 port map( A1 => n11878, A2 => n9795, B1 => n12260, B2 => 
                           n12492, ZN => n1637);
   U10914 : OAI22_X1 port map( A1 => n11878, A2 => n9794, B1 => n12260, B2 => 
                           n12496, ZN => n1638);
   U10915 : OAI22_X1 port map( A1 => n11878, A2 => n9793, B1 => n12260, B2 => 
                           n12500, ZN => n1639);
   U10916 : OAI22_X1 port map( A1 => n11878, A2 => n9792, B1 => n12260, B2 => 
                           n12504, ZN => n1640);
   U10917 : OAI22_X1 port map( A1 => n11878, A2 => n9791, B1 => n12260, B2 => 
                           n12508, ZN => n1641);
   U10918 : OAI22_X1 port map( A1 => n11878, A2 => n9790, B1 => n12260, B2 => 
                           n12516, ZN => n1642);
   U10919 : OAI21_X1 port map( B1 => n11870, B2 => n4742, A => n11973, ZN => 
                           n1483);
   U10920 : OAI21_X1 port map( B1 => n11872, B2 => n4744, A => n11973, ZN => 
                           n1485);
   U10921 : OAI21_X1 port map( B1 => n11872, B2 => n4746, A => n11973, ZN => 
                           n1487);
   U10922 : OAI21_X1 port map( B1 => n11872, B2 => n4748, A => n11973, ZN => 
                           n1489);
   U10923 : OAI21_X1 port map( B1 => n11872, B2 => n4750, A => n11973, ZN => 
                           n1491);
   U10924 : OAI21_X1 port map( B1 => n11872, B2 => n4752, A => n11973, ZN => 
                           n1493);
   U10925 : OAI21_X1 port map( B1 => n11872, B2 => n4754, A => n11973, ZN => 
                           n1495);
   U10926 : OAI21_X1 port map( B1 => n11872, B2 => n4756, A => n11973, ZN => 
                           n1497);
   U10927 : OAI21_X1 port map( B1 => n11871, B2 => n4758, A => n11973, ZN => 
                           n1499);
   U10928 : OAI21_X1 port map( B1 => n11871, B2 => n4760, A => n11973, ZN => 
                           n1501);
   U10929 : OAI21_X1 port map( B1 => n11871, B2 => n4762, A => n11973, ZN => 
                           n1503);
   U10930 : OAI21_X1 port map( B1 => n11871, B2 => n4764, A => n11973, ZN => 
                           n1505);
   U10931 : OAI21_X1 port map( B1 => n11871, B2 => n4766, A => n11974, ZN => 
                           n1507);
   U10932 : OAI21_X1 port map( B1 => n11871, B2 => n4768, A => n11974, ZN => 
                           n1509);
   U10933 : OAI21_X1 port map( B1 => n11871, B2 => n4770, A => n11974, ZN => 
                           n1511);
   U10934 : OAI21_X1 port map( B1 => n11871, B2 => n4772, A => n11974, ZN => 
                           n1513);
   U10935 : OAI21_X1 port map( B1 => n11871, B2 => n4774, A => n11974, ZN => 
                           n1515);
   U10936 : OAI21_X1 port map( B1 => n11871, B2 => n4776, A => n11974, ZN => 
                           n1517);
   U10937 : OAI21_X1 port map( B1 => n11871, B2 => n4778, A => n11974, ZN => 
                           n1519);
   U10938 : OAI21_X1 port map( B1 => n11870, B2 => n4780, A => n11974, ZN => 
                           n1521);
   U10939 : OAI21_X1 port map( B1 => n11870, B2 => n4782, A => n11974, ZN => 
                           n1523);
   U10940 : OAI21_X1 port map( B1 => n11870, B2 => n4784, A => n11974, ZN => 
                           n1525);
   U10941 : OAI21_X1 port map( B1 => n11870, B2 => n4786, A => n11974, ZN => 
                           n1527);
   U10942 : OAI21_X1 port map( B1 => n11870, B2 => n4788, A => n11974, ZN => 
                           n1529);
   U10943 : OAI21_X1 port map( B1 => n11871, B2 => n4790, A => n11975, ZN => 
                           n1531);
   U10944 : OAI21_X1 port map( B1 => n11871, B2 => n4792, A => n11975, ZN => 
                           n1533);
   U10945 : OAI21_X1 port map( B1 => n11870, B2 => n4794, A => n11975, ZN => 
                           n1535);
   U10946 : OAI21_X1 port map( B1 => n11870, B2 => n4796, A => n11975, ZN => 
                           n1537);
   U10947 : OAI21_X1 port map( B1 => n11870, B2 => n4798, A => n11975, ZN => 
                           n1539);
   U10948 : OAI21_X1 port map( B1 => n11870, B2 => n4800, A => n11975, ZN => 
                           n1541);
   U10949 : OAI21_X1 port map( B1 => n11870, B2 => n4802, A => n11975, ZN => 
                           n1543);
   U10950 : OAI21_X1 port map( B1 => n11870, B2 => n4804, A => n11975, ZN => 
                           n1545);
   U10951 : OAI21_X1 port map( B1 => n11873, B2 => n4806, A => n12117, ZN => 
                           n1547);
   U10952 : OAI21_X1 port map( B1 => n11875, B2 => n4808, A => n12117, ZN => 
                           n1549);
   U10953 : OAI21_X1 port map( B1 => n11875, B2 => n4810, A => n12117, ZN => 
                           n1551);
   U10954 : OAI21_X1 port map( B1 => n11875, B2 => n4812, A => n12117, ZN => 
                           n1553);
   U10955 : OAI21_X1 port map( B1 => n11875, B2 => n4814, A => n12117, ZN => 
                           n1555);
   U10956 : OAI21_X1 port map( B1 => n11875, B2 => n4816, A => n12117, ZN => 
                           n1557);
   U10957 : OAI21_X1 port map( B1 => n11875, B2 => n4818, A => n12117, ZN => 
                           n1559);
   U10958 : OAI21_X1 port map( B1 => n11875, B2 => n4820, A => n12117, ZN => 
                           n1561);
   U10959 : OAI21_X1 port map( B1 => n11874, B2 => n4822, A => n12117, ZN => 
                           n1563);
   U10960 : OAI21_X1 port map( B1 => n11874, B2 => n4824, A => n12117, ZN => 
                           n1565);
   U10961 : OAI21_X1 port map( B1 => n11874, B2 => n4826, A => n12117, ZN => 
                           n1567);
   U10962 : OAI21_X1 port map( B1 => n11874, B2 => n4828, A => n12117, ZN => 
                           n1569);
   U10963 : OAI21_X1 port map( B1 => n11874, B2 => n4830, A => n12118, ZN => 
                           n1571);
   U10964 : OAI21_X1 port map( B1 => n11874, B2 => n4832, A => n12118, ZN => 
                           n1573);
   U10965 : OAI21_X1 port map( B1 => n11874, B2 => n4834, A => n12118, ZN => 
                           n1575);
   U10966 : OAI21_X1 port map( B1 => n11874, B2 => n4836, A => n12118, ZN => 
                           n1577);
   U10967 : OAI21_X1 port map( B1 => n11874, B2 => n4838, A => n12118, ZN => 
                           n1579);
   U10968 : OAI21_X1 port map( B1 => n11874, B2 => n4840, A => n12118, ZN => 
                           n1581);
   U10969 : OAI21_X1 port map( B1 => n11874, B2 => n4842, A => n12118, ZN => 
                           n1583);
   U10970 : OAI21_X1 port map( B1 => n11873, B2 => n4844, A => n12118, ZN => 
                           n1585);
   U10971 : OAI21_X1 port map( B1 => n11873, B2 => n4846, A => n12118, ZN => 
                           n1587);
   U10972 : OAI21_X1 port map( B1 => n11873, B2 => n4848, A => n12118, ZN => 
                           n1589);
   U10973 : OAI21_X1 port map( B1 => n11873, B2 => n4850, A => n12118, ZN => 
                           n1591);
   U10974 : OAI21_X1 port map( B1 => n11873, B2 => n4852, A => n12118, ZN => 
                           n1593);
   U10975 : OAI21_X1 port map( B1 => n11874, B2 => n4854, A => n12119, ZN => 
                           n1595);
   U10976 : OAI21_X1 port map( B1 => n11874, B2 => n4856, A => n12119, ZN => 
                           n1597);
   U10977 : OAI21_X1 port map( B1 => n11873, B2 => n4858, A => n12119, ZN => 
                           n1599);
   U10978 : OAI21_X1 port map( B1 => n11873, B2 => n4860, A => n12119, ZN => 
                           n1601);
   U10979 : OAI21_X1 port map( B1 => n11873, B2 => n4862, A => n12119, ZN => 
                           n1603);
   U10980 : OAI21_X1 port map( B1 => n11873, B2 => n4864, A => n12119, ZN => 
                           n1605);
   U10981 : OAI21_X1 port map( B1 => n11873, B2 => n4866, A => n12119, ZN => 
                           n1607);
   U10982 : OAI21_X1 port map( B1 => n11873, B2 => n4868, A => n12119, ZN => 
                           n1609);
   U10983 : NOR2_X1 port map( A1 => ADD_RD2(4), A2 => ADD_RD2(3), ZN => n11095)
                           ;
   U10984 : NOR2_X1 port map( A1 => n8794, A2 => ADD_RD2(4), ZN => n11094);
   U10985 : NOR2_X1 port map( A1 => ADD_RD1(4), A2 => ADD_RD1(3), ZN => n10495)
                           ;
   U10986 : NOR2_X1 port map( A1 => n8790, A2 => ADD_RD1(4), ZN => n10494);
   U10987 : NOR3_X1 port map( A1 => n8796, A2 => ADD_RD2(2), A3 => n8797, ZN =>
                           n11072);
   U10988 : NOR3_X1 port map( A1 => n8792, A2 => ADD_RD1(2), A3 => n8793, ZN =>
                           n10472);
   U10989 : NOR3_X1 port map( A1 => ADD_RD2(0), A2 => ADD_RD2(1), A3 => n8795, 
                           ZN => n11069);
   U10990 : NOR3_X1 port map( A1 => ADD_RD1(0), A2 => ADD_RD1(1), A3 => n8791, 
                           ZN => n10469);
   U10991 : NOR3_X1 port map( A1 => ADD_RD2(1), A2 => ADD_RD2(2), A3 => n8797, 
                           ZN => n11073);
   U10992 : NOR3_X1 port map( A1 => ADD_RD1(1), A2 => ADD_RD1(2), A3 => n8793, 
                           ZN => n10473);
   U10993 : NOR3_X1 port map( A1 => ADD_RD2(0), A2 => ADD_RD2(2), A3 => n8796, 
                           ZN => n11075);
   U10994 : NOR3_X1 port map( A1 => ADD_RD2(1), A2 => ADD_RD2(2), A3 => 
                           ADD_RD2(0), ZN => n11071);
   U10995 : NOR3_X1 port map( A1 => ADD_RD1(0), A2 => ADD_RD1(2), A3 => n8792, 
                           ZN => n10475);
   U10996 : NOR3_X1 port map( A1 => ADD_RD1(1), A2 => ADD_RD1(2), A3 => 
                           ADD_RD1(0), ZN => n10471);
   U10997 : NOR3_X1 port map( A1 => n8796, A2 => ADD_RD2(0), A3 => n8795, ZN =>
                           n11070);
   U10998 : NOR3_X1 port map( A1 => n8792, A2 => ADD_RD1(0), A3 => n8791, ZN =>
                           n10470);
   U10999 : NOR3_X1 port map( A1 => n8795, A2 => ADD_RD2(1), A3 => n8797, ZN =>
                           n11076);
   U11000 : NOR3_X1 port map( A1 => n8791, A2 => ADD_RD1(1), A3 => n8793, ZN =>
                           n10476);
   U11001 : NOR3_X1 port map( A1 => n8782, A2 => ADD_WR(4), A3 => n8783, ZN => 
                           n9863);
   U11002 : INV_X1 port map( A => ENABLE, ZN => n8782);
   U11003 : NAND2_X1 port map( A1 => ADD_WR(0), A2 => n8786, ZN => n9858);
   U11004 : NAND2_X1 port map( A1 => ADD_WR(1), A2 => ADD_WR(0), ZN => n9862);
   U11005 : NAND2_X1 port map( A1 => ADD_WR(1), A2 => n8789, ZN => n9860);
   U11006 : INV_X1 port map( A => WR, ZN => n8783);
   U11007 : XNOR2_X1 port map( A => n8789, B => ADD_RD2(0), ZN => n11088);
   U11008 : XNOR2_X1 port map( A => n8789, B => ADD_RD1(0), ZN => n10488);
   U11009 : XNOR2_X1 port map( A => ADD_WR(4), B => ADD_RD2(4), ZN => n11083);
   U11010 : XNOR2_X1 port map( A => ADD_WR(4), B => ADD_RD1(4), ZN => n10483);
   U11011 : NAND4_X1 port map( A1 => n11083, A2 => n8787, A3 => n11084, A4 => 
                           n11085, ZN => n11082);
   U11012 : INV_X1 port map( A => n11088, ZN => n8787);
   U11013 : NAND4_X1 port map( A1 => n10483, A2 => n8788, A3 => n10484, A4 => 
                           n10485, ZN => n10482);
   U11014 : INV_X1 port map( A => n10488, ZN => n8788);
   U11015 : AND2_X1 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(4), ZN => n11077)
                           ;
   U11016 : AND2_X1 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(4), ZN => n10477)
                           ;
   U11017 : AND2_X1 port map( A1 => ADD_RD2(4), A2 => n8794, ZN => n11068);
   U11018 : AND2_X1 port map( A1 => ADD_RD1(4), A2 => n8790, ZN => n10468);
   U11019 : INV_X1 port map( A => ADD_RD2(2), ZN => n8795);
   U11020 : INV_X1 port map( A => ADD_RD1(2), ZN => n8791);
   U11021 : INV_X1 port map( A => ADD_WR(0), ZN => n8789);
   U11022 : INV_X1 port map( A => ADD_RD2(0), ZN => n8797);
   U11023 : INV_X1 port map( A => ADD_RD1(0), ZN => n8793);
   U11024 : INV_X1 port map( A => ADD_RD2(1), ZN => n8796);
   U11025 : INV_X1 port map( A => ADD_RD1(1), ZN => n8792);
   U11026 : AND3_X1 port map( A1 => WR, A2 => ENABLE, A3 => ADD_WR(4), ZN => 
                           n9884);
   U11027 : INV_X1 port map( A => ADD_WR(3), ZN => n8784);
   U11028 : INV_X1 port map( A => ADD_WR(2), ZN => n8785);
   U11029 : INV_X1 port map( A => ADD_WR(1), ZN => n8786);
   U11030 : NAND2_X1 port map( A1 => DATAIN(0), A2 => n12519, ZN => n9854);
   U11031 : NAND2_X1 port map( A1 => DATAIN(1), A2 => n12519, ZN => n9853);
   U11032 : NAND2_X1 port map( A1 => DATAIN(2), A2 => n12519, ZN => n9852);
   U11033 : NAND2_X1 port map( A1 => DATAIN(3), A2 => n12519, ZN => n9851);
   U11034 : NAND2_X1 port map( A1 => DATAIN(4), A2 => n12519, ZN => n9850);
   U11035 : NAND2_X1 port map( A1 => DATAIN(5), A2 => n12519, ZN => n9849);
   U11036 : NAND2_X1 port map( A1 => DATAIN(6), A2 => n12519, ZN => n9848);
   U11037 : NAND2_X1 port map( A1 => DATAIN(7), A2 => n12519, ZN => n9847);
   U11038 : NAND2_X1 port map( A1 => DATAIN(8), A2 => n12518, ZN => n9846);
   U11039 : NAND2_X1 port map( A1 => DATAIN(9), A2 => n12518, ZN => n9845);
   U11040 : NAND2_X1 port map( A1 => DATAIN(10), A2 => n12518, ZN => n9844);
   U11041 : NAND2_X1 port map( A1 => DATAIN(11), A2 => n12518, ZN => n9843);
   U11042 : NAND2_X1 port map( A1 => DATAIN(12), A2 => n12518, ZN => n9842);
   U11043 : NAND2_X1 port map( A1 => DATAIN(13), A2 => n12518, ZN => n9841);
   U11044 : NAND2_X1 port map( A1 => DATAIN(14), A2 => n12518, ZN => n9840);
   U11045 : NAND2_X1 port map( A1 => DATAIN(15), A2 => n12518, ZN => n9839);
   U11046 : NAND2_X1 port map( A1 => DATAIN(16), A2 => n12518, ZN => n9838);
   U11047 : NAND2_X1 port map( A1 => DATAIN(17), A2 => n12518, ZN => n9837);
   U11048 : NAND2_X1 port map( A1 => DATAIN(18), A2 => n12518, ZN => n9836);
   U11049 : NAND2_X1 port map( A1 => DATAIN(19), A2 => n12518, ZN => n9835);
   U11050 : NAND2_X1 port map( A1 => DATAIN(20), A2 => n12517, ZN => n9834);
   U11051 : NAND2_X1 port map( A1 => DATAIN(21), A2 => n12517, ZN => n9833);
   U11052 : NAND2_X1 port map( A1 => DATAIN(22), A2 => n12517, ZN => n9832);
   U11053 : NAND2_X1 port map( A1 => DATAIN(23), A2 => n12517, ZN => n9831);
   U11054 : NAND2_X1 port map( A1 => DATAIN(24), A2 => n12517, ZN => n9830);
   U11055 : NAND2_X1 port map( A1 => DATAIN(25), A2 => n12517, ZN => n9829);
   U11056 : NAND2_X1 port map( A1 => DATAIN(26), A2 => n12517, ZN => n9828);
   U11057 : NAND2_X1 port map( A1 => DATAIN(27), A2 => n12517, ZN => n9827);
   U11058 : NAND2_X1 port map( A1 => DATAIN(28), A2 => n12517, ZN => n9826);
   U11059 : NAND2_X1 port map( A1 => DATAIN(29), A2 => n12517, ZN => n9825);
   U11060 : NAND2_X1 port map( A1 => DATAIN(30), A2 => n12517, ZN => n9824);
   U11061 : NAND2_X1 port map( A1 => DATAIN(31), A2 => n12517, ZN => n9822);
   U11062 : OR2_X1 port map( A1 => n10521, A2 => RD2, ZN => n10552);
   U11063 : OR2_X1 port map( A1 => n9921, A2 => RD1, ZN => n9952);
   U11064 : INV_X1 port map( A => ADD_RD2(3), ZN => n8794);
   U11065 : INV_X1 port map( A => ADD_RD1(3), ZN => n8790);
   U11066 : INV_X1 port map( A => RESET, ZN => n8781);
   U11067 : INV_X1 port map( A => n10521, ZN => n12059);
   U11068 : OAI211_X1 port map( C1 => RD2, C2 => n8783, A => n12519, B => 
                           ENABLE, ZN => n10521);
   U11069 : INV_X1 port map( A => n9921, ZN => n12203);
   U11070 : OAI211_X1 port map( C1 => RD1, C2 => n8783, A => n12519, B => 
                           ENABLE, ZN => n9921);

end SYN_Behavioral;
